////
//// Part of the ISPD 2013 Discrete Gate Sizing Contest Benchmark Suite. 
//// Please cite the following paper if you refer to these benchmarks in a publication:
//// M. M. Ozdal, C. Amin, A. Ayupov, S. Burns, G. Wilke, C. Zhuo, 
//// "An Improved Benchmark Suite for the ISPD-2013 Discrete Cell Sizing Contest"
//// Proc. ACM International Symposium on Physical Design, 2013.
////
//// This benchmark was generated for the ISPD 2013 contest using Cadence C-to-Silicon Compiler and Encounter Digital Implementation System 
////

module fft (
ispd_clk,
rst,
x_in_0_0,
x_in_0_1,
x_in_0_10,
x_in_0_11,
x_in_0_12,
x_in_0_13,
x_in_0_14,
x_in_0_15,
x_in_0_2,
x_in_0_3,
x_in_0_4,
x_in_0_5,
x_in_0_6,
x_in_0_7,
x_in_0_8,
x_in_0_9,
x_in_10_0,
x_in_10_1,
x_in_10_10,
x_in_10_11,
x_in_10_12,
x_in_10_13,
x_in_10_14,
x_in_10_15,
x_in_10_2,
x_in_10_3,
x_in_10_4,
x_in_10_5,
x_in_10_6,
x_in_10_7,
x_in_10_8,
x_in_10_9,
x_in_11_0,
x_in_11_1,
x_in_11_10,
x_in_11_11,
x_in_11_12,
x_in_11_13,
x_in_11_14,
x_in_11_15,
x_in_11_2,
x_in_11_3,
x_in_11_4,
x_in_11_5,
x_in_11_6,
x_in_11_7,
x_in_11_8,
x_in_11_9,
x_in_12_0,
x_in_12_1,
x_in_12_10,
x_in_12_11,
x_in_12_12,
x_in_12_13,
x_in_12_14,
x_in_12_15,
x_in_12_2,
x_in_12_3,
x_in_12_4,
x_in_12_5,
x_in_12_6,
x_in_12_7,
x_in_12_8,
x_in_12_9,
x_in_13_0,
x_in_13_1,
x_in_13_10,
x_in_13_11,
x_in_13_12,
x_in_13_13,
x_in_13_14,
x_in_13_15,
x_in_13_2,
x_in_13_3,
x_in_13_4,
x_in_13_5,
x_in_13_6,
x_in_13_7,
x_in_13_8,
x_in_13_9,
x_in_14_0,
x_in_14_1,
x_in_14_10,
x_in_14_11,
x_in_14_12,
x_in_14_13,
x_in_14_14,
x_in_14_15,
x_in_14_2,
x_in_14_3,
x_in_14_4,
x_in_14_5,
x_in_14_6,
x_in_14_7,
x_in_14_8,
x_in_14_9,
x_in_15_0,
x_in_15_1,
x_in_15_10,
x_in_15_11,
x_in_15_12,
x_in_15_13,
x_in_15_14,
x_in_15_15,
x_in_15_2,
x_in_15_3,
x_in_15_4,
x_in_15_5,
x_in_15_6,
x_in_15_7,
x_in_15_8,
x_in_15_9,
x_in_16_0,
x_in_16_1,
x_in_16_10,
x_in_16_11,
x_in_16_12,
x_in_16_13,
x_in_16_14,
x_in_16_15,
x_in_16_2,
x_in_16_3,
x_in_16_4,
x_in_16_5,
x_in_16_6,
x_in_16_7,
x_in_16_8,
x_in_16_9,
x_in_17_0,
x_in_17_1,
x_in_17_10,
x_in_17_11,
x_in_17_12,
x_in_17_13,
x_in_17_14,
x_in_17_15,
x_in_17_2,
x_in_17_3,
x_in_17_4,
x_in_17_5,
x_in_17_6,
x_in_17_7,
x_in_17_8,
x_in_17_9,
x_in_18_0,
x_in_18_1,
x_in_18_10,
x_in_18_11,
x_in_18_12,
x_in_18_13,
x_in_18_14,
x_in_18_15,
x_in_18_2,
x_in_18_3,
x_in_18_4,
x_in_18_5,
x_in_18_6,
x_in_18_7,
x_in_18_8,
x_in_18_9,
x_in_19_0,
x_in_19_1,
x_in_19_10,
x_in_19_11,
x_in_19_12,
x_in_19_13,
x_in_19_14,
x_in_19_15,
x_in_19_2,
x_in_19_3,
x_in_19_4,
x_in_19_5,
x_in_19_6,
x_in_19_7,
x_in_19_8,
x_in_19_9,
x_in_1_0,
x_in_1_1,
x_in_1_10,
x_in_1_11,
x_in_1_12,
x_in_1_13,
x_in_1_14,
x_in_1_15,
x_in_1_2,
x_in_1_3,
x_in_1_4,
x_in_1_5,
x_in_1_6,
x_in_1_7,
x_in_1_8,
x_in_1_9,
x_in_20_0,
x_in_20_1,
x_in_20_10,
x_in_20_11,
x_in_20_12,
x_in_20_13,
x_in_20_14,
x_in_20_15,
x_in_20_2,
x_in_20_3,
x_in_20_4,
x_in_20_5,
x_in_20_6,
x_in_20_7,
x_in_20_8,
x_in_20_9,
x_in_21_0,
x_in_21_1,
x_in_21_10,
x_in_21_11,
x_in_21_12,
x_in_21_13,
x_in_21_14,
x_in_21_15,
x_in_21_2,
x_in_21_3,
x_in_21_4,
x_in_21_5,
x_in_21_6,
x_in_21_7,
x_in_21_8,
x_in_21_9,
x_in_22_0,
x_in_22_1,
x_in_22_10,
x_in_22_11,
x_in_22_12,
x_in_22_13,
x_in_22_14,
x_in_22_15,
x_in_22_2,
x_in_22_3,
x_in_22_4,
x_in_22_5,
x_in_22_6,
x_in_22_7,
x_in_22_8,
x_in_22_9,
x_in_23_0,
x_in_23_1,
x_in_23_10,
x_in_23_11,
x_in_23_12,
x_in_23_13,
x_in_23_14,
x_in_23_15,
x_in_23_2,
x_in_23_3,
x_in_23_4,
x_in_23_5,
x_in_23_6,
x_in_23_7,
x_in_23_8,
x_in_23_9,
x_in_24_0,
x_in_24_1,
x_in_24_10,
x_in_24_11,
x_in_24_12,
x_in_24_13,
x_in_24_14,
x_in_24_15,
x_in_24_2,
x_in_24_3,
x_in_24_4,
x_in_24_5,
x_in_24_6,
x_in_24_7,
x_in_24_8,
x_in_24_9,
x_in_25_0,
x_in_25_1,
x_in_25_10,
x_in_25_11,
x_in_25_12,
x_in_25_13,
x_in_25_14,
x_in_25_15,
x_in_25_2,
x_in_25_3,
x_in_25_4,
x_in_25_5,
x_in_25_6,
x_in_25_7,
x_in_25_8,
x_in_25_9,
x_in_26_0,
x_in_26_1,
x_in_26_10,
x_in_26_11,
x_in_26_12,
x_in_26_13,
x_in_26_14,
x_in_26_15,
x_in_26_2,
x_in_26_3,
x_in_26_4,
x_in_26_5,
x_in_26_6,
x_in_26_7,
x_in_26_8,
x_in_26_9,
x_in_27_0,
x_in_27_1,
x_in_27_10,
x_in_27_11,
x_in_27_12,
x_in_27_13,
x_in_27_14,
x_in_27_15,
x_in_27_2,
x_in_27_3,
x_in_27_4,
x_in_27_5,
x_in_27_6,
x_in_27_7,
x_in_27_8,
x_in_27_9,
x_in_28_0,
x_in_28_1,
x_in_28_10,
x_in_28_11,
x_in_28_12,
x_in_28_13,
x_in_28_14,
x_in_28_15,
x_in_28_2,
x_in_28_3,
x_in_28_4,
x_in_28_5,
x_in_28_6,
x_in_28_7,
x_in_28_8,
x_in_28_9,
x_in_29_0,
x_in_29_1,
x_in_29_10,
x_in_29_11,
x_in_29_12,
x_in_29_13,
x_in_29_14,
x_in_29_15,
x_in_29_2,
x_in_29_3,
x_in_29_4,
x_in_29_5,
x_in_29_6,
x_in_29_7,
x_in_29_8,
x_in_29_9,
x_in_2_0,
x_in_2_1,
x_in_2_10,
x_in_2_11,
x_in_2_12,
x_in_2_13,
x_in_2_14,
x_in_2_15,
x_in_2_2,
x_in_2_3,
x_in_2_4,
x_in_2_5,
x_in_2_6,
x_in_2_7,
x_in_2_8,
x_in_2_9,
x_in_30_0,
x_in_30_1,
x_in_30_10,
x_in_30_11,
x_in_30_12,
x_in_30_13,
x_in_30_14,
x_in_30_15,
x_in_30_2,
x_in_30_3,
x_in_30_4,
x_in_30_5,
x_in_30_6,
x_in_30_7,
x_in_30_8,
x_in_30_9,
x_in_31_0,
x_in_31_1,
x_in_31_10,
x_in_31_11,
x_in_31_12,
x_in_31_13,
x_in_31_14,
x_in_31_15,
x_in_31_2,
x_in_31_3,
x_in_31_4,
x_in_31_5,
x_in_31_6,
x_in_31_7,
x_in_31_8,
x_in_31_9,
x_in_32_0,
x_in_32_1,
x_in_32_10,
x_in_32_11,
x_in_32_12,
x_in_32_13,
x_in_32_14,
x_in_32_15,
x_in_32_2,
x_in_32_3,
x_in_32_4,
x_in_32_5,
x_in_32_6,
x_in_32_7,
x_in_32_8,
x_in_32_9,
x_in_33_0,
x_in_33_1,
x_in_33_10,
x_in_33_11,
x_in_33_12,
x_in_33_13,
x_in_33_14,
x_in_33_15,
x_in_33_2,
x_in_33_3,
x_in_33_4,
x_in_33_5,
x_in_33_6,
x_in_33_7,
x_in_33_8,
x_in_33_9,
x_in_34_0,
x_in_34_1,
x_in_34_10,
x_in_34_11,
x_in_34_12,
x_in_34_13,
x_in_34_14,
x_in_34_15,
x_in_34_2,
x_in_34_3,
x_in_34_4,
x_in_34_5,
x_in_34_6,
x_in_34_7,
x_in_34_8,
x_in_34_9,
x_in_35_0,
x_in_35_1,
x_in_35_10,
x_in_35_11,
x_in_35_12,
x_in_35_13,
x_in_35_14,
x_in_35_15,
x_in_35_2,
x_in_35_3,
x_in_35_4,
x_in_35_5,
x_in_35_6,
x_in_35_7,
x_in_35_8,
x_in_35_9,
x_in_36_0,
x_in_36_1,
x_in_36_10,
x_in_36_11,
x_in_36_12,
x_in_36_13,
x_in_36_14,
x_in_36_15,
x_in_36_2,
x_in_36_3,
x_in_36_4,
x_in_36_5,
x_in_36_6,
x_in_36_7,
x_in_36_8,
x_in_36_9,
x_in_37_0,
x_in_37_1,
x_in_37_10,
x_in_37_11,
x_in_37_12,
x_in_37_13,
x_in_37_14,
x_in_37_15,
x_in_37_2,
x_in_37_3,
x_in_37_4,
x_in_37_5,
x_in_37_6,
x_in_37_7,
x_in_37_8,
x_in_37_9,
x_in_38_0,
x_in_38_1,
x_in_38_10,
x_in_38_11,
x_in_38_12,
x_in_38_13,
x_in_38_14,
x_in_38_15,
x_in_38_2,
x_in_38_3,
x_in_38_4,
x_in_38_5,
x_in_38_6,
x_in_38_7,
x_in_38_8,
x_in_38_9,
x_in_39_0,
x_in_39_1,
x_in_39_10,
x_in_39_11,
x_in_39_12,
x_in_39_13,
x_in_39_14,
x_in_39_15,
x_in_39_2,
x_in_39_3,
x_in_39_4,
x_in_39_5,
x_in_39_6,
x_in_39_7,
x_in_39_8,
x_in_39_9,
x_in_3_0,
x_in_3_1,
x_in_3_10,
x_in_3_11,
x_in_3_12,
x_in_3_13,
x_in_3_14,
x_in_3_15,
x_in_3_2,
x_in_3_3,
x_in_3_4,
x_in_3_5,
x_in_3_6,
x_in_3_7,
x_in_3_8,
x_in_3_9,
x_in_40_0,
x_in_40_1,
x_in_40_10,
x_in_40_11,
x_in_40_12,
x_in_40_13,
x_in_40_14,
x_in_40_15,
x_in_40_2,
x_in_40_3,
x_in_40_4,
x_in_40_5,
x_in_40_6,
x_in_40_7,
x_in_40_8,
x_in_40_9,
x_in_41_0,
x_in_41_1,
x_in_41_10,
x_in_41_11,
x_in_41_12,
x_in_41_13,
x_in_41_14,
x_in_41_15,
x_in_41_2,
x_in_41_3,
x_in_41_4,
x_in_41_5,
x_in_41_6,
x_in_41_7,
x_in_41_8,
x_in_41_9,
x_in_42_0,
x_in_42_1,
x_in_42_10,
x_in_42_11,
x_in_42_12,
x_in_42_13,
x_in_42_14,
x_in_42_15,
x_in_42_2,
x_in_42_3,
x_in_42_4,
x_in_42_5,
x_in_42_6,
x_in_42_7,
x_in_42_8,
x_in_42_9,
x_in_43_0,
x_in_43_1,
x_in_43_10,
x_in_43_11,
x_in_43_12,
x_in_43_13,
x_in_43_14,
x_in_43_15,
x_in_43_2,
x_in_43_3,
x_in_43_4,
x_in_43_5,
x_in_43_6,
x_in_43_7,
x_in_43_8,
x_in_43_9,
x_in_44_0,
x_in_44_1,
x_in_44_10,
x_in_44_11,
x_in_44_12,
x_in_44_13,
x_in_44_14,
x_in_44_15,
x_in_44_2,
x_in_44_3,
x_in_44_4,
x_in_44_5,
x_in_44_6,
x_in_44_7,
x_in_44_8,
x_in_44_9,
x_in_45_0,
x_in_45_1,
x_in_45_10,
x_in_45_11,
x_in_45_12,
x_in_45_13,
x_in_45_14,
x_in_45_15,
x_in_45_2,
x_in_45_3,
x_in_45_4,
x_in_45_5,
x_in_45_6,
x_in_45_7,
x_in_45_8,
x_in_45_9,
x_in_46_0,
x_in_46_1,
x_in_46_10,
x_in_46_11,
x_in_46_12,
x_in_46_13,
x_in_46_14,
x_in_46_15,
x_in_46_2,
x_in_46_3,
x_in_46_4,
x_in_46_5,
x_in_46_6,
x_in_46_7,
x_in_46_8,
x_in_46_9,
x_in_47_0,
x_in_47_1,
x_in_47_10,
x_in_47_11,
x_in_47_12,
x_in_47_13,
x_in_47_14,
x_in_47_15,
x_in_47_2,
x_in_47_3,
x_in_47_4,
x_in_47_5,
x_in_47_6,
x_in_47_7,
x_in_47_8,
x_in_47_9,
x_in_48_0,
x_in_48_1,
x_in_48_10,
x_in_48_11,
x_in_48_12,
x_in_48_13,
x_in_48_14,
x_in_48_15,
x_in_48_2,
x_in_48_3,
x_in_48_4,
x_in_48_5,
x_in_48_6,
x_in_48_7,
x_in_48_8,
x_in_48_9,
x_in_49_0,
x_in_49_1,
x_in_49_10,
x_in_49_11,
x_in_49_12,
x_in_49_13,
x_in_49_14,
x_in_49_15,
x_in_49_2,
x_in_49_3,
x_in_49_4,
x_in_49_5,
x_in_49_6,
x_in_49_7,
x_in_49_8,
x_in_49_9,
x_in_4_0,
x_in_4_1,
x_in_4_10,
x_in_4_11,
x_in_4_12,
x_in_4_13,
x_in_4_14,
x_in_4_15,
x_in_4_2,
x_in_4_3,
x_in_4_4,
x_in_4_5,
x_in_4_6,
x_in_4_7,
x_in_4_8,
x_in_4_9,
x_in_50_0,
x_in_50_1,
x_in_50_10,
x_in_50_11,
x_in_50_12,
x_in_50_13,
x_in_50_14,
x_in_50_15,
x_in_50_2,
x_in_50_3,
x_in_50_4,
x_in_50_5,
x_in_50_6,
x_in_50_7,
x_in_50_8,
x_in_50_9,
x_in_51_0,
x_in_51_1,
x_in_51_10,
x_in_51_11,
x_in_51_12,
x_in_51_13,
x_in_51_14,
x_in_51_15,
x_in_51_2,
x_in_51_3,
x_in_51_4,
x_in_51_5,
x_in_51_6,
x_in_51_7,
x_in_51_8,
x_in_51_9,
x_in_52_0,
x_in_52_1,
x_in_52_10,
x_in_52_11,
x_in_52_12,
x_in_52_13,
x_in_52_14,
x_in_52_15,
x_in_52_2,
x_in_52_3,
x_in_52_4,
x_in_52_5,
x_in_52_6,
x_in_52_7,
x_in_52_8,
x_in_52_9,
x_in_53_0,
x_in_53_1,
x_in_53_10,
x_in_53_11,
x_in_53_12,
x_in_53_13,
x_in_53_14,
x_in_53_15,
x_in_53_2,
x_in_53_3,
x_in_53_4,
x_in_53_5,
x_in_53_6,
x_in_53_7,
x_in_53_8,
x_in_53_9,
x_in_54_0,
x_in_54_1,
x_in_54_10,
x_in_54_11,
x_in_54_12,
x_in_54_13,
x_in_54_14,
x_in_54_15,
x_in_54_2,
x_in_54_3,
x_in_54_4,
x_in_54_5,
x_in_54_6,
x_in_54_7,
x_in_54_8,
x_in_54_9,
x_in_55_0,
x_in_55_1,
x_in_55_10,
x_in_55_11,
x_in_55_12,
x_in_55_13,
x_in_55_14,
x_in_55_15,
x_in_55_2,
x_in_55_3,
x_in_55_4,
x_in_55_5,
x_in_55_6,
x_in_55_7,
x_in_55_8,
x_in_55_9,
x_in_56_0,
x_in_56_1,
x_in_56_10,
x_in_56_11,
x_in_56_12,
x_in_56_13,
x_in_56_14,
x_in_56_15,
x_in_56_2,
x_in_56_3,
x_in_56_4,
x_in_56_5,
x_in_56_6,
x_in_56_7,
x_in_56_8,
x_in_56_9,
x_in_57_0,
x_in_57_1,
x_in_57_10,
x_in_57_11,
x_in_57_12,
x_in_57_13,
x_in_57_14,
x_in_57_15,
x_in_57_2,
x_in_57_3,
x_in_57_4,
x_in_57_5,
x_in_57_6,
x_in_57_7,
x_in_57_8,
x_in_57_9,
x_in_58_0,
x_in_58_1,
x_in_58_10,
x_in_58_11,
x_in_58_12,
x_in_58_13,
x_in_58_14,
x_in_58_15,
x_in_58_2,
x_in_58_3,
x_in_58_4,
x_in_58_5,
x_in_58_6,
x_in_58_7,
x_in_58_8,
x_in_58_9,
x_in_59_0,
x_in_59_1,
x_in_59_10,
x_in_59_11,
x_in_59_12,
x_in_59_13,
x_in_59_14,
x_in_59_15,
x_in_59_2,
x_in_59_3,
x_in_59_4,
x_in_59_5,
x_in_59_6,
x_in_59_7,
x_in_59_8,
x_in_59_9,
x_in_5_0,
x_in_5_1,
x_in_5_10,
x_in_5_11,
x_in_5_12,
x_in_5_13,
x_in_5_14,
x_in_5_15,
x_in_5_2,
x_in_5_3,
x_in_5_4,
x_in_5_5,
x_in_5_6,
x_in_5_7,
x_in_5_8,
x_in_5_9,
x_in_60_0,
x_in_60_1,
x_in_60_10,
x_in_60_11,
x_in_60_12,
x_in_60_13,
x_in_60_14,
x_in_60_15,
x_in_60_2,
x_in_60_3,
x_in_60_4,
x_in_60_5,
x_in_60_6,
x_in_60_7,
x_in_60_8,
x_in_60_9,
x_in_61_0,
x_in_61_1,
x_in_61_10,
x_in_61_11,
x_in_61_12,
x_in_61_13,
x_in_61_14,
x_in_61_15,
x_in_61_2,
x_in_61_3,
x_in_61_4,
x_in_61_5,
x_in_61_6,
x_in_61_7,
x_in_61_8,
x_in_61_9,
x_in_62_0,
x_in_62_1,
x_in_62_10,
x_in_62_11,
x_in_62_12,
x_in_62_13,
x_in_62_14,
x_in_62_15,
x_in_62_2,
x_in_62_3,
x_in_62_4,
x_in_62_5,
x_in_62_6,
x_in_62_7,
x_in_62_8,
x_in_62_9,
x_in_63_0,
x_in_63_1,
x_in_63_10,
x_in_63_11,
x_in_63_12,
x_in_63_13,
x_in_63_14,
x_in_63_15,
x_in_63_2,
x_in_63_3,
x_in_63_4,
x_in_63_5,
x_in_63_6,
x_in_63_7,
x_in_63_8,
x_in_63_9,
x_in_6_0,
x_in_6_1,
x_in_6_10,
x_in_6_11,
x_in_6_12,
x_in_6_13,
x_in_6_14,
x_in_6_15,
x_in_6_2,
x_in_6_3,
x_in_6_4,
x_in_6_5,
x_in_6_6,
x_in_6_7,
x_in_6_8,
x_in_6_9,
x_in_7_0,
x_in_7_1,
x_in_7_10,
x_in_7_11,
x_in_7_12,
x_in_7_13,
x_in_7_14,
x_in_7_15,
x_in_7_2,
x_in_7_3,
x_in_7_4,
x_in_7_5,
x_in_7_6,
x_in_7_7,
x_in_7_8,
x_in_7_9,
x_in_8_0,
x_in_8_1,
x_in_8_10,
x_in_8_11,
x_in_8_12,
x_in_8_13,
x_in_8_14,
x_in_8_15,
x_in_8_2,
x_in_8_3,
x_in_8_4,
x_in_8_5,
x_in_8_6,
x_in_8_7,
x_in_8_8,
x_in_8_9,
x_in_9_0,
x_in_9_1,
x_in_9_10,
x_in_9_11,
x_in_9_12,
x_in_9_13,
x_in_9_14,
x_in_9_15,
x_in_9_2,
x_in_9_3,
x_in_9_4,
x_in_9_5,
x_in_9_6,
x_in_9_7,
x_in_9_8,
x_in_9_9,
x_out_0_0,
x_out_0_1,
x_out_0_10,
x_out_0_11,
x_out_0_12,
x_out_0_13,
x_out_0_14,
x_out_0_15,
x_out_0_2,
x_out_0_3,
x_out_0_4,
x_out_0_5,
x_out_0_6,
x_out_0_7,
x_out_0_8,
x_out_0_9,
x_out_10_0,
x_out_10_1,
x_out_10_10,
x_out_10_11,
x_out_10_12,
x_out_10_13,
x_out_10_14,
x_out_10_15,
x_out_10_18,
x_out_10_19,
x_out_10_2,
x_out_10_20,
x_out_10_21,
x_out_10_22,
x_out_10_23,
x_out_10_24,
x_out_10_25,
x_out_10_26,
x_out_10_27,
x_out_10_28,
x_out_10_29,
x_out_10_3,
x_out_10_30,
x_out_10_31,
x_out_10_32,
x_out_10_33,
x_out_10_4,
x_out_10_5,
x_out_10_6,
x_out_10_7,
x_out_10_8,
x_out_10_9,
x_out_11_0,
x_out_11_1,
x_out_11_10,
x_out_11_11,
x_out_11_12,
x_out_11_13,
x_out_11_14,
x_out_11_15,
x_out_11_18,
x_out_11_19,
x_out_11_2,
x_out_11_20,
x_out_11_21,
x_out_11_22,
x_out_11_23,
x_out_11_24,
x_out_11_25,
x_out_11_26,
x_out_11_27,
x_out_11_28,
x_out_11_29,
x_out_11_3,
x_out_11_30,
x_out_11_31,
x_out_11_32,
x_out_11_33,
x_out_11_4,
x_out_11_5,
x_out_11_6,
x_out_11_7,
x_out_11_8,
x_out_11_9,
x_out_12_0,
x_out_12_1,
x_out_12_10,
x_out_12_11,
x_out_12_12,
x_out_12_13,
x_out_12_14,
x_out_12_15,
x_out_12_18,
x_out_12_19,
x_out_12_2,
x_out_12_20,
x_out_12_21,
x_out_12_22,
x_out_12_23,
x_out_12_24,
x_out_12_25,
x_out_12_26,
x_out_12_27,
x_out_12_28,
x_out_12_29,
x_out_12_3,
x_out_12_30,
x_out_12_31,
x_out_12_32,
x_out_12_33,
x_out_12_4,
x_out_12_5,
x_out_12_6,
x_out_12_7,
x_out_12_8,
x_out_12_9,
x_out_13_0,
x_out_13_1,
x_out_13_10,
x_out_13_11,
x_out_13_12,
x_out_13_13,
x_out_13_14,
x_out_13_15,
x_out_13_18,
x_out_13_19,
x_out_13_2,
x_out_13_20,
x_out_13_21,
x_out_13_22,
x_out_13_23,
x_out_13_24,
x_out_13_25,
x_out_13_26,
x_out_13_27,
x_out_13_28,
x_out_13_29,
x_out_13_3,
x_out_13_30,
x_out_13_31,
x_out_13_32,
x_out_13_33,
x_out_13_4,
x_out_13_5,
x_out_13_6,
x_out_13_7,
x_out_13_8,
x_out_13_9,
x_out_14_0,
x_out_14_1,
x_out_14_10,
x_out_14_11,
x_out_14_12,
x_out_14_13,
x_out_14_14,
x_out_14_15,
x_out_14_18,
x_out_14_19,
x_out_14_2,
x_out_14_20,
x_out_14_21,
x_out_14_22,
x_out_14_23,
x_out_14_24,
x_out_14_25,
x_out_14_26,
x_out_14_27,
x_out_14_28,
x_out_14_29,
x_out_14_3,
x_out_14_30,
x_out_14_31,
x_out_14_32,
x_out_14_33,
x_out_14_4,
x_out_14_5,
x_out_14_6,
x_out_14_7,
x_out_14_8,
x_out_14_9,
x_out_15_0,
x_out_15_1,
x_out_15_10,
x_out_15_11,
x_out_15_12,
x_out_15_13,
x_out_15_14,
x_out_15_15,
x_out_15_18,
x_out_15_19,
x_out_15_2,
x_out_15_20,
x_out_15_21,
x_out_15_22,
x_out_15_23,
x_out_15_24,
x_out_15_25,
x_out_15_26,
x_out_15_27,
x_out_15_28,
x_out_15_29,
x_out_15_3,
x_out_15_30,
x_out_15_31,
x_out_15_32,
x_out_15_33,
x_out_15_4,
x_out_15_5,
x_out_15_6,
x_out_15_7,
x_out_15_8,
x_out_15_9,
x_out_16_0,
x_out_16_1,
x_out_16_10,
x_out_16_11,
x_out_16_12,
x_out_16_13,
x_out_16_14,
x_out_16_15,
x_out_16_18,
x_out_16_19,
x_out_16_2,
x_out_16_20,
x_out_16_21,
x_out_16_22,
x_out_16_23,
x_out_16_24,
x_out_16_25,
x_out_16_26,
x_out_16_27,
x_out_16_28,
x_out_16_29,
x_out_16_3,
x_out_16_30,
x_out_16_31,
x_out_16_32,
x_out_16_33,
x_out_16_4,
x_out_16_5,
x_out_16_6,
x_out_16_7,
x_out_16_8,
x_out_16_9,
x_out_17_0,
x_out_17_1,
x_out_17_10,
x_out_17_11,
x_out_17_12,
x_out_17_13,
x_out_17_14,
x_out_17_15,
x_out_17_18,
x_out_17_19,
x_out_17_2,
x_out_17_20,
x_out_17_21,
x_out_17_22,
x_out_17_23,
x_out_17_24,
x_out_17_25,
x_out_17_26,
x_out_17_27,
x_out_17_28,
x_out_17_29,
x_out_17_3,
x_out_17_30,
x_out_17_31,
x_out_17_32,
x_out_17_33,
x_out_17_4,
x_out_17_5,
x_out_17_6,
x_out_17_7,
x_out_17_8,
x_out_17_9,
x_out_18_0,
x_out_18_1,
x_out_18_10,
x_out_18_11,
x_out_18_12,
x_out_18_13,
x_out_18_14,
x_out_18_15,
x_out_18_18,
x_out_18_19,
x_out_18_2,
x_out_18_20,
x_out_18_21,
x_out_18_22,
x_out_18_23,
x_out_18_24,
x_out_18_25,
x_out_18_26,
x_out_18_27,
x_out_18_28,
x_out_18_29,
x_out_18_3,
x_out_18_30,
x_out_18_31,
x_out_18_32,
x_out_18_33,
x_out_18_4,
x_out_18_5,
x_out_18_6,
x_out_18_7,
x_out_18_8,
x_out_18_9,
x_out_19_0,
x_out_19_1,
x_out_19_10,
x_out_19_11,
x_out_19_12,
x_out_19_13,
x_out_19_14,
x_out_19_15,
x_out_19_18,
x_out_19_19,
x_out_19_2,
x_out_19_20,
x_out_19_21,
x_out_19_22,
x_out_19_23,
x_out_19_24,
x_out_19_25,
x_out_19_26,
x_out_19_27,
x_out_19_28,
x_out_19_29,
x_out_19_3,
x_out_19_30,
x_out_19_31,
x_out_19_32,
x_out_19_33,
x_out_19_4,
x_out_19_5,
x_out_19_6,
x_out_19_7,
x_out_19_8,
x_out_19_9,
x_out_1_0,
x_out_1_1,
x_out_1_10,
x_out_1_11,
x_out_1_12,
x_out_1_13,
x_out_1_14,
x_out_1_15,
x_out_1_18,
x_out_1_19,
x_out_1_2,
x_out_1_20,
x_out_1_21,
x_out_1_22,
x_out_1_23,
x_out_1_24,
x_out_1_25,
x_out_1_26,
x_out_1_27,
x_out_1_28,
x_out_1_29,
x_out_1_3,
x_out_1_30,
x_out_1_31,
x_out_1_32,
x_out_1_33,
x_out_1_4,
x_out_1_5,
x_out_1_6,
x_out_1_7,
x_out_1_8,
x_out_1_9,
x_out_20_0,
x_out_20_1,
x_out_20_10,
x_out_20_11,
x_out_20_12,
x_out_20_13,
x_out_20_14,
x_out_20_15,
x_out_20_2,
x_out_20_3,
x_out_20_4,
x_out_20_5,
x_out_20_6,
x_out_20_7,
x_out_20_8,
x_out_20_9,
x_out_21_0,
x_out_21_1,
x_out_21_10,
x_out_21_11,
x_out_21_12,
x_out_21_13,
x_out_21_14,
x_out_21_15,
x_out_21_18,
x_out_21_19,
x_out_21_2,
x_out_21_20,
x_out_21_21,
x_out_21_22,
x_out_21_23,
x_out_21_24,
x_out_21_25,
x_out_21_26,
x_out_21_27,
x_out_21_28,
x_out_21_29,
x_out_21_3,
x_out_21_30,
x_out_21_31,
x_out_21_32,
x_out_21_33,
x_out_21_4,
x_out_21_5,
x_out_21_6,
x_out_21_7,
x_out_21_8,
x_out_21_9,
x_out_22_0,
x_out_22_1,
x_out_22_10,
x_out_22_11,
x_out_22_12,
x_out_22_13,
x_out_22_14,
x_out_22_15,
x_out_22_18,
x_out_22_19,
x_out_22_2,
x_out_22_20,
x_out_22_21,
x_out_22_22,
x_out_22_23,
x_out_22_24,
x_out_22_25,
x_out_22_26,
x_out_22_27,
x_out_22_28,
x_out_22_29,
x_out_22_3,
x_out_22_30,
x_out_22_31,
x_out_22_32,
x_out_22_33,
x_out_22_4,
x_out_22_5,
x_out_22_6,
x_out_22_7,
x_out_22_8,
x_out_22_9,
x_out_23_0,
x_out_23_1,
x_out_23_10,
x_out_23_11,
x_out_23_12,
x_out_23_13,
x_out_23_14,
x_out_23_15,
x_out_23_18,
x_out_23_19,
x_out_23_2,
x_out_23_20,
x_out_23_21,
x_out_23_22,
x_out_23_23,
x_out_23_24,
x_out_23_25,
x_out_23_26,
x_out_23_27,
x_out_23_28,
x_out_23_29,
x_out_23_3,
x_out_23_30,
x_out_23_31,
x_out_23_32,
x_out_23_33,
x_out_23_4,
x_out_23_5,
x_out_23_6,
x_out_23_7,
x_out_23_8,
x_out_23_9,
x_out_24_0,
x_out_24_1,
x_out_24_10,
x_out_24_11,
x_out_24_12,
x_out_24_13,
x_out_24_14,
x_out_24_15,
x_out_24_18,
x_out_24_19,
x_out_24_2,
x_out_24_20,
x_out_24_21,
x_out_24_22,
x_out_24_23,
x_out_24_24,
x_out_24_25,
x_out_24_26,
x_out_24_27,
x_out_24_28,
x_out_24_29,
x_out_24_3,
x_out_24_30,
x_out_24_31,
x_out_24_32,
x_out_24_33,
x_out_24_4,
x_out_24_5,
x_out_24_6,
x_out_24_7,
x_out_24_8,
x_out_24_9,
x_out_25_0,
x_out_25_1,
x_out_25_10,
x_out_25_11,
x_out_25_12,
x_out_25_13,
x_out_25_14,
x_out_25_15,
x_out_25_18,
x_out_25_19,
x_out_25_2,
x_out_25_20,
x_out_25_21,
x_out_25_22,
x_out_25_23,
x_out_25_24,
x_out_25_25,
x_out_25_26,
x_out_25_27,
x_out_25_28,
x_out_25_29,
x_out_25_3,
x_out_25_30,
x_out_25_31,
x_out_25_32,
x_out_25_33,
x_out_25_4,
x_out_25_5,
x_out_25_6,
x_out_25_7,
x_out_25_8,
x_out_25_9,
x_out_26_0,
x_out_26_1,
x_out_26_10,
x_out_26_11,
x_out_26_12,
x_out_26_13,
x_out_26_14,
x_out_26_15,
x_out_26_18,
x_out_26_19,
x_out_26_2,
x_out_26_20,
x_out_26_21,
x_out_26_22,
x_out_26_23,
x_out_26_24,
x_out_26_25,
x_out_26_26,
x_out_26_27,
x_out_26_28,
x_out_26_29,
x_out_26_3,
x_out_26_30,
x_out_26_31,
x_out_26_32,
x_out_26_33,
x_out_26_4,
x_out_26_5,
x_out_26_6,
x_out_26_7,
x_out_26_8,
x_out_26_9,
x_out_27_0,
x_out_27_1,
x_out_27_10,
x_out_27_11,
x_out_27_12,
x_out_27_13,
x_out_27_14,
x_out_27_15,
x_out_27_18,
x_out_27_19,
x_out_27_2,
x_out_27_20,
x_out_27_21,
x_out_27_22,
x_out_27_23,
x_out_27_24,
x_out_27_25,
x_out_27_26,
x_out_27_27,
x_out_27_28,
x_out_27_29,
x_out_27_3,
x_out_27_30,
x_out_27_31,
x_out_27_32,
x_out_27_33,
x_out_27_4,
x_out_27_5,
x_out_27_6,
x_out_27_7,
x_out_27_8,
x_out_27_9,
x_out_28_0,
x_out_28_1,
x_out_28_10,
x_out_28_11,
x_out_28_12,
x_out_28_13,
x_out_28_14,
x_out_28_15,
x_out_28_18,
x_out_28_19,
x_out_28_2,
x_out_28_20,
x_out_28_21,
x_out_28_22,
x_out_28_23,
x_out_28_24,
x_out_28_25,
x_out_28_26,
x_out_28_27,
x_out_28_28,
x_out_28_29,
x_out_28_3,
x_out_28_30,
x_out_28_31,
x_out_28_32,
x_out_28_33,
x_out_28_4,
x_out_28_5,
x_out_28_6,
x_out_28_7,
x_out_28_8,
x_out_28_9,
x_out_29_0,
x_out_29_1,
x_out_29_10,
x_out_29_11,
x_out_29_12,
x_out_29_13,
x_out_29_14,
x_out_29_15,
x_out_29_18,
x_out_29_19,
x_out_29_2,
x_out_29_20,
x_out_29_21,
x_out_29_22,
x_out_29_23,
x_out_29_24,
x_out_29_25,
x_out_29_26,
x_out_29_27,
x_out_29_28,
x_out_29_29,
x_out_29_3,
x_out_29_30,
x_out_29_31,
x_out_29_32,
x_out_29_33,
x_out_29_4,
x_out_29_5,
x_out_29_6,
x_out_29_7,
x_out_29_8,
x_out_29_9,
x_out_2_0,
x_out_2_1,
x_out_2_10,
x_out_2_11,
x_out_2_12,
x_out_2_13,
x_out_2_14,
x_out_2_15,
x_out_2_18,
x_out_2_19,
x_out_2_2,
x_out_2_20,
x_out_2_21,
x_out_2_22,
x_out_2_23,
x_out_2_24,
x_out_2_25,
x_out_2_26,
x_out_2_27,
x_out_2_28,
x_out_2_29,
x_out_2_3,
x_out_2_30,
x_out_2_31,
x_out_2_32,
x_out_2_33,
x_out_2_4,
x_out_2_5,
x_out_2_6,
x_out_2_7,
x_out_2_8,
x_out_2_9,
x_out_30_0,
x_out_30_1,
x_out_30_10,
x_out_30_11,
x_out_30_12,
x_out_30_13,
x_out_30_14,
x_out_30_15,
x_out_30_18,
x_out_30_19,
x_out_30_2,
x_out_30_20,
x_out_30_21,
x_out_30_22,
x_out_30_23,
x_out_30_24,
x_out_30_25,
x_out_30_26,
x_out_30_27,
x_out_30_28,
x_out_30_29,
x_out_30_3,
x_out_30_30,
x_out_30_31,
x_out_30_32,
x_out_30_33,
x_out_30_4,
x_out_30_5,
x_out_30_6,
x_out_30_7,
x_out_30_8,
x_out_30_9,
x_out_31_0,
x_out_31_1,
x_out_31_10,
x_out_31_11,
x_out_31_12,
x_out_31_13,
x_out_31_14,
x_out_31_15,
x_out_31_18,
x_out_31_19,
x_out_31_2,
x_out_31_20,
x_out_31_21,
x_out_31_22,
x_out_31_23,
x_out_31_24,
x_out_31_25,
x_out_31_26,
x_out_31_27,
x_out_31_28,
x_out_31_29,
x_out_31_3,
x_out_31_30,
x_out_31_31,
x_out_31_32,
x_out_31_33,
x_out_31_4,
x_out_31_5,
x_out_31_6,
x_out_31_7,
x_out_31_8,
x_out_31_9,
x_out_32_0,
x_out_32_1,
x_out_32_10,
x_out_32_11,
x_out_32_12,
x_out_32_13,
x_out_32_14,
x_out_32_15,
x_out_32_2,
x_out_32_3,
x_out_32_4,
x_out_32_5,
x_out_32_6,
x_out_32_7,
x_out_32_8,
x_out_32_9,
x_out_33_0,
x_out_33_1,
x_out_33_10,
x_out_33_11,
x_out_33_12,
x_out_33_13,
x_out_33_14,
x_out_33_15,
x_out_33_18,
x_out_33_19,
x_out_33_2,
x_out_33_20,
x_out_33_21,
x_out_33_22,
x_out_33_23,
x_out_33_24,
x_out_33_25,
x_out_33_26,
x_out_33_27,
x_out_33_28,
x_out_33_29,
x_out_33_3,
x_out_33_30,
x_out_33_31,
x_out_33_32,
x_out_33_33,
x_out_33_4,
x_out_33_5,
x_out_33_6,
x_out_33_7,
x_out_33_8,
x_out_33_9,
x_out_34_0,
x_out_34_1,
x_out_34_10,
x_out_34_11,
x_out_34_12,
x_out_34_13,
x_out_34_14,
x_out_34_15,
x_out_34_18,
x_out_34_19,
x_out_34_2,
x_out_34_20,
x_out_34_21,
x_out_34_22,
x_out_34_23,
x_out_34_24,
x_out_34_25,
x_out_34_26,
x_out_34_27,
x_out_34_28,
x_out_34_29,
x_out_34_3,
x_out_34_30,
x_out_34_31,
x_out_34_32,
x_out_34_33,
x_out_34_4,
x_out_34_5,
x_out_34_6,
x_out_34_7,
x_out_34_8,
x_out_34_9,
x_out_35_0,
x_out_35_1,
x_out_35_10,
x_out_35_11,
x_out_35_12,
x_out_35_13,
x_out_35_14,
x_out_35_15,
x_out_35_18,
x_out_35_19,
x_out_35_2,
x_out_35_20,
x_out_35_21,
x_out_35_22,
x_out_35_23,
x_out_35_24,
x_out_35_25,
x_out_35_26,
x_out_35_27,
x_out_35_28,
x_out_35_29,
x_out_35_3,
x_out_35_30,
x_out_35_31,
x_out_35_32,
x_out_35_33,
x_out_35_4,
x_out_35_5,
x_out_35_6,
x_out_35_7,
x_out_35_8,
x_out_35_9,
x_out_36_0,
x_out_36_1,
x_out_36_10,
x_out_36_11,
x_out_36_12,
x_out_36_13,
x_out_36_14,
x_out_36_15,
x_out_36_18,
x_out_36_19,
x_out_36_2,
x_out_36_20,
x_out_36_21,
x_out_36_22,
x_out_36_23,
x_out_36_24,
x_out_36_25,
x_out_36_26,
x_out_36_27,
x_out_36_28,
x_out_36_29,
x_out_36_3,
x_out_36_30,
x_out_36_31,
x_out_36_32,
x_out_36_33,
x_out_36_4,
x_out_36_5,
x_out_36_6,
x_out_36_7,
x_out_36_8,
x_out_36_9,
x_out_37_0,
x_out_37_1,
x_out_37_10,
x_out_37_11,
x_out_37_12,
x_out_37_13,
x_out_37_14,
x_out_37_15,
x_out_37_18,
x_out_37_19,
x_out_37_2,
x_out_37_20,
x_out_37_21,
x_out_37_22,
x_out_37_23,
x_out_37_24,
x_out_37_25,
x_out_37_26,
x_out_37_27,
x_out_37_28,
x_out_37_29,
x_out_37_3,
x_out_37_30,
x_out_37_31,
x_out_37_32,
x_out_37_33,
x_out_37_4,
x_out_37_5,
x_out_37_6,
x_out_37_7,
x_out_37_8,
x_out_37_9,
x_out_38_0,
x_out_38_1,
x_out_38_10,
x_out_38_11,
x_out_38_12,
x_out_38_13,
x_out_38_14,
x_out_38_15,
x_out_38_18,
x_out_38_19,
x_out_38_2,
x_out_38_20,
x_out_38_21,
x_out_38_22,
x_out_38_23,
x_out_38_24,
x_out_38_25,
x_out_38_26,
x_out_38_27,
x_out_38_28,
x_out_38_29,
x_out_38_3,
x_out_38_30,
x_out_38_31,
x_out_38_32,
x_out_38_33,
x_out_38_4,
x_out_38_5,
x_out_38_6,
x_out_38_7,
x_out_38_8,
x_out_38_9,
x_out_39_0,
x_out_39_1,
x_out_39_10,
x_out_39_11,
x_out_39_12,
x_out_39_13,
x_out_39_14,
x_out_39_15,
x_out_39_18,
x_out_39_19,
x_out_39_2,
x_out_39_20,
x_out_39_21,
x_out_39_22,
x_out_39_23,
x_out_39_24,
x_out_39_25,
x_out_39_26,
x_out_39_27,
x_out_39_28,
x_out_39_29,
x_out_39_3,
x_out_39_30,
x_out_39_31,
x_out_39_32,
x_out_39_33,
x_out_39_4,
x_out_39_5,
x_out_39_6,
x_out_39_7,
x_out_39_8,
x_out_39_9,
x_out_3_0,
x_out_3_1,
x_out_3_10,
x_out_3_11,
x_out_3_12,
x_out_3_13,
x_out_3_14,
x_out_3_15,
x_out_3_18,
x_out_3_19,
x_out_3_2,
x_out_3_20,
x_out_3_21,
x_out_3_22,
x_out_3_23,
x_out_3_24,
x_out_3_25,
x_out_3_26,
x_out_3_27,
x_out_3_28,
x_out_3_29,
x_out_3_3,
x_out_3_30,
x_out_3_31,
x_out_3_32,
x_out_3_33,
x_out_3_4,
x_out_3_5,
x_out_3_6,
x_out_3_7,
x_out_3_8,
x_out_3_9,
x_out_40_0,
x_out_40_1,
x_out_40_10,
x_out_40_11,
x_out_40_12,
x_out_40_13,
x_out_40_14,
x_out_40_15,
x_out_40_18,
x_out_40_19,
x_out_40_2,
x_out_40_20,
x_out_40_21,
x_out_40_22,
x_out_40_23,
x_out_40_24,
x_out_40_25,
x_out_40_26,
x_out_40_27,
x_out_40_28,
x_out_40_29,
x_out_40_3,
x_out_40_30,
x_out_40_31,
x_out_40_32,
x_out_40_33,
x_out_40_4,
x_out_40_5,
x_out_40_6,
x_out_40_7,
x_out_40_8,
x_out_40_9,
x_out_41_0,
x_out_41_1,
x_out_41_10,
x_out_41_11,
x_out_41_12,
x_out_41_13,
x_out_41_14,
x_out_41_15,
x_out_41_18,
x_out_41_19,
x_out_41_2,
x_out_41_20,
x_out_41_21,
x_out_41_22,
x_out_41_23,
x_out_41_24,
x_out_41_25,
x_out_41_26,
x_out_41_27,
x_out_41_28,
x_out_41_29,
x_out_41_3,
x_out_41_30,
x_out_41_31,
x_out_41_32,
x_out_41_33,
x_out_41_4,
x_out_41_5,
x_out_41_6,
x_out_41_7,
x_out_41_8,
x_out_41_9,
x_out_42_0,
x_out_42_1,
x_out_42_10,
x_out_42_11,
x_out_42_12,
x_out_42_13,
x_out_42_14,
x_out_42_15,
x_out_42_18,
x_out_42_19,
x_out_42_2,
x_out_42_20,
x_out_42_21,
x_out_42_22,
x_out_42_23,
x_out_42_24,
x_out_42_25,
x_out_42_26,
x_out_42_27,
x_out_42_28,
x_out_42_29,
x_out_42_3,
x_out_42_30,
x_out_42_31,
x_out_42_32,
x_out_42_33,
x_out_42_4,
x_out_42_5,
x_out_42_6,
x_out_42_7,
x_out_42_8,
x_out_42_9,
x_out_43_0,
x_out_43_1,
x_out_43_10,
x_out_43_11,
x_out_43_12,
x_out_43_13,
x_out_43_14,
x_out_43_15,
x_out_43_18,
x_out_43_19,
x_out_43_2,
x_out_43_20,
x_out_43_21,
x_out_43_22,
x_out_43_23,
x_out_43_24,
x_out_43_25,
x_out_43_26,
x_out_43_27,
x_out_43_28,
x_out_43_29,
x_out_43_3,
x_out_43_30,
x_out_43_31,
x_out_43_32,
x_out_43_33,
x_out_43_4,
x_out_43_5,
x_out_43_6,
x_out_43_7,
x_out_43_8,
x_out_43_9,
x_out_44_0,
x_out_44_1,
x_out_44_10,
x_out_44_11,
x_out_44_12,
x_out_44_13,
x_out_44_14,
x_out_44_15,
x_out_44_18,
x_out_44_19,
x_out_44_2,
x_out_44_20,
x_out_44_21,
x_out_44_22,
x_out_44_23,
x_out_44_24,
x_out_44_25,
x_out_44_26,
x_out_44_27,
x_out_44_28,
x_out_44_29,
x_out_44_3,
x_out_44_30,
x_out_44_31,
x_out_44_32,
x_out_44_33,
x_out_44_4,
x_out_44_5,
x_out_44_6,
x_out_44_7,
x_out_44_8,
x_out_44_9,
x_out_45_0,
x_out_45_1,
x_out_45_10,
x_out_45_11,
x_out_45_12,
x_out_45_13,
x_out_45_14,
x_out_45_15,
x_out_45_18,
x_out_45_19,
x_out_45_2,
x_out_45_20,
x_out_45_21,
x_out_45_22,
x_out_45_23,
x_out_45_24,
x_out_45_25,
x_out_45_26,
x_out_45_27,
x_out_45_28,
x_out_45_29,
x_out_45_3,
x_out_45_30,
x_out_45_31,
x_out_45_32,
x_out_45_33,
x_out_45_4,
x_out_45_5,
x_out_45_6,
x_out_45_7,
x_out_45_8,
x_out_45_9,
x_out_46_0,
x_out_46_1,
x_out_46_10,
x_out_46_11,
x_out_46_12,
x_out_46_13,
x_out_46_14,
x_out_46_15,
x_out_46_18,
x_out_46_19,
x_out_46_2,
x_out_46_20,
x_out_46_21,
x_out_46_22,
x_out_46_23,
x_out_46_24,
x_out_46_25,
x_out_46_26,
x_out_46_27,
x_out_46_28,
x_out_46_29,
x_out_46_3,
x_out_46_30,
x_out_46_31,
x_out_46_32,
x_out_46_33,
x_out_46_4,
x_out_46_5,
x_out_46_6,
x_out_46_7,
x_out_46_8,
x_out_46_9,
x_out_47_0,
x_out_47_1,
x_out_47_10,
x_out_47_11,
x_out_47_12,
x_out_47_13,
x_out_47_14,
x_out_47_15,
x_out_47_18,
x_out_47_19,
x_out_47_2,
x_out_47_20,
x_out_47_21,
x_out_47_22,
x_out_47_23,
x_out_47_24,
x_out_47_25,
x_out_47_26,
x_out_47_27,
x_out_47_28,
x_out_47_29,
x_out_47_3,
x_out_47_30,
x_out_47_31,
x_out_47_32,
x_out_47_33,
x_out_47_4,
x_out_47_5,
x_out_47_6,
x_out_47_7,
x_out_47_8,
x_out_47_9,
x_out_48_0,
x_out_48_1,
x_out_48_10,
x_out_48_11,
x_out_48_12,
x_out_48_13,
x_out_48_14,
x_out_48_15,
x_out_48_18,
x_out_48_19,
x_out_48_2,
x_out_48_20,
x_out_48_21,
x_out_48_22,
x_out_48_23,
x_out_48_24,
x_out_48_25,
x_out_48_26,
x_out_48_27,
x_out_48_28,
x_out_48_29,
x_out_48_3,
x_out_48_30,
x_out_48_31,
x_out_48_32,
x_out_48_33,
x_out_48_4,
x_out_48_5,
x_out_48_6,
x_out_48_7,
x_out_48_8,
x_out_48_9,
x_out_49_0,
x_out_49_1,
x_out_49_10,
x_out_49_11,
x_out_49_12,
x_out_49_13,
x_out_49_14,
x_out_49_15,
x_out_49_18,
x_out_49_19,
x_out_49_2,
x_out_49_20,
x_out_49_21,
x_out_49_22,
x_out_49_23,
x_out_49_24,
x_out_49_25,
x_out_49_26,
x_out_49_27,
x_out_49_28,
x_out_49_29,
x_out_49_3,
x_out_49_30,
x_out_49_31,
x_out_49_32,
x_out_49_33,
x_out_49_4,
x_out_49_5,
x_out_49_6,
x_out_49_7,
x_out_49_8,
x_out_49_9,
x_out_4_0,
x_out_4_1,
x_out_4_10,
x_out_4_11,
x_out_4_12,
x_out_4_13,
x_out_4_14,
x_out_4_15,
x_out_4_18,
x_out_4_19,
x_out_4_2,
x_out_4_20,
x_out_4_21,
x_out_4_22,
x_out_4_23,
x_out_4_24,
x_out_4_25,
x_out_4_26,
x_out_4_27,
x_out_4_28,
x_out_4_29,
x_out_4_3,
x_out_4_30,
x_out_4_31,
x_out_4_32,
x_out_4_33,
x_out_4_4,
x_out_4_5,
x_out_4_6,
x_out_4_7,
x_out_4_8,
x_out_4_9,
x_out_50_0,
x_out_50_1,
x_out_50_10,
x_out_50_11,
x_out_50_12,
x_out_50_13,
x_out_50_14,
x_out_50_15,
x_out_50_18,
x_out_50_19,
x_out_50_2,
x_out_50_20,
x_out_50_21,
x_out_50_22,
x_out_50_23,
x_out_50_24,
x_out_50_25,
x_out_50_26,
x_out_50_27,
x_out_50_28,
x_out_50_29,
x_out_50_3,
x_out_50_30,
x_out_50_31,
x_out_50_32,
x_out_50_33,
x_out_50_4,
x_out_50_5,
x_out_50_6,
x_out_50_7,
x_out_50_8,
x_out_50_9,
x_out_51_0,
x_out_51_1,
x_out_51_10,
x_out_51_11,
x_out_51_12,
x_out_51_13,
x_out_51_14,
x_out_51_15,
x_out_51_18,
x_out_51_19,
x_out_51_2,
x_out_51_20,
x_out_51_21,
x_out_51_22,
x_out_51_23,
x_out_51_24,
x_out_51_25,
x_out_51_26,
x_out_51_27,
x_out_51_28,
x_out_51_29,
x_out_51_3,
x_out_51_30,
x_out_51_31,
x_out_51_32,
x_out_51_33,
x_out_51_4,
x_out_51_5,
x_out_51_6,
x_out_51_7,
x_out_51_8,
x_out_51_9,
x_out_52_0,
x_out_52_1,
x_out_52_10,
x_out_52_11,
x_out_52_12,
x_out_52_13,
x_out_52_14,
x_out_52_15,
x_out_52_2,
x_out_52_3,
x_out_52_4,
x_out_52_5,
x_out_52_6,
x_out_52_7,
x_out_52_8,
x_out_52_9,
x_out_53_0,
x_out_53_1,
x_out_53_10,
x_out_53_11,
x_out_53_12,
x_out_53_13,
x_out_53_14,
x_out_53_15,
x_out_53_18,
x_out_53_19,
x_out_53_2,
x_out_53_20,
x_out_53_21,
x_out_53_22,
x_out_53_23,
x_out_53_24,
x_out_53_25,
x_out_53_26,
x_out_53_27,
x_out_53_28,
x_out_53_29,
x_out_53_3,
x_out_53_30,
x_out_53_31,
x_out_53_32,
x_out_53_33,
x_out_53_4,
x_out_53_5,
x_out_53_6,
x_out_53_7,
x_out_53_8,
x_out_53_9,
x_out_54_0,
x_out_54_1,
x_out_54_10,
x_out_54_11,
x_out_54_12,
x_out_54_13,
x_out_54_14,
x_out_54_15,
x_out_54_18,
x_out_54_19,
x_out_54_2,
x_out_54_20,
x_out_54_21,
x_out_54_22,
x_out_54_23,
x_out_54_24,
x_out_54_25,
x_out_54_26,
x_out_54_27,
x_out_54_28,
x_out_54_29,
x_out_54_3,
x_out_54_30,
x_out_54_31,
x_out_54_32,
x_out_54_33,
x_out_54_4,
x_out_54_5,
x_out_54_6,
x_out_54_7,
x_out_54_8,
x_out_54_9,
x_out_55_0,
x_out_55_1,
x_out_55_10,
x_out_55_11,
x_out_55_12,
x_out_55_13,
x_out_55_14,
x_out_55_15,
x_out_55_18,
x_out_55_19,
x_out_55_2,
x_out_55_20,
x_out_55_21,
x_out_55_22,
x_out_55_23,
x_out_55_24,
x_out_55_25,
x_out_55_26,
x_out_55_27,
x_out_55_28,
x_out_55_29,
x_out_55_3,
x_out_55_30,
x_out_55_31,
x_out_55_32,
x_out_55_33,
x_out_55_4,
x_out_55_5,
x_out_55_6,
x_out_55_7,
x_out_55_8,
x_out_55_9,
x_out_56_0,
x_out_56_1,
x_out_56_10,
x_out_56_11,
x_out_56_12,
x_out_56_13,
x_out_56_14,
x_out_56_15,
x_out_56_18,
x_out_56_19,
x_out_56_2,
x_out_56_20,
x_out_56_21,
x_out_56_22,
x_out_56_23,
x_out_56_24,
x_out_56_25,
x_out_56_26,
x_out_56_27,
x_out_56_28,
x_out_56_29,
x_out_56_3,
x_out_56_30,
x_out_56_31,
x_out_56_32,
x_out_56_33,
x_out_56_4,
x_out_56_5,
x_out_56_6,
x_out_56_7,
x_out_56_8,
x_out_56_9,
x_out_57_0,
x_out_57_1,
x_out_57_10,
x_out_57_11,
x_out_57_12,
x_out_57_13,
x_out_57_14,
x_out_57_15,
x_out_57_18,
x_out_57_19,
x_out_57_2,
x_out_57_20,
x_out_57_21,
x_out_57_22,
x_out_57_23,
x_out_57_24,
x_out_57_25,
x_out_57_26,
x_out_57_27,
x_out_57_28,
x_out_57_29,
x_out_57_3,
x_out_57_30,
x_out_57_31,
x_out_57_32,
x_out_57_33,
x_out_57_4,
x_out_57_5,
x_out_57_6,
x_out_57_7,
x_out_57_8,
x_out_57_9,
x_out_58_0,
x_out_58_1,
x_out_58_10,
x_out_58_11,
x_out_58_12,
x_out_58_13,
x_out_58_14,
x_out_58_15,
x_out_58_18,
x_out_58_19,
x_out_58_2,
x_out_58_20,
x_out_58_21,
x_out_58_22,
x_out_58_23,
x_out_58_24,
x_out_58_25,
x_out_58_26,
x_out_58_27,
x_out_58_28,
x_out_58_29,
x_out_58_3,
x_out_58_30,
x_out_58_31,
x_out_58_32,
x_out_58_33,
x_out_58_4,
x_out_58_5,
x_out_58_6,
x_out_58_7,
x_out_58_8,
x_out_58_9,
x_out_59_0,
x_out_59_1,
x_out_59_10,
x_out_59_11,
x_out_59_12,
x_out_59_13,
x_out_59_14,
x_out_59_15,
x_out_59_18,
x_out_59_19,
x_out_59_2,
x_out_59_20,
x_out_59_21,
x_out_59_22,
x_out_59_23,
x_out_59_24,
x_out_59_25,
x_out_59_26,
x_out_59_27,
x_out_59_28,
x_out_59_29,
x_out_59_3,
x_out_59_30,
x_out_59_31,
x_out_59_32,
x_out_59_33,
x_out_59_4,
x_out_59_5,
x_out_59_6,
x_out_59_7,
x_out_59_8,
x_out_59_9,
x_out_5_0,
x_out_5_1,
x_out_5_10,
x_out_5_11,
x_out_5_12,
x_out_5_13,
x_out_5_14,
x_out_5_15,
x_out_5_18,
x_out_5_19,
x_out_5_2,
x_out_5_20,
x_out_5_21,
x_out_5_22,
x_out_5_23,
x_out_5_24,
x_out_5_25,
x_out_5_26,
x_out_5_27,
x_out_5_28,
x_out_5_29,
x_out_5_3,
x_out_5_30,
x_out_5_31,
x_out_5_32,
x_out_5_33,
x_out_5_4,
x_out_5_5,
x_out_5_6,
x_out_5_7,
x_out_5_8,
x_out_5_9,
x_out_60_0,
x_out_60_1,
x_out_60_10,
x_out_60_11,
x_out_60_12,
x_out_60_13,
x_out_60_14,
x_out_60_15,
x_out_60_18,
x_out_60_19,
x_out_60_2,
x_out_60_20,
x_out_60_21,
x_out_60_22,
x_out_60_23,
x_out_60_24,
x_out_60_25,
x_out_60_26,
x_out_60_27,
x_out_60_28,
x_out_60_29,
x_out_60_3,
x_out_60_30,
x_out_60_31,
x_out_60_32,
x_out_60_33,
x_out_60_4,
x_out_60_5,
x_out_60_6,
x_out_60_7,
x_out_60_8,
x_out_60_9,
x_out_61_0,
x_out_61_1,
x_out_61_10,
x_out_61_11,
x_out_61_12,
x_out_61_13,
x_out_61_14,
x_out_61_15,
x_out_61_18,
x_out_61_19,
x_out_61_2,
x_out_61_20,
x_out_61_21,
x_out_61_22,
x_out_61_23,
x_out_61_24,
x_out_61_25,
x_out_61_26,
x_out_61_27,
x_out_61_28,
x_out_61_29,
x_out_61_3,
x_out_61_30,
x_out_61_31,
x_out_61_32,
x_out_61_33,
x_out_61_4,
x_out_61_5,
x_out_61_6,
x_out_61_7,
x_out_61_8,
x_out_61_9,
x_out_62_0,
x_out_62_1,
x_out_62_10,
x_out_62_11,
x_out_62_12,
x_out_62_13,
x_out_62_14,
x_out_62_15,
x_out_62_18,
x_out_62_19,
x_out_62_2,
x_out_62_20,
x_out_62_21,
x_out_62_22,
x_out_62_23,
x_out_62_24,
x_out_62_25,
x_out_62_26,
x_out_62_27,
x_out_62_28,
x_out_62_29,
x_out_62_3,
x_out_62_30,
x_out_62_31,
x_out_62_32,
x_out_62_33,
x_out_62_4,
x_out_62_5,
x_out_62_6,
x_out_62_7,
x_out_62_8,
x_out_62_9,
x_out_63_0,
x_out_63_1,
x_out_63_10,
x_out_63_11,
x_out_63_12,
x_out_63_13,
x_out_63_14,
x_out_63_15,
x_out_63_18,
x_out_63_19,
x_out_63_2,
x_out_63_20,
x_out_63_21,
x_out_63_22,
x_out_63_23,
x_out_63_24,
x_out_63_25,
x_out_63_26,
x_out_63_27,
x_out_63_28,
x_out_63_29,
x_out_63_3,
x_out_63_30,
x_out_63_31,
x_out_63_32,
x_out_63_33,
x_out_63_4,
x_out_63_5,
x_out_63_6,
x_out_63_7,
x_out_63_8,
x_out_63_9,
x_out_6_0,
x_out_6_1,
x_out_6_10,
x_out_6_11,
x_out_6_12,
x_out_6_13,
x_out_6_14,
x_out_6_15,
x_out_6_18,
x_out_6_19,
x_out_6_2,
x_out_6_20,
x_out_6_21,
x_out_6_22,
x_out_6_23,
x_out_6_24,
x_out_6_25,
x_out_6_26,
x_out_6_27,
x_out_6_28,
x_out_6_29,
x_out_6_3,
x_out_6_30,
x_out_6_31,
x_out_6_32,
x_out_6_33,
x_out_6_4,
x_out_6_5,
x_out_6_6,
x_out_6_7,
x_out_6_8,
x_out_6_9,
x_out_7_0,
x_out_7_1,
x_out_7_10,
x_out_7_11,
x_out_7_12,
x_out_7_13,
x_out_7_14,
x_out_7_15,
x_out_7_18,
x_out_7_19,
x_out_7_2,
x_out_7_20,
x_out_7_21,
x_out_7_22,
x_out_7_23,
x_out_7_24,
x_out_7_25,
x_out_7_26,
x_out_7_27,
x_out_7_28,
x_out_7_29,
x_out_7_3,
x_out_7_30,
x_out_7_31,
x_out_7_32,
x_out_7_33,
x_out_7_4,
x_out_7_5,
x_out_7_6,
x_out_7_7,
x_out_7_8,
x_out_7_9,
x_out_8_0,
x_out_8_1,
x_out_8_10,
x_out_8_11,
x_out_8_12,
x_out_8_13,
x_out_8_14,
x_out_8_15,
x_out_8_18,
x_out_8_19,
x_out_8_2,
x_out_8_20,
x_out_8_21,
x_out_8_22,
x_out_8_23,
x_out_8_24,
x_out_8_25,
x_out_8_26,
x_out_8_27,
x_out_8_28,
x_out_8_29,
x_out_8_3,
x_out_8_30,
x_out_8_31,
x_out_8_32,
x_out_8_33,
x_out_8_4,
x_out_8_5,
x_out_8_6,
x_out_8_7,
x_out_8_8,
x_out_8_9,
x_out_9_0,
x_out_9_1,
x_out_9_10,
x_out_9_11,
x_out_9_12,
x_out_9_13,
x_out_9_14,
x_out_9_15,
x_out_9_18,
x_out_9_19,
x_out_9_2,
x_out_9_20,
x_out_9_21,
x_out_9_22,
x_out_9_23,
x_out_9_24,
x_out_9_25,
x_out_9_26,
x_out_9_27,
x_out_9_28,
x_out_9_29,
x_out_9_3,
x_out_9_30,
x_out_9_31,
x_out_9_32,
x_out_9_33,
x_out_9_4,
x_out_9_5,
x_out_9_6,
x_out_9_7,
x_out_9_8,
x_out_9_9
);

// Start PIs
input ispd_clk;
input rst;
input x_in_0_0;
input x_in_0_1;
input x_in_0_10;
input x_in_0_11;
input x_in_0_12;
input x_in_0_13;
input x_in_0_14;
input x_in_0_15;
input x_in_0_2;
input x_in_0_3;
input x_in_0_4;
input x_in_0_5;
input x_in_0_6;
input x_in_0_7;
input x_in_0_8;
input x_in_0_9;
input x_in_10_0;
input x_in_10_1;
input x_in_10_10;
input x_in_10_11;
input x_in_10_12;
input x_in_10_13;
input x_in_10_14;
input x_in_10_15;
input x_in_10_2;
input x_in_10_3;
input x_in_10_4;
input x_in_10_5;
input x_in_10_6;
input x_in_10_7;
input x_in_10_8;
input x_in_10_9;
input x_in_11_0;
input x_in_11_1;
input x_in_11_10;
input x_in_11_11;
input x_in_11_12;
input x_in_11_13;
input x_in_11_14;
input x_in_11_15;
input x_in_11_2;
input x_in_11_3;
input x_in_11_4;
input x_in_11_5;
input x_in_11_6;
input x_in_11_7;
input x_in_11_8;
input x_in_11_9;
input x_in_12_0;
input x_in_12_1;
input x_in_12_10;
input x_in_12_11;
input x_in_12_12;
input x_in_12_13;
input x_in_12_14;
input x_in_12_15;
input x_in_12_2;
input x_in_12_3;
input x_in_12_4;
input x_in_12_5;
input x_in_12_6;
input x_in_12_7;
input x_in_12_8;
input x_in_12_9;
input x_in_13_0;
input x_in_13_1;
input x_in_13_10;
input x_in_13_11;
input x_in_13_12;
input x_in_13_13;
input x_in_13_14;
input x_in_13_15;
input x_in_13_2;
input x_in_13_3;
input x_in_13_4;
input x_in_13_5;
input x_in_13_6;
input x_in_13_7;
input x_in_13_8;
input x_in_13_9;
input x_in_14_0;
input x_in_14_1;
input x_in_14_10;
input x_in_14_11;
input x_in_14_12;
input x_in_14_13;
input x_in_14_14;
input x_in_14_15;
input x_in_14_2;
input x_in_14_3;
input x_in_14_4;
input x_in_14_5;
input x_in_14_6;
input x_in_14_7;
input x_in_14_8;
input x_in_14_9;
input x_in_15_0;
input x_in_15_1;
input x_in_15_10;
input x_in_15_11;
input x_in_15_12;
input x_in_15_13;
input x_in_15_14;
input x_in_15_15;
input x_in_15_2;
input x_in_15_3;
input x_in_15_4;
input x_in_15_5;
input x_in_15_6;
input x_in_15_7;
input x_in_15_8;
input x_in_15_9;
input x_in_16_0;
input x_in_16_1;
input x_in_16_10;
input x_in_16_11;
input x_in_16_12;
input x_in_16_13;
input x_in_16_14;
input x_in_16_15;
input x_in_16_2;
input x_in_16_3;
input x_in_16_4;
input x_in_16_5;
input x_in_16_6;
input x_in_16_7;
input x_in_16_8;
input x_in_16_9;
input x_in_17_0;
input x_in_17_1;
input x_in_17_10;
input x_in_17_11;
input x_in_17_12;
input x_in_17_13;
input x_in_17_14;
input x_in_17_15;
input x_in_17_2;
input x_in_17_3;
input x_in_17_4;
input x_in_17_5;
input x_in_17_6;
input x_in_17_7;
input x_in_17_8;
input x_in_17_9;
input x_in_18_0;
input x_in_18_1;
input x_in_18_10;
input x_in_18_11;
input x_in_18_12;
input x_in_18_13;
input x_in_18_14;
input x_in_18_15;
input x_in_18_2;
input x_in_18_3;
input x_in_18_4;
input x_in_18_5;
input x_in_18_6;
input x_in_18_7;
input x_in_18_8;
input x_in_18_9;
input x_in_19_0;
input x_in_19_1;
input x_in_19_10;
input x_in_19_11;
input x_in_19_12;
input x_in_19_13;
input x_in_19_14;
input x_in_19_15;
input x_in_19_2;
input x_in_19_3;
input x_in_19_4;
input x_in_19_5;
input x_in_19_6;
input x_in_19_7;
input x_in_19_8;
input x_in_19_9;
input x_in_1_0;
input x_in_1_1;
input x_in_1_10;
input x_in_1_11;
input x_in_1_12;
input x_in_1_13;
input x_in_1_14;
input x_in_1_15;
input x_in_1_2;
input x_in_1_3;
input x_in_1_4;
input x_in_1_5;
input x_in_1_6;
input x_in_1_7;
input x_in_1_8;
input x_in_1_9;
input x_in_20_0;
input x_in_20_1;
input x_in_20_10;
input x_in_20_11;
input x_in_20_12;
input x_in_20_13;
input x_in_20_14;
input x_in_20_15;
input x_in_20_2;
input x_in_20_3;
input x_in_20_4;
input x_in_20_5;
input x_in_20_6;
input x_in_20_7;
input x_in_20_8;
input x_in_20_9;
input x_in_21_0;
input x_in_21_1;
input x_in_21_10;
input x_in_21_11;
input x_in_21_12;
input x_in_21_13;
input x_in_21_14;
input x_in_21_15;
input x_in_21_2;
input x_in_21_3;
input x_in_21_4;
input x_in_21_5;
input x_in_21_6;
input x_in_21_7;
input x_in_21_8;
input x_in_21_9;
input x_in_22_0;
input x_in_22_1;
input x_in_22_10;
input x_in_22_11;
input x_in_22_12;
input x_in_22_13;
input x_in_22_14;
input x_in_22_15;
input x_in_22_2;
input x_in_22_3;
input x_in_22_4;
input x_in_22_5;
input x_in_22_6;
input x_in_22_7;
input x_in_22_8;
input x_in_22_9;
input x_in_23_0;
input x_in_23_1;
input x_in_23_10;
input x_in_23_11;
input x_in_23_12;
input x_in_23_13;
input x_in_23_14;
input x_in_23_15;
input x_in_23_2;
input x_in_23_3;
input x_in_23_4;
input x_in_23_5;
input x_in_23_6;
input x_in_23_7;
input x_in_23_8;
input x_in_23_9;
input x_in_24_0;
input x_in_24_1;
input x_in_24_10;
input x_in_24_11;
input x_in_24_12;
input x_in_24_13;
input x_in_24_14;
input x_in_24_15;
input x_in_24_2;
input x_in_24_3;
input x_in_24_4;
input x_in_24_5;
input x_in_24_6;
input x_in_24_7;
input x_in_24_8;
input x_in_24_9;
input x_in_25_0;
input x_in_25_1;
input x_in_25_10;
input x_in_25_11;
input x_in_25_12;
input x_in_25_13;
input x_in_25_14;
input x_in_25_15;
input x_in_25_2;
input x_in_25_3;
input x_in_25_4;
input x_in_25_5;
input x_in_25_6;
input x_in_25_7;
input x_in_25_8;
input x_in_25_9;
input x_in_26_0;
input x_in_26_1;
input x_in_26_10;
input x_in_26_11;
input x_in_26_12;
input x_in_26_13;
input x_in_26_14;
input x_in_26_15;
input x_in_26_2;
input x_in_26_3;
input x_in_26_4;
input x_in_26_5;
input x_in_26_6;
input x_in_26_7;
input x_in_26_8;
input x_in_26_9;
input x_in_27_0;
input x_in_27_1;
input x_in_27_10;
input x_in_27_11;
input x_in_27_12;
input x_in_27_13;
input x_in_27_14;
input x_in_27_15;
input x_in_27_2;
input x_in_27_3;
input x_in_27_4;
input x_in_27_5;
input x_in_27_6;
input x_in_27_7;
input x_in_27_8;
input x_in_27_9;
input x_in_28_0;
input x_in_28_1;
input x_in_28_10;
input x_in_28_11;
input x_in_28_12;
input x_in_28_13;
input x_in_28_14;
input x_in_28_15;
input x_in_28_2;
input x_in_28_3;
input x_in_28_4;
input x_in_28_5;
input x_in_28_6;
input x_in_28_7;
input x_in_28_8;
input x_in_28_9;
input x_in_29_0;
input x_in_29_1;
input x_in_29_10;
input x_in_29_11;
input x_in_29_12;
input x_in_29_13;
input x_in_29_14;
input x_in_29_15;
input x_in_29_2;
input x_in_29_3;
input x_in_29_4;
input x_in_29_5;
input x_in_29_6;
input x_in_29_7;
input x_in_29_8;
input x_in_29_9;
input x_in_2_0;
input x_in_2_1;
input x_in_2_10;
input x_in_2_11;
input x_in_2_12;
input x_in_2_13;
input x_in_2_14;
input x_in_2_15;
input x_in_2_2;
input x_in_2_3;
input x_in_2_4;
input x_in_2_5;
input x_in_2_6;
input x_in_2_7;
input x_in_2_8;
input x_in_2_9;
input x_in_30_0;
input x_in_30_1;
input x_in_30_10;
input x_in_30_11;
input x_in_30_12;
input x_in_30_13;
input x_in_30_14;
input x_in_30_15;
input x_in_30_2;
input x_in_30_3;
input x_in_30_4;
input x_in_30_5;
input x_in_30_6;
input x_in_30_7;
input x_in_30_8;
input x_in_30_9;
input x_in_31_0;
input x_in_31_1;
input x_in_31_10;
input x_in_31_11;
input x_in_31_12;
input x_in_31_13;
input x_in_31_14;
input x_in_31_15;
input x_in_31_2;
input x_in_31_3;
input x_in_31_4;
input x_in_31_5;
input x_in_31_6;
input x_in_31_7;
input x_in_31_8;
input x_in_31_9;
input x_in_32_0;
input x_in_32_1;
input x_in_32_10;
input x_in_32_11;
input x_in_32_12;
input x_in_32_13;
input x_in_32_14;
input x_in_32_15;
input x_in_32_2;
input x_in_32_3;
input x_in_32_4;
input x_in_32_5;
input x_in_32_6;
input x_in_32_7;
input x_in_32_8;
input x_in_32_9;
input x_in_33_0;
input x_in_33_1;
input x_in_33_10;
input x_in_33_11;
input x_in_33_12;
input x_in_33_13;
input x_in_33_14;
input x_in_33_15;
input x_in_33_2;
input x_in_33_3;
input x_in_33_4;
input x_in_33_5;
input x_in_33_6;
input x_in_33_7;
input x_in_33_8;
input x_in_33_9;
input x_in_34_0;
input x_in_34_1;
input x_in_34_10;
input x_in_34_11;
input x_in_34_12;
input x_in_34_13;
input x_in_34_14;
input x_in_34_15;
input x_in_34_2;
input x_in_34_3;
input x_in_34_4;
input x_in_34_5;
input x_in_34_6;
input x_in_34_7;
input x_in_34_8;
input x_in_34_9;
input x_in_35_0;
input x_in_35_1;
input x_in_35_10;
input x_in_35_11;
input x_in_35_12;
input x_in_35_13;
input x_in_35_14;
input x_in_35_15;
input x_in_35_2;
input x_in_35_3;
input x_in_35_4;
input x_in_35_5;
input x_in_35_6;
input x_in_35_7;
input x_in_35_8;
input x_in_35_9;
input x_in_36_0;
input x_in_36_1;
input x_in_36_10;
input x_in_36_11;
input x_in_36_12;
input x_in_36_13;
input x_in_36_14;
input x_in_36_15;
input x_in_36_2;
input x_in_36_3;
input x_in_36_4;
input x_in_36_5;
input x_in_36_6;
input x_in_36_7;
input x_in_36_8;
input x_in_36_9;
input x_in_37_0;
input x_in_37_1;
input x_in_37_10;
input x_in_37_11;
input x_in_37_12;
input x_in_37_13;
input x_in_37_14;
input x_in_37_15;
input x_in_37_2;
input x_in_37_3;
input x_in_37_4;
input x_in_37_5;
input x_in_37_6;
input x_in_37_7;
input x_in_37_8;
input x_in_37_9;
input x_in_38_0;
input x_in_38_1;
input x_in_38_10;
input x_in_38_11;
input x_in_38_12;
input x_in_38_13;
input x_in_38_14;
input x_in_38_15;
input x_in_38_2;
input x_in_38_3;
input x_in_38_4;
input x_in_38_5;
input x_in_38_6;
input x_in_38_7;
input x_in_38_8;
input x_in_38_9;
input x_in_39_0;
input x_in_39_1;
input x_in_39_10;
input x_in_39_11;
input x_in_39_12;
input x_in_39_13;
input x_in_39_14;
input x_in_39_15;
input x_in_39_2;
input x_in_39_3;
input x_in_39_4;
input x_in_39_5;
input x_in_39_6;
input x_in_39_7;
input x_in_39_8;
input x_in_39_9;
input x_in_3_0;
input x_in_3_1;
input x_in_3_10;
input x_in_3_11;
input x_in_3_12;
input x_in_3_13;
input x_in_3_14;
input x_in_3_15;
input x_in_3_2;
input x_in_3_3;
input x_in_3_4;
input x_in_3_5;
input x_in_3_6;
input x_in_3_7;
input x_in_3_8;
input x_in_3_9;
input x_in_40_0;
input x_in_40_1;
input x_in_40_10;
input x_in_40_11;
input x_in_40_12;
input x_in_40_13;
input x_in_40_14;
input x_in_40_15;
input x_in_40_2;
input x_in_40_3;
input x_in_40_4;
input x_in_40_5;
input x_in_40_6;
input x_in_40_7;
input x_in_40_8;
input x_in_40_9;
input x_in_41_0;
input x_in_41_1;
input x_in_41_10;
input x_in_41_11;
input x_in_41_12;
input x_in_41_13;
input x_in_41_14;
input x_in_41_15;
input x_in_41_2;
input x_in_41_3;
input x_in_41_4;
input x_in_41_5;
input x_in_41_6;
input x_in_41_7;
input x_in_41_8;
input x_in_41_9;
input x_in_42_0;
input x_in_42_1;
input x_in_42_10;
input x_in_42_11;
input x_in_42_12;
input x_in_42_13;
input x_in_42_14;
input x_in_42_15;
input x_in_42_2;
input x_in_42_3;
input x_in_42_4;
input x_in_42_5;
input x_in_42_6;
input x_in_42_7;
input x_in_42_8;
input x_in_42_9;
input x_in_43_0;
input x_in_43_1;
input x_in_43_10;
input x_in_43_11;
input x_in_43_12;
input x_in_43_13;
input x_in_43_14;
input x_in_43_15;
input x_in_43_2;
input x_in_43_3;
input x_in_43_4;
input x_in_43_5;
input x_in_43_6;
input x_in_43_7;
input x_in_43_8;
input x_in_43_9;
input x_in_44_0;
input x_in_44_1;
input x_in_44_10;
input x_in_44_11;
input x_in_44_12;
input x_in_44_13;
input x_in_44_14;
input x_in_44_15;
input x_in_44_2;
input x_in_44_3;
input x_in_44_4;
input x_in_44_5;
input x_in_44_6;
input x_in_44_7;
input x_in_44_8;
input x_in_44_9;
input x_in_45_0;
input x_in_45_1;
input x_in_45_10;
input x_in_45_11;
input x_in_45_12;
input x_in_45_13;
input x_in_45_14;
input x_in_45_15;
input x_in_45_2;
input x_in_45_3;
input x_in_45_4;
input x_in_45_5;
input x_in_45_6;
input x_in_45_7;
input x_in_45_8;
input x_in_45_9;
input x_in_46_0;
input x_in_46_1;
input x_in_46_10;
input x_in_46_11;
input x_in_46_12;
input x_in_46_13;
input x_in_46_14;
input x_in_46_15;
input x_in_46_2;
input x_in_46_3;
input x_in_46_4;
input x_in_46_5;
input x_in_46_6;
input x_in_46_7;
input x_in_46_8;
input x_in_46_9;
input x_in_47_0;
input x_in_47_1;
input x_in_47_10;
input x_in_47_11;
input x_in_47_12;
input x_in_47_13;
input x_in_47_14;
input x_in_47_15;
input x_in_47_2;
input x_in_47_3;
input x_in_47_4;
input x_in_47_5;
input x_in_47_6;
input x_in_47_7;
input x_in_47_8;
input x_in_47_9;
input x_in_48_0;
input x_in_48_1;
input x_in_48_10;
input x_in_48_11;
input x_in_48_12;
input x_in_48_13;
input x_in_48_14;
input x_in_48_15;
input x_in_48_2;
input x_in_48_3;
input x_in_48_4;
input x_in_48_5;
input x_in_48_6;
input x_in_48_7;
input x_in_48_8;
input x_in_48_9;
input x_in_49_0;
input x_in_49_1;
input x_in_49_10;
input x_in_49_11;
input x_in_49_12;
input x_in_49_13;
input x_in_49_14;
input x_in_49_15;
input x_in_49_2;
input x_in_49_3;
input x_in_49_4;
input x_in_49_5;
input x_in_49_6;
input x_in_49_7;
input x_in_49_8;
input x_in_49_9;
input x_in_4_0;
input x_in_4_1;
input x_in_4_10;
input x_in_4_11;
input x_in_4_12;
input x_in_4_13;
input x_in_4_14;
input x_in_4_15;
input x_in_4_2;
input x_in_4_3;
input x_in_4_4;
input x_in_4_5;
input x_in_4_6;
input x_in_4_7;
input x_in_4_8;
input x_in_4_9;
input x_in_50_0;
input x_in_50_1;
input x_in_50_10;
input x_in_50_11;
input x_in_50_12;
input x_in_50_13;
input x_in_50_14;
input x_in_50_15;
input x_in_50_2;
input x_in_50_3;
input x_in_50_4;
input x_in_50_5;
input x_in_50_6;
input x_in_50_7;
input x_in_50_8;
input x_in_50_9;
input x_in_51_0;
input x_in_51_1;
input x_in_51_10;
input x_in_51_11;
input x_in_51_12;
input x_in_51_13;
input x_in_51_14;
input x_in_51_15;
input x_in_51_2;
input x_in_51_3;
input x_in_51_4;
input x_in_51_5;
input x_in_51_6;
input x_in_51_7;
input x_in_51_8;
input x_in_51_9;
input x_in_52_0;
input x_in_52_1;
input x_in_52_10;
input x_in_52_11;
input x_in_52_12;
input x_in_52_13;
input x_in_52_14;
input x_in_52_15;
input x_in_52_2;
input x_in_52_3;
input x_in_52_4;
input x_in_52_5;
input x_in_52_6;
input x_in_52_7;
input x_in_52_8;
input x_in_52_9;
input x_in_53_0;
input x_in_53_1;
input x_in_53_10;
input x_in_53_11;
input x_in_53_12;
input x_in_53_13;
input x_in_53_14;
input x_in_53_15;
input x_in_53_2;
input x_in_53_3;
input x_in_53_4;
input x_in_53_5;
input x_in_53_6;
input x_in_53_7;
input x_in_53_8;
input x_in_53_9;
input x_in_54_0;
input x_in_54_1;
input x_in_54_10;
input x_in_54_11;
input x_in_54_12;
input x_in_54_13;
input x_in_54_14;
input x_in_54_15;
input x_in_54_2;
input x_in_54_3;
input x_in_54_4;
input x_in_54_5;
input x_in_54_6;
input x_in_54_7;
input x_in_54_8;
input x_in_54_9;
input x_in_55_0;
input x_in_55_1;
input x_in_55_10;
input x_in_55_11;
input x_in_55_12;
input x_in_55_13;
input x_in_55_14;
input x_in_55_15;
input x_in_55_2;
input x_in_55_3;
input x_in_55_4;
input x_in_55_5;
input x_in_55_6;
input x_in_55_7;
input x_in_55_8;
input x_in_55_9;
input x_in_56_0;
input x_in_56_1;
input x_in_56_10;
input x_in_56_11;
input x_in_56_12;
input x_in_56_13;
input x_in_56_14;
input x_in_56_15;
input x_in_56_2;
input x_in_56_3;
input x_in_56_4;
input x_in_56_5;
input x_in_56_6;
input x_in_56_7;
input x_in_56_8;
input x_in_56_9;
input x_in_57_0;
input x_in_57_1;
input x_in_57_10;
input x_in_57_11;
input x_in_57_12;
input x_in_57_13;
input x_in_57_14;
input x_in_57_15;
input x_in_57_2;
input x_in_57_3;
input x_in_57_4;
input x_in_57_5;
input x_in_57_6;
input x_in_57_7;
input x_in_57_8;
input x_in_57_9;
input x_in_58_0;
input x_in_58_1;
input x_in_58_10;
input x_in_58_11;
input x_in_58_12;
input x_in_58_13;
input x_in_58_14;
input x_in_58_15;
input x_in_58_2;
input x_in_58_3;
input x_in_58_4;
input x_in_58_5;
input x_in_58_6;
input x_in_58_7;
input x_in_58_8;
input x_in_58_9;
input x_in_59_0;
input x_in_59_1;
input x_in_59_10;
input x_in_59_11;
input x_in_59_12;
input x_in_59_13;
input x_in_59_14;
input x_in_59_15;
input x_in_59_2;
input x_in_59_3;
input x_in_59_4;
input x_in_59_5;
input x_in_59_6;
input x_in_59_7;
input x_in_59_8;
input x_in_59_9;
input x_in_5_0;
input x_in_5_1;
input x_in_5_10;
input x_in_5_11;
input x_in_5_12;
input x_in_5_13;
input x_in_5_14;
input x_in_5_15;
input x_in_5_2;
input x_in_5_3;
input x_in_5_4;
input x_in_5_5;
input x_in_5_6;
input x_in_5_7;
input x_in_5_8;
input x_in_5_9;
input x_in_60_0;
input x_in_60_1;
input x_in_60_10;
input x_in_60_11;
input x_in_60_12;
input x_in_60_13;
input x_in_60_14;
input x_in_60_15;
input x_in_60_2;
input x_in_60_3;
input x_in_60_4;
input x_in_60_5;
input x_in_60_6;
input x_in_60_7;
input x_in_60_8;
input x_in_60_9;
input x_in_61_0;
input x_in_61_1;
input x_in_61_10;
input x_in_61_11;
input x_in_61_12;
input x_in_61_13;
input x_in_61_14;
input x_in_61_15;
input x_in_61_2;
input x_in_61_3;
input x_in_61_4;
input x_in_61_5;
input x_in_61_6;
input x_in_61_7;
input x_in_61_8;
input x_in_61_9;
input x_in_62_0;
input x_in_62_1;
input x_in_62_10;
input x_in_62_11;
input x_in_62_12;
input x_in_62_13;
input x_in_62_14;
input x_in_62_15;
input x_in_62_2;
input x_in_62_3;
input x_in_62_4;
input x_in_62_5;
input x_in_62_6;
input x_in_62_7;
input x_in_62_8;
input x_in_62_9;
input x_in_63_0;
input x_in_63_1;
input x_in_63_10;
input x_in_63_11;
input x_in_63_12;
input x_in_63_13;
input x_in_63_14;
input x_in_63_15;
input x_in_63_2;
input x_in_63_3;
input x_in_63_4;
input x_in_63_5;
input x_in_63_6;
input x_in_63_7;
input x_in_63_8;
input x_in_63_9;
input x_in_6_0;
input x_in_6_1;
input x_in_6_10;
input x_in_6_11;
input x_in_6_12;
input x_in_6_13;
input x_in_6_14;
input x_in_6_15;
input x_in_6_2;
input x_in_6_3;
input x_in_6_4;
input x_in_6_5;
input x_in_6_6;
input x_in_6_7;
input x_in_6_8;
input x_in_6_9;
input x_in_7_0;
input x_in_7_1;
input x_in_7_10;
input x_in_7_11;
input x_in_7_12;
input x_in_7_13;
input x_in_7_14;
input x_in_7_15;
input x_in_7_2;
input x_in_7_3;
input x_in_7_4;
input x_in_7_5;
input x_in_7_6;
input x_in_7_7;
input x_in_7_8;
input x_in_7_9;
input x_in_8_0;
input x_in_8_1;
input x_in_8_10;
input x_in_8_11;
input x_in_8_12;
input x_in_8_13;
input x_in_8_14;
input x_in_8_15;
input x_in_8_2;
input x_in_8_3;
input x_in_8_4;
input x_in_8_5;
input x_in_8_6;
input x_in_8_7;
input x_in_8_8;
input x_in_8_9;
input x_in_9_0;
input x_in_9_1;
input x_in_9_10;
input x_in_9_11;
input x_in_9_12;
input x_in_9_13;
input x_in_9_14;
input x_in_9_15;
input x_in_9_2;
input x_in_9_3;
input x_in_9_4;
input x_in_9_5;
input x_in_9_6;
input x_in_9_7;
input x_in_9_8;
input x_in_9_9;

// Start POs
output x_out_0_0;
output x_out_0_1;
output x_out_0_10;
output x_out_0_11;
output x_out_0_12;
output x_out_0_13;
output x_out_0_14;
output x_out_0_15;
output x_out_0_2;
output x_out_0_3;
output x_out_0_4;
output x_out_0_5;
output x_out_0_6;
output x_out_0_7;
output x_out_0_8;
output x_out_0_9;
output x_out_10_0;
output x_out_10_1;
output x_out_10_10;
output x_out_10_11;
output x_out_10_12;
output x_out_10_13;
output x_out_10_14;
output x_out_10_15;
output x_out_10_18;
output x_out_10_19;
output x_out_10_2;
output x_out_10_20;
output x_out_10_21;
output x_out_10_22;
output x_out_10_23;
output x_out_10_24;
output x_out_10_25;
output x_out_10_26;
output x_out_10_27;
output x_out_10_28;
output x_out_10_29;
output x_out_10_3;
output x_out_10_30;
output x_out_10_31;
output x_out_10_32;
output x_out_10_33;
output x_out_10_4;
output x_out_10_5;
output x_out_10_6;
output x_out_10_7;
output x_out_10_8;
output x_out_10_9;
output x_out_11_0;
output x_out_11_1;
output x_out_11_10;
output x_out_11_11;
output x_out_11_12;
output x_out_11_13;
output x_out_11_14;
output x_out_11_15;
output x_out_11_18;
output x_out_11_19;
output x_out_11_2;
output x_out_11_20;
output x_out_11_21;
output x_out_11_22;
output x_out_11_23;
output x_out_11_24;
output x_out_11_25;
output x_out_11_26;
output x_out_11_27;
output x_out_11_28;
output x_out_11_29;
output x_out_11_3;
output x_out_11_30;
output x_out_11_31;
output x_out_11_32;
output x_out_11_33;
output x_out_11_4;
output x_out_11_5;
output x_out_11_6;
output x_out_11_7;
output x_out_11_8;
output x_out_11_9;
output x_out_12_0;
output x_out_12_1;
output x_out_12_10;
output x_out_12_11;
output x_out_12_12;
output x_out_12_13;
output x_out_12_14;
output x_out_12_15;
output x_out_12_18;
output x_out_12_19;
output x_out_12_2;
output x_out_12_20;
output x_out_12_21;
output x_out_12_22;
output x_out_12_23;
output x_out_12_24;
output x_out_12_25;
output x_out_12_26;
output x_out_12_27;
output x_out_12_28;
output x_out_12_29;
output x_out_12_3;
output x_out_12_30;
output x_out_12_31;
output x_out_12_32;
output x_out_12_33;
output x_out_12_4;
output x_out_12_5;
output x_out_12_6;
output x_out_12_7;
output x_out_12_8;
output x_out_12_9;
output x_out_13_0;
output x_out_13_1;
output x_out_13_10;
output x_out_13_11;
output x_out_13_12;
output x_out_13_13;
output x_out_13_14;
output x_out_13_15;
output x_out_13_18;
output x_out_13_19;
output x_out_13_2;
output x_out_13_20;
output x_out_13_21;
output x_out_13_22;
output x_out_13_23;
output x_out_13_24;
output x_out_13_25;
output x_out_13_26;
output x_out_13_27;
output x_out_13_28;
output x_out_13_29;
output x_out_13_3;
output x_out_13_30;
output x_out_13_31;
output x_out_13_32;
output x_out_13_33;
output x_out_13_4;
output x_out_13_5;
output x_out_13_6;
output x_out_13_7;
output x_out_13_8;
output x_out_13_9;
output x_out_14_0;
output x_out_14_1;
output x_out_14_10;
output x_out_14_11;
output x_out_14_12;
output x_out_14_13;
output x_out_14_14;
output x_out_14_15;
output x_out_14_18;
output x_out_14_19;
output x_out_14_2;
output x_out_14_20;
output x_out_14_21;
output x_out_14_22;
output x_out_14_23;
output x_out_14_24;
output x_out_14_25;
output x_out_14_26;
output x_out_14_27;
output x_out_14_28;
output x_out_14_29;
output x_out_14_3;
output x_out_14_30;
output x_out_14_31;
output x_out_14_32;
output x_out_14_33;
output x_out_14_4;
output x_out_14_5;
output x_out_14_6;
output x_out_14_7;
output x_out_14_8;
output x_out_14_9;
output x_out_15_0;
output x_out_15_1;
output x_out_15_10;
output x_out_15_11;
output x_out_15_12;
output x_out_15_13;
output x_out_15_14;
output x_out_15_15;
output x_out_15_18;
output x_out_15_19;
output x_out_15_2;
output x_out_15_20;
output x_out_15_21;
output x_out_15_22;
output x_out_15_23;
output x_out_15_24;
output x_out_15_25;
output x_out_15_26;
output x_out_15_27;
output x_out_15_28;
output x_out_15_29;
output x_out_15_3;
output x_out_15_30;
output x_out_15_31;
output x_out_15_32;
output x_out_15_33;
output x_out_15_4;
output x_out_15_5;
output x_out_15_6;
output x_out_15_7;
output x_out_15_8;
output x_out_15_9;
output x_out_16_0;
output x_out_16_1;
output x_out_16_10;
output x_out_16_11;
output x_out_16_12;
output x_out_16_13;
output x_out_16_14;
output x_out_16_15;
output x_out_16_18;
output x_out_16_19;
output x_out_16_2;
output x_out_16_20;
output x_out_16_21;
output x_out_16_22;
output x_out_16_23;
output x_out_16_24;
output x_out_16_25;
output x_out_16_26;
output x_out_16_27;
output x_out_16_28;
output x_out_16_29;
output x_out_16_3;
output x_out_16_30;
output x_out_16_31;
output x_out_16_32;
output x_out_16_33;
output x_out_16_4;
output x_out_16_5;
output x_out_16_6;
output x_out_16_7;
output x_out_16_8;
output x_out_16_9;
output x_out_17_0;
output x_out_17_1;
output x_out_17_10;
output x_out_17_11;
output x_out_17_12;
output x_out_17_13;
output x_out_17_14;
output x_out_17_15;
output x_out_17_18;
output x_out_17_19;
output x_out_17_2;
output x_out_17_20;
output x_out_17_21;
output x_out_17_22;
output x_out_17_23;
output x_out_17_24;
output x_out_17_25;
output x_out_17_26;
output x_out_17_27;
output x_out_17_28;
output x_out_17_29;
output x_out_17_3;
output x_out_17_30;
output x_out_17_31;
output x_out_17_32;
output x_out_17_33;
output x_out_17_4;
output x_out_17_5;
output x_out_17_6;
output x_out_17_7;
output x_out_17_8;
output x_out_17_9;
output x_out_18_0;
output x_out_18_1;
output x_out_18_10;
output x_out_18_11;
output x_out_18_12;
output x_out_18_13;
output x_out_18_14;
output x_out_18_15;
output x_out_18_18;
output x_out_18_19;
output x_out_18_2;
output x_out_18_20;
output x_out_18_21;
output x_out_18_22;
output x_out_18_23;
output x_out_18_24;
output x_out_18_25;
output x_out_18_26;
output x_out_18_27;
output x_out_18_28;
output x_out_18_29;
output x_out_18_3;
output x_out_18_30;
output x_out_18_31;
output x_out_18_32;
output x_out_18_33;
output x_out_18_4;
output x_out_18_5;
output x_out_18_6;
output x_out_18_7;
output x_out_18_8;
output x_out_18_9;
output x_out_19_0;
output x_out_19_1;
output x_out_19_10;
output x_out_19_11;
output x_out_19_12;
output x_out_19_13;
output x_out_19_14;
output x_out_19_15;
output x_out_19_18;
output x_out_19_19;
output x_out_19_2;
output x_out_19_20;
output x_out_19_21;
output x_out_19_22;
output x_out_19_23;
output x_out_19_24;
output x_out_19_25;
output x_out_19_26;
output x_out_19_27;
output x_out_19_28;
output x_out_19_29;
output x_out_19_3;
output x_out_19_30;
output x_out_19_31;
output x_out_19_32;
output x_out_19_33;
output x_out_19_4;
output x_out_19_5;
output x_out_19_6;
output x_out_19_7;
output x_out_19_8;
output x_out_19_9;
output x_out_1_0;
output x_out_1_1;
output x_out_1_10;
output x_out_1_11;
output x_out_1_12;
output x_out_1_13;
output x_out_1_14;
output x_out_1_15;
output x_out_1_18;
output x_out_1_19;
output x_out_1_2;
output x_out_1_20;
output x_out_1_21;
output x_out_1_22;
output x_out_1_23;
output x_out_1_24;
output x_out_1_25;
output x_out_1_26;
output x_out_1_27;
output x_out_1_28;
output x_out_1_29;
output x_out_1_3;
output x_out_1_30;
output x_out_1_31;
output x_out_1_32;
output x_out_1_33;
output x_out_1_4;
output x_out_1_5;
output x_out_1_6;
output x_out_1_7;
output x_out_1_8;
output x_out_1_9;
output x_out_20_0;
output x_out_20_1;
output x_out_20_10;
output x_out_20_11;
output x_out_20_12;
output x_out_20_13;
output x_out_20_14;
output x_out_20_15;
output x_out_20_2;
output x_out_20_3;
output x_out_20_4;
output x_out_20_5;
output x_out_20_6;
output x_out_20_7;
output x_out_20_8;
output x_out_20_9;
output x_out_21_0;
output x_out_21_1;
output x_out_21_10;
output x_out_21_11;
output x_out_21_12;
output x_out_21_13;
output x_out_21_14;
output x_out_21_15;
output x_out_21_18;
output x_out_21_19;
output x_out_21_2;
output x_out_21_20;
output x_out_21_21;
output x_out_21_22;
output x_out_21_23;
output x_out_21_24;
output x_out_21_25;
output x_out_21_26;
output x_out_21_27;
output x_out_21_28;
output x_out_21_29;
output x_out_21_3;
output x_out_21_30;
output x_out_21_31;
output x_out_21_32;
output x_out_21_33;
output x_out_21_4;
output x_out_21_5;
output x_out_21_6;
output x_out_21_7;
output x_out_21_8;
output x_out_21_9;
output x_out_22_0;
output x_out_22_1;
output x_out_22_10;
output x_out_22_11;
output x_out_22_12;
output x_out_22_13;
output x_out_22_14;
output x_out_22_15;
output x_out_22_18;
output x_out_22_19;
output x_out_22_2;
output x_out_22_20;
output x_out_22_21;
output x_out_22_22;
output x_out_22_23;
output x_out_22_24;
output x_out_22_25;
output x_out_22_26;
output x_out_22_27;
output x_out_22_28;
output x_out_22_29;
output x_out_22_3;
output x_out_22_30;
output x_out_22_31;
output x_out_22_32;
output x_out_22_33;
output x_out_22_4;
output x_out_22_5;
output x_out_22_6;
output x_out_22_7;
output x_out_22_8;
output x_out_22_9;
output x_out_23_0;
output x_out_23_1;
output x_out_23_10;
output x_out_23_11;
output x_out_23_12;
output x_out_23_13;
output x_out_23_14;
output x_out_23_15;
output x_out_23_18;
output x_out_23_19;
output x_out_23_2;
output x_out_23_20;
output x_out_23_21;
output x_out_23_22;
output x_out_23_23;
output x_out_23_24;
output x_out_23_25;
output x_out_23_26;
output x_out_23_27;
output x_out_23_28;
output x_out_23_29;
output x_out_23_3;
output x_out_23_30;
output x_out_23_31;
output x_out_23_32;
output x_out_23_33;
output x_out_23_4;
output x_out_23_5;
output x_out_23_6;
output x_out_23_7;
output x_out_23_8;
output x_out_23_9;
output x_out_24_0;
output x_out_24_1;
output x_out_24_10;
output x_out_24_11;
output x_out_24_12;
output x_out_24_13;
output x_out_24_14;
output x_out_24_15;
output x_out_24_18;
output x_out_24_19;
output x_out_24_2;
output x_out_24_20;
output x_out_24_21;
output x_out_24_22;
output x_out_24_23;
output x_out_24_24;
output x_out_24_25;
output x_out_24_26;
output x_out_24_27;
output x_out_24_28;
output x_out_24_29;
output x_out_24_3;
output x_out_24_30;
output x_out_24_31;
output x_out_24_32;
output x_out_24_33;
output x_out_24_4;
output x_out_24_5;
output x_out_24_6;
output x_out_24_7;
output x_out_24_8;
output x_out_24_9;
output x_out_25_0;
output x_out_25_1;
output x_out_25_10;
output x_out_25_11;
output x_out_25_12;
output x_out_25_13;
output x_out_25_14;
output x_out_25_15;
output x_out_25_18;
output x_out_25_19;
output x_out_25_2;
output x_out_25_20;
output x_out_25_21;
output x_out_25_22;
output x_out_25_23;
output x_out_25_24;
output x_out_25_25;
output x_out_25_26;
output x_out_25_27;
output x_out_25_28;
output x_out_25_29;
output x_out_25_3;
output x_out_25_30;
output x_out_25_31;
output x_out_25_32;
output x_out_25_33;
output x_out_25_4;
output x_out_25_5;
output x_out_25_6;
output x_out_25_7;
output x_out_25_8;
output x_out_25_9;
output x_out_26_0;
output x_out_26_1;
output x_out_26_10;
output x_out_26_11;
output x_out_26_12;
output x_out_26_13;
output x_out_26_14;
output x_out_26_15;
output x_out_26_18;
output x_out_26_19;
output x_out_26_2;
output x_out_26_20;
output x_out_26_21;
output x_out_26_22;
output x_out_26_23;
output x_out_26_24;
output x_out_26_25;
output x_out_26_26;
output x_out_26_27;
output x_out_26_28;
output x_out_26_29;
output x_out_26_3;
output x_out_26_30;
output x_out_26_31;
output x_out_26_32;
output x_out_26_33;
output x_out_26_4;
output x_out_26_5;
output x_out_26_6;
output x_out_26_7;
output x_out_26_8;
output x_out_26_9;
output x_out_27_0;
output x_out_27_1;
output x_out_27_10;
output x_out_27_11;
output x_out_27_12;
output x_out_27_13;
output x_out_27_14;
output x_out_27_15;
output x_out_27_18;
output x_out_27_19;
output x_out_27_2;
output x_out_27_20;
output x_out_27_21;
output x_out_27_22;
output x_out_27_23;
output x_out_27_24;
output x_out_27_25;
output x_out_27_26;
output x_out_27_27;
output x_out_27_28;
output x_out_27_29;
output x_out_27_3;
output x_out_27_30;
output x_out_27_31;
output x_out_27_32;
output x_out_27_33;
output x_out_27_4;
output x_out_27_5;
output x_out_27_6;
output x_out_27_7;
output x_out_27_8;
output x_out_27_9;
output x_out_28_0;
output x_out_28_1;
output x_out_28_10;
output x_out_28_11;
output x_out_28_12;
output x_out_28_13;
output x_out_28_14;
output x_out_28_15;
output x_out_28_18;
output x_out_28_19;
output x_out_28_2;
output x_out_28_20;
output x_out_28_21;
output x_out_28_22;
output x_out_28_23;
output x_out_28_24;
output x_out_28_25;
output x_out_28_26;
output x_out_28_27;
output x_out_28_28;
output x_out_28_29;
output x_out_28_3;
output x_out_28_30;
output x_out_28_31;
output x_out_28_32;
output x_out_28_33;
output x_out_28_4;
output x_out_28_5;
output x_out_28_6;
output x_out_28_7;
output x_out_28_8;
output x_out_28_9;
output x_out_29_0;
output x_out_29_1;
output x_out_29_10;
output x_out_29_11;
output x_out_29_12;
output x_out_29_13;
output x_out_29_14;
output x_out_29_15;
output x_out_29_18;
output x_out_29_19;
output x_out_29_2;
output x_out_29_20;
output x_out_29_21;
output x_out_29_22;
output x_out_29_23;
output x_out_29_24;
output x_out_29_25;
output x_out_29_26;
output x_out_29_27;
output x_out_29_28;
output x_out_29_29;
output x_out_29_3;
output x_out_29_30;
output x_out_29_31;
output x_out_29_32;
output x_out_29_33;
output x_out_29_4;
output x_out_29_5;
output x_out_29_6;
output x_out_29_7;
output x_out_29_8;
output x_out_29_9;
output x_out_2_0;
output x_out_2_1;
output x_out_2_10;
output x_out_2_11;
output x_out_2_12;
output x_out_2_13;
output x_out_2_14;
output x_out_2_15;
output x_out_2_18;
output x_out_2_19;
output x_out_2_2;
output x_out_2_20;
output x_out_2_21;
output x_out_2_22;
output x_out_2_23;
output x_out_2_24;
output x_out_2_25;
output x_out_2_26;
output x_out_2_27;
output x_out_2_28;
output x_out_2_29;
output x_out_2_3;
output x_out_2_30;
output x_out_2_31;
output x_out_2_32;
output x_out_2_33;
output x_out_2_4;
output x_out_2_5;
output x_out_2_6;
output x_out_2_7;
output x_out_2_8;
output x_out_2_9;
output x_out_30_0;
output x_out_30_1;
output x_out_30_10;
output x_out_30_11;
output x_out_30_12;
output x_out_30_13;
output x_out_30_14;
output x_out_30_15;
output x_out_30_18;
output x_out_30_19;
output x_out_30_2;
output x_out_30_20;
output x_out_30_21;
output x_out_30_22;
output x_out_30_23;
output x_out_30_24;
output x_out_30_25;
output x_out_30_26;
output x_out_30_27;
output x_out_30_28;
output x_out_30_29;
output x_out_30_3;
output x_out_30_30;
output x_out_30_31;
output x_out_30_32;
output x_out_30_33;
output x_out_30_4;
output x_out_30_5;
output x_out_30_6;
output x_out_30_7;
output x_out_30_8;
output x_out_30_9;
output x_out_31_0;
output x_out_31_1;
output x_out_31_10;
output x_out_31_11;
output x_out_31_12;
output x_out_31_13;
output x_out_31_14;
output x_out_31_15;
output x_out_31_18;
output x_out_31_19;
output x_out_31_2;
output x_out_31_20;
output x_out_31_21;
output x_out_31_22;
output x_out_31_23;
output x_out_31_24;
output x_out_31_25;
output x_out_31_26;
output x_out_31_27;
output x_out_31_28;
output x_out_31_29;
output x_out_31_3;
output x_out_31_30;
output x_out_31_31;
output x_out_31_32;
output x_out_31_33;
output x_out_31_4;
output x_out_31_5;
output x_out_31_6;
output x_out_31_7;
output x_out_31_8;
output x_out_31_9;
output x_out_32_0;
output x_out_32_1;
output x_out_32_10;
output x_out_32_11;
output x_out_32_12;
output x_out_32_13;
output x_out_32_14;
output x_out_32_15;
output x_out_32_2;
output x_out_32_3;
output x_out_32_4;
output x_out_32_5;
output x_out_32_6;
output x_out_32_7;
output x_out_32_8;
output x_out_32_9;
output x_out_33_0;
output x_out_33_1;
output x_out_33_10;
output x_out_33_11;
output x_out_33_12;
output x_out_33_13;
output x_out_33_14;
output x_out_33_15;
output x_out_33_18;
output x_out_33_19;
output x_out_33_2;
output x_out_33_20;
output x_out_33_21;
output x_out_33_22;
output x_out_33_23;
output x_out_33_24;
output x_out_33_25;
output x_out_33_26;
output x_out_33_27;
output x_out_33_28;
output x_out_33_29;
output x_out_33_3;
output x_out_33_30;
output x_out_33_31;
output x_out_33_32;
output x_out_33_33;
output x_out_33_4;
output x_out_33_5;
output x_out_33_6;
output x_out_33_7;
output x_out_33_8;
output x_out_33_9;
output x_out_34_0;
output x_out_34_1;
output x_out_34_10;
output x_out_34_11;
output x_out_34_12;
output x_out_34_13;
output x_out_34_14;
output x_out_34_15;
output x_out_34_18;
output x_out_34_19;
output x_out_34_2;
output x_out_34_20;
output x_out_34_21;
output x_out_34_22;
output x_out_34_23;
output x_out_34_24;
output x_out_34_25;
output x_out_34_26;
output x_out_34_27;
output x_out_34_28;
output x_out_34_29;
output x_out_34_3;
output x_out_34_30;
output x_out_34_31;
output x_out_34_32;
output x_out_34_33;
output x_out_34_4;
output x_out_34_5;
output x_out_34_6;
output x_out_34_7;
output x_out_34_8;
output x_out_34_9;
output x_out_35_0;
output x_out_35_1;
output x_out_35_10;
output x_out_35_11;
output x_out_35_12;
output x_out_35_13;
output x_out_35_14;
output x_out_35_15;
output x_out_35_18;
output x_out_35_19;
output x_out_35_2;
output x_out_35_20;
output x_out_35_21;
output x_out_35_22;
output x_out_35_23;
output x_out_35_24;
output x_out_35_25;
output x_out_35_26;
output x_out_35_27;
output x_out_35_28;
output x_out_35_29;
output x_out_35_3;
output x_out_35_30;
output x_out_35_31;
output x_out_35_32;
output x_out_35_33;
output x_out_35_4;
output x_out_35_5;
output x_out_35_6;
output x_out_35_7;
output x_out_35_8;
output x_out_35_9;
output x_out_36_0;
output x_out_36_1;
output x_out_36_10;
output x_out_36_11;
output x_out_36_12;
output x_out_36_13;
output x_out_36_14;
output x_out_36_15;
output x_out_36_18;
output x_out_36_19;
output x_out_36_2;
output x_out_36_20;
output x_out_36_21;
output x_out_36_22;
output x_out_36_23;
output x_out_36_24;
output x_out_36_25;
output x_out_36_26;
output x_out_36_27;
output x_out_36_28;
output x_out_36_29;
output x_out_36_3;
output x_out_36_30;
output x_out_36_31;
output x_out_36_32;
output x_out_36_33;
output x_out_36_4;
output x_out_36_5;
output x_out_36_6;
output x_out_36_7;
output x_out_36_8;
output x_out_36_9;
output x_out_37_0;
output x_out_37_1;
output x_out_37_10;
output x_out_37_11;
output x_out_37_12;
output x_out_37_13;
output x_out_37_14;
output x_out_37_15;
output x_out_37_18;
output x_out_37_19;
output x_out_37_2;
output x_out_37_20;
output x_out_37_21;
output x_out_37_22;
output x_out_37_23;
output x_out_37_24;
output x_out_37_25;
output x_out_37_26;
output x_out_37_27;
output x_out_37_28;
output x_out_37_29;
output x_out_37_3;
output x_out_37_30;
output x_out_37_31;
output x_out_37_32;
output x_out_37_33;
output x_out_37_4;
output x_out_37_5;
output x_out_37_6;
output x_out_37_7;
output x_out_37_8;
output x_out_37_9;
output x_out_38_0;
output x_out_38_1;
output x_out_38_10;
output x_out_38_11;
output x_out_38_12;
output x_out_38_13;
output x_out_38_14;
output x_out_38_15;
output x_out_38_18;
output x_out_38_19;
output x_out_38_2;
output x_out_38_20;
output x_out_38_21;
output x_out_38_22;
output x_out_38_23;
output x_out_38_24;
output x_out_38_25;
output x_out_38_26;
output x_out_38_27;
output x_out_38_28;
output x_out_38_29;
output x_out_38_3;
output x_out_38_30;
output x_out_38_31;
output x_out_38_32;
output x_out_38_33;
output x_out_38_4;
output x_out_38_5;
output x_out_38_6;
output x_out_38_7;
output x_out_38_8;
output x_out_38_9;
output x_out_39_0;
output x_out_39_1;
output x_out_39_10;
output x_out_39_11;
output x_out_39_12;
output x_out_39_13;
output x_out_39_14;
output x_out_39_15;
output x_out_39_18;
output x_out_39_19;
output x_out_39_2;
output x_out_39_20;
output x_out_39_21;
output x_out_39_22;
output x_out_39_23;
output x_out_39_24;
output x_out_39_25;
output x_out_39_26;
output x_out_39_27;
output x_out_39_28;
output x_out_39_29;
output x_out_39_3;
output x_out_39_30;
output x_out_39_31;
output x_out_39_32;
output x_out_39_33;
output x_out_39_4;
output x_out_39_5;
output x_out_39_6;
output x_out_39_7;
output x_out_39_8;
output x_out_39_9;
output x_out_3_0;
output x_out_3_1;
output x_out_3_10;
output x_out_3_11;
output x_out_3_12;
output x_out_3_13;
output x_out_3_14;
output x_out_3_15;
output x_out_3_18;
output x_out_3_19;
output x_out_3_2;
output x_out_3_20;
output x_out_3_21;
output x_out_3_22;
output x_out_3_23;
output x_out_3_24;
output x_out_3_25;
output x_out_3_26;
output x_out_3_27;
output x_out_3_28;
output x_out_3_29;
output x_out_3_3;
output x_out_3_30;
output x_out_3_31;
output x_out_3_32;
output x_out_3_33;
output x_out_3_4;
output x_out_3_5;
output x_out_3_6;
output x_out_3_7;
output x_out_3_8;
output x_out_3_9;
output x_out_40_0;
output x_out_40_1;
output x_out_40_10;
output x_out_40_11;
output x_out_40_12;
output x_out_40_13;
output x_out_40_14;
output x_out_40_15;
output x_out_40_18;
output x_out_40_19;
output x_out_40_2;
output x_out_40_20;
output x_out_40_21;
output x_out_40_22;
output x_out_40_23;
output x_out_40_24;
output x_out_40_25;
output x_out_40_26;
output x_out_40_27;
output x_out_40_28;
output x_out_40_29;
output x_out_40_3;
output x_out_40_30;
output x_out_40_31;
output x_out_40_32;
output x_out_40_33;
output x_out_40_4;
output x_out_40_5;
output x_out_40_6;
output x_out_40_7;
output x_out_40_8;
output x_out_40_9;
output x_out_41_0;
output x_out_41_1;
output x_out_41_10;
output x_out_41_11;
output x_out_41_12;
output x_out_41_13;
output x_out_41_14;
output x_out_41_15;
output x_out_41_18;
output x_out_41_19;
output x_out_41_2;
output x_out_41_20;
output x_out_41_21;
output x_out_41_22;
output x_out_41_23;
output x_out_41_24;
output x_out_41_25;
output x_out_41_26;
output x_out_41_27;
output x_out_41_28;
output x_out_41_29;
output x_out_41_3;
output x_out_41_30;
output x_out_41_31;
output x_out_41_32;
output x_out_41_33;
output x_out_41_4;
output x_out_41_5;
output x_out_41_6;
output x_out_41_7;
output x_out_41_8;
output x_out_41_9;
output x_out_42_0;
output x_out_42_1;
output x_out_42_10;
output x_out_42_11;
output x_out_42_12;
output x_out_42_13;
output x_out_42_14;
output x_out_42_15;
output x_out_42_18;
output x_out_42_19;
output x_out_42_2;
output x_out_42_20;
output x_out_42_21;
output x_out_42_22;
output x_out_42_23;
output x_out_42_24;
output x_out_42_25;
output x_out_42_26;
output x_out_42_27;
output x_out_42_28;
output x_out_42_29;
output x_out_42_3;
output x_out_42_30;
output x_out_42_31;
output x_out_42_32;
output x_out_42_33;
output x_out_42_4;
output x_out_42_5;
output x_out_42_6;
output x_out_42_7;
output x_out_42_8;
output x_out_42_9;
output x_out_43_0;
output x_out_43_1;
output x_out_43_10;
output x_out_43_11;
output x_out_43_12;
output x_out_43_13;
output x_out_43_14;
output x_out_43_15;
output x_out_43_18;
output x_out_43_19;
output x_out_43_2;
output x_out_43_20;
output x_out_43_21;
output x_out_43_22;
output x_out_43_23;
output x_out_43_24;
output x_out_43_25;
output x_out_43_26;
output x_out_43_27;
output x_out_43_28;
output x_out_43_29;
output x_out_43_3;
output x_out_43_30;
output x_out_43_31;
output x_out_43_32;
output x_out_43_33;
output x_out_43_4;
output x_out_43_5;
output x_out_43_6;
output x_out_43_7;
output x_out_43_8;
output x_out_43_9;
output x_out_44_0;
output x_out_44_1;
output x_out_44_10;
output x_out_44_11;
output x_out_44_12;
output x_out_44_13;
output x_out_44_14;
output x_out_44_15;
output x_out_44_18;
output x_out_44_19;
output x_out_44_2;
output x_out_44_20;
output x_out_44_21;
output x_out_44_22;
output x_out_44_23;
output x_out_44_24;
output x_out_44_25;
output x_out_44_26;
output x_out_44_27;
output x_out_44_28;
output x_out_44_29;
output x_out_44_3;
output x_out_44_30;
output x_out_44_31;
output x_out_44_32;
output x_out_44_33;
output x_out_44_4;
output x_out_44_5;
output x_out_44_6;
output x_out_44_7;
output x_out_44_8;
output x_out_44_9;
output x_out_45_0;
output x_out_45_1;
output x_out_45_10;
output x_out_45_11;
output x_out_45_12;
output x_out_45_13;
output x_out_45_14;
output x_out_45_15;
output x_out_45_18;
output x_out_45_19;
output x_out_45_2;
output x_out_45_20;
output x_out_45_21;
output x_out_45_22;
output x_out_45_23;
output x_out_45_24;
output x_out_45_25;
output x_out_45_26;
output x_out_45_27;
output x_out_45_28;
output x_out_45_29;
output x_out_45_3;
output x_out_45_30;
output x_out_45_31;
output x_out_45_32;
output x_out_45_33;
output x_out_45_4;
output x_out_45_5;
output x_out_45_6;
output x_out_45_7;
output x_out_45_8;
output x_out_45_9;
output x_out_46_0;
output x_out_46_1;
output x_out_46_10;
output x_out_46_11;
output x_out_46_12;
output x_out_46_13;
output x_out_46_14;
output x_out_46_15;
output x_out_46_18;
output x_out_46_19;
output x_out_46_2;
output x_out_46_20;
output x_out_46_21;
output x_out_46_22;
output x_out_46_23;
output x_out_46_24;
output x_out_46_25;
output x_out_46_26;
output x_out_46_27;
output x_out_46_28;
output x_out_46_29;
output x_out_46_3;
output x_out_46_30;
output x_out_46_31;
output x_out_46_32;
output x_out_46_33;
output x_out_46_4;
output x_out_46_5;
output x_out_46_6;
output x_out_46_7;
output x_out_46_8;
output x_out_46_9;
output x_out_47_0;
output x_out_47_1;
output x_out_47_10;
output x_out_47_11;
output x_out_47_12;
output x_out_47_13;
output x_out_47_14;
output x_out_47_15;
output x_out_47_18;
output x_out_47_19;
output x_out_47_2;
output x_out_47_20;
output x_out_47_21;
output x_out_47_22;
output x_out_47_23;
output x_out_47_24;
output x_out_47_25;
output x_out_47_26;
output x_out_47_27;
output x_out_47_28;
output x_out_47_29;
output x_out_47_3;
output x_out_47_30;
output x_out_47_31;
output x_out_47_32;
output x_out_47_33;
output x_out_47_4;
output x_out_47_5;
output x_out_47_6;
output x_out_47_7;
output x_out_47_8;
output x_out_47_9;
output x_out_48_0;
output x_out_48_1;
output x_out_48_10;
output x_out_48_11;
output x_out_48_12;
output x_out_48_13;
output x_out_48_14;
output x_out_48_15;
output x_out_48_18;
output x_out_48_19;
output x_out_48_2;
output x_out_48_20;
output x_out_48_21;
output x_out_48_22;
output x_out_48_23;
output x_out_48_24;
output x_out_48_25;
output x_out_48_26;
output x_out_48_27;
output x_out_48_28;
output x_out_48_29;
output x_out_48_3;
output x_out_48_30;
output x_out_48_31;
output x_out_48_32;
output x_out_48_33;
output x_out_48_4;
output x_out_48_5;
output x_out_48_6;
output x_out_48_7;
output x_out_48_8;
output x_out_48_9;
output x_out_49_0;
output x_out_49_1;
output x_out_49_10;
output x_out_49_11;
output x_out_49_12;
output x_out_49_13;
output x_out_49_14;
output x_out_49_15;
output x_out_49_18;
output x_out_49_19;
output x_out_49_2;
output x_out_49_20;
output x_out_49_21;
output x_out_49_22;
output x_out_49_23;
output x_out_49_24;
output x_out_49_25;
output x_out_49_26;
output x_out_49_27;
output x_out_49_28;
output x_out_49_29;
output x_out_49_3;
output x_out_49_30;
output x_out_49_31;
output x_out_49_32;
output x_out_49_33;
output x_out_49_4;
output x_out_49_5;
output x_out_49_6;
output x_out_49_7;
output x_out_49_8;
output x_out_49_9;
output x_out_4_0;
output x_out_4_1;
output x_out_4_10;
output x_out_4_11;
output x_out_4_12;
output x_out_4_13;
output x_out_4_14;
output x_out_4_15;
output x_out_4_18;
output x_out_4_19;
output x_out_4_2;
output x_out_4_20;
output x_out_4_21;
output x_out_4_22;
output x_out_4_23;
output x_out_4_24;
output x_out_4_25;
output x_out_4_26;
output x_out_4_27;
output x_out_4_28;
output x_out_4_29;
output x_out_4_3;
output x_out_4_30;
output x_out_4_31;
output x_out_4_32;
output x_out_4_33;
output x_out_4_4;
output x_out_4_5;
output x_out_4_6;
output x_out_4_7;
output x_out_4_8;
output x_out_4_9;
output x_out_50_0;
output x_out_50_1;
output x_out_50_10;
output x_out_50_11;
output x_out_50_12;
output x_out_50_13;
output x_out_50_14;
output x_out_50_15;
output x_out_50_18;
output x_out_50_19;
output x_out_50_2;
output x_out_50_20;
output x_out_50_21;
output x_out_50_22;
output x_out_50_23;
output x_out_50_24;
output x_out_50_25;
output x_out_50_26;
output x_out_50_27;
output x_out_50_28;
output x_out_50_29;
output x_out_50_3;
output x_out_50_30;
output x_out_50_31;
output x_out_50_32;
output x_out_50_33;
output x_out_50_4;
output x_out_50_5;
output x_out_50_6;
output x_out_50_7;
output x_out_50_8;
output x_out_50_9;
output x_out_51_0;
output x_out_51_1;
output x_out_51_10;
output x_out_51_11;
output x_out_51_12;
output x_out_51_13;
output x_out_51_14;
output x_out_51_15;
output x_out_51_18;
output x_out_51_19;
output x_out_51_2;
output x_out_51_20;
output x_out_51_21;
output x_out_51_22;
output x_out_51_23;
output x_out_51_24;
output x_out_51_25;
output x_out_51_26;
output x_out_51_27;
output x_out_51_28;
output x_out_51_29;
output x_out_51_3;
output x_out_51_30;
output x_out_51_31;
output x_out_51_32;
output x_out_51_33;
output x_out_51_4;
output x_out_51_5;
output x_out_51_6;
output x_out_51_7;
output x_out_51_8;
output x_out_51_9;
output x_out_52_0;
output x_out_52_1;
output x_out_52_10;
output x_out_52_11;
output x_out_52_12;
output x_out_52_13;
output x_out_52_14;
output x_out_52_15;
output x_out_52_2;
output x_out_52_3;
output x_out_52_4;
output x_out_52_5;
output x_out_52_6;
output x_out_52_7;
output x_out_52_8;
output x_out_52_9;
output x_out_53_0;
output x_out_53_1;
output x_out_53_10;
output x_out_53_11;
output x_out_53_12;
output x_out_53_13;
output x_out_53_14;
output x_out_53_15;
output x_out_53_18;
output x_out_53_19;
output x_out_53_2;
output x_out_53_20;
output x_out_53_21;
output x_out_53_22;
output x_out_53_23;
output x_out_53_24;
output x_out_53_25;
output x_out_53_26;
output x_out_53_27;
output x_out_53_28;
output x_out_53_29;
output x_out_53_3;
output x_out_53_30;
output x_out_53_31;
output x_out_53_32;
output x_out_53_33;
output x_out_53_4;
output x_out_53_5;
output x_out_53_6;
output x_out_53_7;
output x_out_53_8;
output x_out_53_9;
output x_out_54_0;
output x_out_54_1;
output x_out_54_10;
output x_out_54_11;
output x_out_54_12;
output x_out_54_13;
output x_out_54_14;
output x_out_54_15;
output x_out_54_18;
output x_out_54_19;
output x_out_54_2;
output x_out_54_20;
output x_out_54_21;
output x_out_54_22;
output x_out_54_23;
output x_out_54_24;
output x_out_54_25;
output x_out_54_26;
output x_out_54_27;
output x_out_54_28;
output x_out_54_29;
output x_out_54_3;
output x_out_54_30;
output x_out_54_31;
output x_out_54_32;
output x_out_54_33;
output x_out_54_4;
output x_out_54_5;
output x_out_54_6;
output x_out_54_7;
output x_out_54_8;
output x_out_54_9;
output x_out_55_0;
output x_out_55_1;
output x_out_55_10;
output x_out_55_11;
output x_out_55_12;
output x_out_55_13;
output x_out_55_14;
output x_out_55_15;
output x_out_55_18;
output x_out_55_19;
output x_out_55_2;
output x_out_55_20;
output x_out_55_21;
output x_out_55_22;
output x_out_55_23;
output x_out_55_24;
output x_out_55_25;
output x_out_55_26;
output x_out_55_27;
output x_out_55_28;
output x_out_55_29;
output x_out_55_3;
output x_out_55_30;
output x_out_55_31;
output x_out_55_32;
output x_out_55_33;
output x_out_55_4;
output x_out_55_5;
output x_out_55_6;
output x_out_55_7;
output x_out_55_8;
output x_out_55_9;
output x_out_56_0;
output x_out_56_1;
output x_out_56_10;
output x_out_56_11;
output x_out_56_12;
output x_out_56_13;
output x_out_56_14;
output x_out_56_15;
output x_out_56_18;
output x_out_56_19;
output x_out_56_2;
output x_out_56_20;
output x_out_56_21;
output x_out_56_22;
output x_out_56_23;
output x_out_56_24;
output x_out_56_25;
output x_out_56_26;
output x_out_56_27;
output x_out_56_28;
output x_out_56_29;
output x_out_56_3;
output x_out_56_30;
output x_out_56_31;
output x_out_56_32;
output x_out_56_33;
output x_out_56_4;
output x_out_56_5;
output x_out_56_6;
output x_out_56_7;
output x_out_56_8;
output x_out_56_9;
output x_out_57_0;
output x_out_57_1;
output x_out_57_10;
output x_out_57_11;
output x_out_57_12;
output x_out_57_13;
output x_out_57_14;
output x_out_57_15;
output x_out_57_18;
output x_out_57_19;
output x_out_57_2;
output x_out_57_20;
output x_out_57_21;
output x_out_57_22;
output x_out_57_23;
output x_out_57_24;
output x_out_57_25;
output x_out_57_26;
output x_out_57_27;
output x_out_57_28;
output x_out_57_29;
output x_out_57_3;
output x_out_57_30;
output x_out_57_31;
output x_out_57_32;
output x_out_57_33;
output x_out_57_4;
output x_out_57_5;
output x_out_57_6;
output x_out_57_7;
output x_out_57_8;
output x_out_57_9;
output x_out_58_0;
output x_out_58_1;
output x_out_58_10;
output x_out_58_11;
output x_out_58_12;
output x_out_58_13;
output x_out_58_14;
output x_out_58_15;
output x_out_58_18;
output x_out_58_19;
output x_out_58_2;
output x_out_58_20;
output x_out_58_21;
output x_out_58_22;
output x_out_58_23;
output x_out_58_24;
output x_out_58_25;
output x_out_58_26;
output x_out_58_27;
output x_out_58_28;
output x_out_58_29;
output x_out_58_3;
output x_out_58_30;
output x_out_58_31;
output x_out_58_32;
output x_out_58_33;
output x_out_58_4;
output x_out_58_5;
output x_out_58_6;
output x_out_58_7;
output x_out_58_8;
output x_out_58_9;
output x_out_59_0;
output x_out_59_1;
output x_out_59_10;
output x_out_59_11;
output x_out_59_12;
output x_out_59_13;
output x_out_59_14;
output x_out_59_15;
output x_out_59_18;
output x_out_59_19;
output x_out_59_2;
output x_out_59_20;
output x_out_59_21;
output x_out_59_22;
output x_out_59_23;
output x_out_59_24;
output x_out_59_25;
output x_out_59_26;
output x_out_59_27;
output x_out_59_28;
output x_out_59_29;
output x_out_59_3;
output x_out_59_30;
output x_out_59_31;
output x_out_59_32;
output x_out_59_33;
output x_out_59_4;
output x_out_59_5;
output x_out_59_6;
output x_out_59_7;
output x_out_59_8;
output x_out_59_9;
output x_out_5_0;
output x_out_5_1;
output x_out_5_10;
output x_out_5_11;
output x_out_5_12;
output x_out_5_13;
output x_out_5_14;
output x_out_5_15;
output x_out_5_18;
output x_out_5_19;
output x_out_5_2;
output x_out_5_20;
output x_out_5_21;
output x_out_5_22;
output x_out_5_23;
output x_out_5_24;
output x_out_5_25;
output x_out_5_26;
output x_out_5_27;
output x_out_5_28;
output x_out_5_29;
output x_out_5_3;
output x_out_5_30;
output x_out_5_31;
output x_out_5_32;
output x_out_5_33;
output x_out_5_4;
output x_out_5_5;
output x_out_5_6;
output x_out_5_7;
output x_out_5_8;
output x_out_5_9;
output x_out_60_0;
output x_out_60_1;
output x_out_60_10;
output x_out_60_11;
output x_out_60_12;
output x_out_60_13;
output x_out_60_14;
output x_out_60_15;
output x_out_60_18;
output x_out_60_19;
output x_out_60_2;
output x_out_60_20;
output x_out_60_21;
output x_out_60_22;
output x_out_60_23;
output x_out_60_24;
output x_out_60_25;
output x_out_60_26;
output x_out_60_27;
output x_out_60_28;
output x_out_60_29;
output x_out_60_3;
output x_out_60_30;
output x_out_60_31;
output x_out_60_32;
output x_out_60_33;
output x_out_60_4;
output x_out_60_5;
output x_out_60_6;
output x_out_60_7;
output x_out_60_8;
output x_out_60_9;
output x_out_61_0;
output x_out_61_1;
output x_out_61_10;
output x_out_61_11;
output x_out_61_12;
output x_out_61_13;
output x_out_61_14;
output x_out_61_15;
output x_out_61_18;
output x_out_61_19;
output x_out_61_2;
output x_out_61_20;
output x_out_61_21;
output x_out_61_22;
output x_out_61_23;
output x_out_61_24;
output x_out_61_25;
output x_out_61_26;
output x_out_61_27;
output x_out_61_28;
output x_out_61_29;
output x_out_61_3;
output x_out_61_30;
output x_out_61_31;
output x_out_61_32;
output x_out_61_33;
output x_out_61_4;
output x_out_61_5;
output x_out_61_6;
output x_out_61_7;
output x_out_61_8;
output x_out_61_9;
output x_out_62_0;
output x_out_62_1;
output x_out_62_10;
output x_out_62_11;
output x_out_62_12;
output x_out_62_13;
output x_out_62_14;
output x_out_62_15;
output x_out_62_18;
output x_out_62_19;
output x_out_62_2;
output x_out_62_20;
output x_out_62_21;
output x_out_62_22;
output x_out_62_23;
output x_out_62_24;
output x_out_62_25;
output x_out_62_26;
output x_out_62_27;
output x_out_62_28;
output x_out_62_29;
output x_out_62_3;
output x_out_62_30;
output x_out_62_31;
output x_out_62_32;
output x_out_62_33;
output x_out_62_4;
output x_out_62_5;
output x_out_62_6;
output x_out_62_7;
output x_out_62_8;
output x_out_62_9;
output x_out_63_0;
output x_out_63_1;
output x_out_63_10;
output x_out_63_11;
output x_out_63_12;
output x_out_63_13;
output x_out_63_14;
output x_out_63_15;
output x_out_63_18;
output x_out_63_19;
output x_out_63_2;
output x_out_63_20;
output x_out_63_21;
output x_out_63_22;
output x_out_63_23;
output x_out_63_24;
output x_out_63_25;
output x_out_63_26;
output x_out_63_27;
output x_out_63_28;
output x_out_63_29;
output x_out_63_3;
output x_out_63_30;
output x_out_63_31;
output x_out_63_32;
output x_out_63_33;
output x_out_63_4;
output x_out_63_5;
output x_out_63_6;
output x_out_63_7;
output x_out_63_8;
output x_out_63_9;
output x_out_6_0;
output x_out_6_1;
output x_out_6_10;
output x_out_6_11;
output x_out_6_12;
output x_out_6_13;
output x_out_6_14;
output x_out_6_15;
output x_out_6_18;
output x_out_6_19;
output x_out_6_2;
output x_out_6_20;
output x_out_6_21;
output x_out_6_22;
output x_out_6_23;
output x_out_6_24;
output x_out_6_25;
output x_out_6_26;
output x_out_6_27;
output x_out_6_28;
output x_out_6_29;
output x_out_6_3;
output x_out_6_30;
output x_out_6_31;
output x_out_6_32;
output x_out_6_33;
output x_out_6_4;
output x_out_6_5;
output x_out_6_6;
output x_out_6_7;
output x_out_6_8;
output x_out_6_9;
output x_out_7_0;
output x_out_7_1;
output x_out_7_10;
output x_out_7_11;
output x_out_7_12;
output x_out_7_13;
output x_out_7_14;
output x_out_7_15;
output x_out_7_18;
output x_out_7_19;
output x_out_7_2;
output x_out_7_20;
output x_out_7_21;
output x_out_7_22;
output x_out_7_23;
output x_out_7_24;
output x_out_7_25;
output x_out_7_26;
output x_out_7_27;
output x_out_7_28;
output x_out_7_29;
output x_out_7_3;
output x_out_7_30;
output x_out_7_31;
output x_out_7_32;
output x_out_7_33;
output x_out_7_4;
output x_out_7_5;
output x_out_7_6;
output x_out_7_7;
output x_out_7_8;
output x_out_7_9;
output x_out_8_0;
output x_out_8_1;
output x_out_8_10;
output x_out_8_11;
output x_out_8_12;
output x_out_8_13;
output x_out_8_14;
output x_out_8_15;
output x_out_8_18;
output x_out_8_19;
output x_out_8_2;
output x_out_8_20;
output x_out_8_21;
output x_out_8_22;
output x_out_8_23;
output x_out_8_24;
output x_out_8_25;
output x_out_8_26;
output x_out_8_27;
output x_out_8_28;
output x_out_8_29;
output x_out_8_3;
output x_out_8_30;
output x_out_8_31;
output x_out_8_32;
output x_out_8_33;
output x_out_8_4;
output x_out_8_5;
output x_out_8_6;
output x_out_8_7;
output x_out_8_8;
output x_out_8_9;
output x_out_9_0;
output x_out_9_1;
output x_out_9_10;
output x_out_9_11;
output x_out_9_12;
output x_out_9_13;
output x_out_9_14;
output x_out_9_15;
output x_out_9_18;
output x_out_9_19;
output x_out_9_2;
output x_out_9_20;
output x_out_9_21;
output x_out_9_22;
output x_out_9_23;
output x_out_9_24;
output x_out_9_25;
output x_out_9_26;
output x_out_9_27;
output x_out_9_28;
output x_out_9_29;
output x_out_9_3;
output x_out_9_30;
output x_out_9_31;
output x_out_9_32;
output x_out_9_33;
output x_out_9_4;
output x_out_9_5;
output x_out_9_6;
output x_out_9_7;
output x_out_9_8;
output x_out_9_9;

// Start wires
wire FE_OFN0_n_17395;
wire FE_OFN1000_n_17200;
wire FE_OFN1001_n_17200;
wire FE_OFN1002_n_19855;
wire FE_OFN1003_n_19855;
wire FE_OFN1004_n_23624;
wire FE_OFN1005_n_23624;
wire FE_OFN1006_n_24950;
wire FE_OFN1007_n_24950;
wire FE_OFN1008_n_27881;
wire FE_OFN1009_n_27881;
wire FE_OFN100_n_27449;
wire FE_OFN1010_n_28328;
wire FE_OFN1011_n_28328;
wire FE_OFN1012_n_28629;
wire FE_OFN1014_n_16571;
wire FE_OFN1015_n_16571;
wire FE_OFN1016_n_17433;
wire FE_OFN1017_n_17433;
wire FE_OFN1018_n_22081;
wire FE_OFN1019_n_22081;
wire FE_OFN101_n_27449;
wire FE_OFN1020_n_28703;
wire FE_OFN1021_n_28703;
wire FE_OFN1028_n_14570;
wire FE_OFN1029_n_14570;
wire FE_OFN102_n_27449;
wire FE_OFN1030_n_19666;
wire FE_OFN1031_n_19666;
wire FE_OFN1034_n_21194;
wire FE_OFN1035_n_21194;
wire FE_OFN1036_n_26168;
wire FE_OFN1037_n_26168;
wire FE_OFN1038_n_27890;
wire FE_OFN1039_n_27890;
wire FE_OFN103_n_27449;
wire FE_OFN1044_n_26162;
wire FE_OFN1045_n_26162;
wire FE_OFN1046_n_27057;
wire FE_OFN1047_n_27057;
wire FE_OFN104_n_27449;
wire FE_OFN1054_n_25805;
wire FE_OFN1055_n_25805;
wire FE_OFN1056_n_18817;
wire FE_OFN1057_n_18817;
wire FE_OFN1058_n_18610;
wire FE_OFN1059_n_18610;
wire FE_OFN105_n_27449;
wire FE_OFN1060_n_19587;
wire FE_OFN1061_n_19587;
wire FE_OFN106_n_27449;
wire FE_OFN1073_n_6399;
wire FE_OFN107_n_27449;
wire FE_OFN1080_n_14273;
wire FE_OFN1081_n_14273;
wire FE_OFN1082_n_8877;
wire FE_OFN1083_n_8877;
wire FE_OFN1084_n_14427;
wire FE_OFN1085_n_14427;
wire FE_OFN1086_n_8974;
wire FE_OFN1087_n_8974;
wire FE_OFN1088_n_8985;
wire FE_OFN1089_n_8985;
wire FE_OFN108_n_27449;
wire FE_OFN1090_n_8621;
wire FE_OFN1091_n_8621;
wire FE_OFN109_n_27449;
wire FE_OFN10_n_29204;
wire FE_OFN1100_n_12369;
wire FE_OFN1101_n_12369;
wire FE_OFN1102_rst;
wire FE_OFN1103_rst;
wire FE_OFN1104_rst;
wire FE_OFN1105_rst;
wire FE_OFN1106_rst;
wire FE_OFN1107_rst;
wire FE_OFN1108_rst;
wire FE_OFN1109_rst;
wire FE_OFN1110_rst;
wire FE_OFN1111_rst;
wire FE_OFN1112_rst;
wire FE_OFN1113_rst;
wire FE_OFN1114_rst;
wire FE_OFN1115_rst;
wire FE_OFN1117_rst;
wire FE_OFN1118_rst;
wire FE_OFN1119_rst;
wire FE_OFN111_n_27449;
wire FE_OFN1120_rst;
wire FE_OFN1121_rst;
wire FE_OFN1122_rst;
wire FE_OFN1123_rst;
wire FE_OFN1124_rst;
wire FE_OFN1125_n_29632;
wire FE_OFN1126_n_29632;
wire FE_OFN1127_n_29567;
wire FE_OFN1128_n_29567;
wire FE_OFN1129_n_6399;
wire FE_OFN1130_n_27986;
wire FE_OFN1131_n_28629;
wire FE_OFN1132_n_28627;
wire FE_OFN1133_n_28782;
wire FE_OFN1134_n_28627;
wire FE_OFN1135_n_28794;
wire FE_OFN1136_n_28794;
wire FE_OFN1137_n_28938;
wire FE_OFN1138_n_28938;
wire FE_OFN1139_n_27012;
wire FE_OFN113_n_27449;
wire FE_OFN1140_n_27012;
wire FE_OFN1141_n_27012;
wire FE_OFN1142_n_27012;
wire FE_OFN1143_n_27012;
wire FE_OFN1144_n_27012;
wire FE_OFN1145_n_4860;
wire FE_OFN1146_n_4860;
wire FE_OFN1147_n_4860;
wire FE_OFN1148_n_6525;
wire FE_OFN1149_n_6525;
wire FE_OFN114_n_27449;
wire FE_OFN1150_n_3069;
wire FE_OFN1151_n_3069;
wire FE_OFN1152_n_3069;
wire FE_OFN1153_n_14586;
wire FE_OFN1154_n_14586;
wire FE_OFN1155_n_14586;
wire FE_OFN1156_n_26184;
wire FE_OFN1157_n_26184;
wire FE_OFN1158_n_26184;
wire FE_OFN1159_n_26184;
wire FE_OFN115_n_27449;
wire FE_OFN1160_n_26184;
wire FE_OFN1161_n_5003;
wire FE_OFN1162_n_5003;
wire FE_OFN1163_n_4162;
wire FE_OFN1164_n_4162;
wire FE_OFN1165_n_4162;
wire FE_OFN1166_n_4162;
wire FE_OFN1167_n_4162;
wire FE_OFN1168_n_4162;
wire FE_OFN1169_n_4860;
wire FE_OFN116_n_27449;
wire FE_OFN1170_n_4860;
wire FE_OFN1171_n_4860;
wire FE_OFN1172_n_4860;
wire FE_OFN1173_n_4860;
wire FE_OFN1174_n_4860;
wire FE_OFN1175_n_28597;
wire FE_OFN1176_n_28597;
wire FE_OFN1177_n_28597;
wire FE_OFN1178_n_17184;
wire FE_OFN1179_n_17184;
wire FE_OFN117_n_27449;
wire FE_OFN1180_rst;
wire FE_OFN1181_rst;
wire FE_OFN1182_rst;
wire FE_OFN1183_n_6701;
wire FE_OFN1184_n_6701;
wire FE_OFN1185_n_12201;
wire FE_OFN1186_n_12201;
wire FE_OFN1187_n_5249;
wire FE_OFN1188_n_5249;
wire FE_OFN1189_n_13090;
wire FE_OFN118_n_27449;
wire FE_OFN1190_n_13090;
wire FE_OFN1191_n_11896;
wire FE_OFN1192_n_11896;
wire FE_OFN1193_n_12908;
wire FE_OFN1194_n_12908;
wire FE_OFN1195_n_12016;
wire FE_OFN1196_n_12016;
wire FE_OFN1197_n_13003;
wire FE_OFN1198_n_13003;
wire FE_OFN1199_n_10340;
wire FE_OFN119_n_27449;
wire FE_OFN11_n_29204;
wire FE_OFN1200_n_10340;
wire FE_OFN1201_n_5312;
wire FE_OFN1202_n_5312;
wire FE_OFN1203_n_11679;
wire FE_OFN1204_n_11679;
wire FE_OFN1205_n_9308;
wire FE_OFN1206_n_9308;
wire FE_OFN1207_n_10456;
wire FE_OFN1208_n_10456;
wire FE_OFN1209_n_10458;
wire FE_OFN120_n_27449;
wire FE_OFN1210_n_10458;
wire FE_OFN1211_n_10465;
wire FE_OFN1212_n_10465;
wire FE_OFN1213_n_10469;
wire FE_OFN1214_n_10469;
wire FE_OFN1215_n_12761;
wire FE_OFN1216_n_12761;
wire FE_OFN1217_n_13369;
wire FE_OFN1218_n_13369;
wire FE_OFN1219_n_8798;
wire FE_OFN121_n_27449;
wire FE_OFN1220_n_8798;
wire FE_OFN1221_n_6089;
wire FE_OFN1222_n_6089;
wire FE_OFN1223_n_29433;
wire FE_OFN1224_n_29433;
wire FE_OFN1225_n_10183;
wire FE_OFN1226_n_10183;
wire FE_OFN1227_n_23261;
wire FE_OFN1228_n_23261;
wire FE_OFN1229_n_24166;
wire FE_OFN122_n_27449;
wire FE_OFN1230_n_24166;
wire FE_OFN1231_n_12068;
wire FE_OFN1232_n_12068;
wire FE_OFN1233_n_4979;
wire FE_OFN1234_n_4979;
wire FE_OFN1235_n_16615;
wire FE_OFN1236_n_16615;
wire FE_OFN1237_n_10491;
wire FE_OFN1238_n_10491;
wire FE_OFN1239_n_10499;
wire FE_OFN123_n_27449;
wire FE_OFN1240_n_10499;
wire FE_OFN1241_n_29553;
wire FE_OFN1242_n_29553;
wire FE_OFN1243_n_12940;
wire FE_OFN1244_n_12940;
wire FE_OFN1245_n_4900;
wire FE_OFN1246_n_4900;
wire FE_OFN1247_n_8470;
wire FE_OFN1248_n_8470;
wire FE_OFN1249_n_5334;
wire FE_OFN124_n_27449;
wire FE_OFN1250_n_5334;
wire FE_OFN1251_n_25296;
wire FE_OFN1252_n_25296;
wire FE_OFN1253_n_12186;
wire FE_OFN1254_n_12186;
wire FE_OFN1255_n_10520;
wire FE_OFN1256_n_10520;
wire FE_OFN1257_n_4905;
wire FE_OFN1258_n_4905;
wire FE_OFN1259_n_6178;
wire FE_OFN125_n_27449;
wire FE_OFN1260_n_6178;
wire FE_OFN1261_n_6197;
wire FE_OFN1262_n_6197;
wire FE_OFN1263_n_29354;
wire FE_OFN1264_n_29354;
wire FE_OFN1265_n_16620;
wire FE_OFN1266_n_16620;
wire FE_OFN1267_n_29314;
wire FE_OFN1268_n_29314;
wire FE_OFN1269_n_29015;
wire FE_OFN126_n_27449;
wire FE_OFN1270_n_29015;
wire FE_OFN1271_n_9600;
wire FE_OFN1272_n_9600;
wire FE_OFN1273_n_8977;
wire FE_OFN1274_n_8977;
wire FE_OFN1275_n_12754;
wire FE_OFN1276_n_12754;
wire FE_OFN1277_n_6116;
wire FE_OFN1278_n_6116;
wire FE_OFN1279_n_8068;
wire FE_OFN127_n_27449;
wire FE_OFN1280_n_8068;
wire FE_OFN128_n_27449;
wire FE_OFN129_n_27449;
wire FE_OFN12_n_29204;
wire FE_OFN130_n_27449;
wire FE_OFN131_n_27449;
wire FE_OFN133_n_27449;
wire FE_OFN134_n_27449;
wire FE_OFN135_n_27449;
wire FE_OFN136_n_27449;
wire FE_OFN138_n_27449;
wire FE_OFN139_n_27449;
wire FE_OFN13_n_29068;
wire FE_OFN141_n_27449;
wire FE_OFN142_n_27449;
wire FE_OFN143_n_7361;
wire FE_OFN144_n_7361;
wire FE_OFN145_n_2667;
wire FE_OFN146_n_2667;
wire FE_OFN147_n_25677;
wire FE_OFN148_n_25677;
wire FE_OFN149_n_25677;
wire FE_OFN14_n_29068;
wire FE_OFN150_n_25677;
wire FE_OFN151_n_22615;
wire FE_OFN152_n_22615;
wire FE_OFN153_n_22615;
wire FE_OFN154_n_22615;
wire FE_OFN155_n_28014;
wire FE_OFN156_n_28014;
wire FE_OFN157_n_28014;
wire FE_OFN158_n_28014;
wire FE_OFN159_n_28014;
wire FE_OFN15_n_29068;
wire FE_OFN160_n_28014;
wire FE_OFN161_n_26454;
wire FE_OFN162_n_26454;
wire FE_OFN164_n_29269;
wire FE_OFN165_n_29269;
wire FE_OFN166_n_29269;
wire FE_OFN169_n_22948;
wire FE_OFN16_n_29617;
wire FE_OFN170_n_22948;
wire FE_OFN171_n_22948;
wire FE_OFN172_n_22948;
wire FE_OFN173_n_22948;
wire FE_OFN174_n_26184;
wire FE_OFN175_n_26184;
wire FE_OFN177_n_27681;
wire FE_OFN179_n_27681;
wire FE_OFN17_n_29617;
wire FE_OFN180_n_27681;
wire FE_OFN181_n_27681;
wire FE_OFN182_n_29402;
wire FE_OFN183_n_29402;
wire FE_OFN184_n_29402;
wire FE_OFN185_n_29496;
wire FE_OFN186_n_29496;
wire FE_OFN187_n_29496;
wire FE_OFN188_n_28362;
wire FE_OFN189_n_28362;
wire FE_OFN18_n_29617;
wire FE_OFN190_n_28362;
wire FE_OFN191_n_28928;
wire FE_OFN192_n_28928;
wire FE_OFN193_n_28928;
wire FE_OFN195_n_5003;
wire FE_OFN196_n_5003;
wire FE_OFN197_n_29637;
wire FE_OFN198_n_29637;
wire FE_OFN199_n_29637;
wire FE_OFN19_n_27452;
wire FE_OFN1_n_17395;
wire FE_OFN200_n_29637;
wire FE_OFN201_n_29637;
wire FE_OFN202_n_28771;
wire FE_OFN203_n_28771;
wire FE_OFN204_n_28771;
wire FE_OFN205_n_28771;
wire FE_OFN206_n_28771;
wire FE_OFN207_n_29661;
wire FE_OFN208_n_29661;
wire FE_OFN209_n_29661;
wire FE_OFN20_n_27452;
wire FE_OFN210_n_29661;
wire FE_OFN211_n_29661;
wire FE_OFN212_n_29661;
wire FE_OFN213_n_29687;
wire FE_OFN214_n_29687;
wire FE_OFN215_n_29687;
wire FE_OFN217_n_29687;
wire FE_OFN218_n_23315;
wire FE_OFN219_n_23315;
wire FE_OFN21_n_27452;
wire FE_OFN220_n_23315;
wire FE_OFN221_n_23315;
wire FE_OFN222_n_21642;
wire FE_OFN223_n_21642;
wire FE_OFN224_n_21642;
wire FE_OFN225_n_21642;
wire FE_OFN226_n_4162;
wire FE_OFN227_n_4162;
wire FE_OFN228_n_4162;
wire FE_OFN230_n_4162;
wire FE_OFN231_n_4162;
wire FE_OFN232_n_4162;
wire FE_OFN234_n_4162;
wire FE_OFN235_n_4162;
wire FE_OFN236_n_4162;
wire FE_OFN237_n_4162;
wire FE_OFN238_n_4162;
wire FE_OFN239_n_4162;
wire FE_OFN23_n_26609;
wire FE_OFN240_n_4162;
wire FE_OFN242_n_4162;
wire FE_OFN243_n_4162;
wire FE_OFN244_n_4162;
wire FE_OFN247_n_4162;
wire FE_OFN248_n_4162;
wire FE_OFN249_n_4162;
wire FE_OFN24_n_11489;
wire FE_OFN251_n_4162;
wire FE_OFN252_n_4280;
wire FE_OFN253_n_4280;
wire FE_OFN254_n_4280;
wire FE_OFN256_n_4280;
wire FE_OFN257_n_4280;
wire FE_OFN258_n_4280;
wire FE_OFN259_n_4280;
wire FE_OFN25_n_11489;
wire FE_OFN260_n_4280;
wire FE_OFN261_n_4280;
wire FE_OFN262_n_4280;
wire FE_OFN264_n_4280;
wire FE_OFN265_n_4280;
wire FE_OFN266_n_4280;
wire FE_OFN267_n_4280;
wire FE_OFN268_n_4280;
wire FE_OFN269_n_4280;
wire FE_OFN26_n_13676;
wire FE_OFN270_n_16028;
wire FE_OFN271_n_16028;
wire FE_OFN272_n_16893;
wire FE_OFN273_n_16893;
wire FE_OFN274_n_16893;
wire FE_OFN275_n_16893;
wire FE_OFN276_n_16893;
wire FE_OFN277_n_16893;
wire FE_OFN278_n_16656;
wire FE_OFN279_n_16656;
wire FE_OFN27_n_13676;
wire FE_OFN280_n_16656;
wire FE_OFN281_n_7349;
wire FE_OFN282_n_7349;
wire FE_OFN283_n_29266;
wire FE_OFN284_n_29266;
wire FE_OFN285_n_29266;
wire FE_OFN286_n_29266;
wire FE_OFN287_n_29266;
wire FE_OFN288_n_29266;
wire FE_OFN289_n_27194;
wire FE_OFN28_n_13676;
wire FE_OFN290_n_27194;
wire FE_OFN291_n_3069;
wire FE_OFN292_n_3069;
wire FE_OFN293_n_3069;
wire FE_OFN294_n_3069;
wire FE_OFN295_n_3069;
wire FE_OFN296_n_3069;
wire FE_OFN297_n_3069;
wire FE_OFN298_n_3069;
wire FE_OFN299_n_3069;
wire FE_OFN29_n_13676;
wire FE_OFN2_n_28682;
wire FE_OFN300_n_3069;
wire FE_OFN301_n_3069;
wire FE_OFN302_n_3069;
wire FE_OFN303_n_3069;
wire FE_OFN304_n_3069;
wire FE_OFN305_n_3069;
wire FE_OFN306_n_3069;
wire FE_OFN307_n_3069;
wire FE_OFN308_n_3069;
wire FE_OFN309_n_3069;
wire FE_OFN30_n_13676;
wire FE_OFN310_n_3069;
wire FE_OFN311_n_3069;
wire FE_OFN312_n_3069;
wire FE_OFN313_n_3069;
wire FE_OFN314_n_3069;
wire FE_OFN315_n_26999;
wire FE_OFN316_n_26999;
wire FE_OFN317_n_27400;
wire FE_OFN318_n_27400;
wire FE_OFN320_n_4860;
wire FE_OFN321_n_4860;
wire FE_OFN322_n_4860;
wire FE_OFN324_n_4860;
wire FE_OFN325_n_4860;
wire FE_OFN326_n_4860;
wire FE_OFN327_n_4860;
wire FE_OFN329_n_4860;
wire FE_OFN32_n_27986;
wire FE_OFN330_n_4860;
wire FE_OFN331_n_4860;
wire FE_OFN332_n_4860;
wire FE_OFN334_n_4860;
wire FE_OFN335_n_4860;
wire FE_OFN336_n_4860;
wire FE_OFN337_n_4860;
wire FE_OFN338_n_4860;
wire FE_OFN339_n_4860;
wire FE_OFN33_n_15183;
wire FE_OFN340_n_4860;
wire FE_OFN341_n_4860;
wire FE_OFN342_n_4860;
wire FE_OFN343_n_4860;
wire FE_OFN344_n_4860;
wire FE_OFN345_n_4860;
wire FE_OFN347_n_4860;
wire FE_OFN349_n_4860;
wire FE_OFN34_n_15183;
wire FE_OFN350_n_4860;
wire FE_OFN352_n_4860;
wire FE_OFN353_n_4860;
wire FE_OFN355_n_4860;
wire FE_OFN357_n_4860;
wire FE_OFN358_n_4860;
wire FE_OFN359_n_4860;
wire FE_OFN35_n_15183;
wire FE_OFN360_n_4860;
wire FE_OFN361_n_4860;
wire FE_OFN363_n_4860;
wire FE_OFN364_n_4860;
wire FE_OFN368_n_26312;
wire FE_OFN369_n_26312;
wire FE_OFN370_n_15817;
wire FE_OFN371_n_15817;
wire FE_OFN372_n_15853;
wire FE_OFN373_n_15853;
wire FE_OFN374_n_14224;
wire FE_OFN375_n_14224;
wire FE_OFN376_n_14285;
wire FE_OFN377_n_14285;
wire FE_OFN378_n_13985;
wire FE_OFN379_n_13985;
wire FE_OFN37_n_17184;
wire FE_OFN380_n_16289;
wire FE_OFN381_n_16289;
wire FE_OFN382_n_16289;
wire FE_OFN383_n_16289;
wire FE_OFN384_n_16289;
wire FE_OFN385_n_16289;
wire FE_OFN386_n_17236;
wire FE_OFN387_n_17236;
wire FE_OFN388_n_16991;
wire FE_OFN389_n_16991;
wire FE_OFN38_n_17184;
wire FE_OFN390_n_15554;
wire FE_OFN391_n_15554;
wire FE_OFN392_n_14663;
wire FE_OFN393_n_14663;
wire FE_OFN394_n_14720;
wire FE_OFN396_n_14720;
wire FE_OFN397_n_8616;
wire FE_OFN398_n_8616;
wire FE_OFN399_n_28303;
wire FE_OFN39_n_25450;
wire FE_OFN3_n_28682;
wire FE_OFN400_n_28303;
wire FE_OFN402_n_28303;
wire FE_OFN404_n_28303;
wire FE_OFN405_n_28303;
wire FE_OFN406_n_28303;
wire FE_OFN407_n_28303;
wire FE_OFN408_n_28303;
wire FE_OFN409_n_28303;
wire FE_OFN40_n_25450;
wire FE_OFN410_n_28303;
wire FE_OFN411_n_28303;
wire FE_OFN412_n_28303;
wire FE_OFN413_n_28303;
wire FE_OFN414_n_28303;
wire FE_OFN416_n_28303;
wire FE_OFN417_n_28303;
wire FE_OFN419_n_16909;
wire FE_OFN41_n_26563;
wire FE_OFN420_n_16909;
wire FE_OFN421_n_16909;
wire FE_OFN422_n_16909;
wire FE_OFN423_n_16296;
wire FE_OFN424_n_16296;
wire FE_OFN425_n_23661;
wire FE_OFN426_n_23661;
wire FE_OFN427_n_17707;
wire FE_OFN428_n_17707;
wire FE_OFN429_n_26458;
wire FE_OFN42_n_26563;
wire FE_OFN430_n_26458;
wire FE_OFN431_n_20518;
wire FE_OFN432_n_20518;
wire FE_OFN433_n_23637;
wire FE_OFN434_n_23637;
wire FE_OFN435_n_26167;
wire FE_OFN436_n_26167;
wire FE_OFN437_n_27889;
wire FE_OFN438_n_27889;
wire FE_OFN43_n_25810;
wire FE_OFN443_n_19118;
wire FE_OFN444_n_19118;
wire FE_OFN445_n_24948;
wire FE_OFN446_n_24948;
wire FE_OFN449_n_17680;
wire FE_OFN44_n_25810;
wire FE_OFN450_n_17680;
wire FE_OFN451_n_23152;
wire FE_OFN452_n_23152;
wire FE_OFN453_n_24837;
wire FE_OFN454_n_24837;
wire FE_OFN455_n_8508;
wire FE_OFN456_n_8508;
wire FE_OFN457_n_5621;
wire FE_OFN458_n_5621;
wire FE_OFN459_n_13371;
wire FE_OFN45_n_17233;
wire FE_OFN460_n_13371;
wire FE_OFN461_n_21334;
wire FE_OFN462_n_21334;
wire FE_OFN46_n_17233;
wire FE_OFN473_n_5257;
wire FE_OFN474_n_5257;
wire FE_OFN477_n_11170;
wire FE_OFN478_n_11170;
wire FE_OFN479_n_12184;
wire FE_OFN47_n_17099;
wire FE_OFN480_n_12184;
wire FE_OFN481_n_13520;
wire FE_OFN482_n_13520;
wire FE_OFN483_n_12038;
wire FE_OFN484_n_12038;
wire FE_OFN485_n_17500;
wire FE_OFN486_n_17500;
wire FE_OFN487_n_27256;
wire FE_OFN488_n_27256;
wire FE_OFN489_n_20516;
wire FE_OFN48_n_17099;
wire FE_OFN490_n_20516;
wire FE_OFN491_n_28765;
wire FE_OFN492_n_28765;
wire FE_OFN493_n_18414;
wire FE_OFN494_n_18414;
wire FE_OFN495_n_21648;
wire FE_OFN496_n_21648;
wire FE_OFN497_n_20677;
wire FE_OFN498_n_20677;
wire FE_OFN4_n_28682;
wire FE_OFN507_n_22083;
wire FE_OFN508_n_22083;
wire FE_OFN511_n_19847;
wire FE_OFN512_n_19847;
wire FE_OFN513_n_23620;
wire FE_OFN514_n_23620;
wire FE_OFN515_n_28406;
wire FE_OFN516_n_28406;
wire FE_OFN517_n_20894;
wire FE_OFN518_n_20894;
wire FE_OFN519_n_22315;
wire FE_OFN51_n_27012;
wire FE_OFN520_n_22315;
wire FE_OFN521_n_25685;
wire FE_OFN522_n_25685;
wire FE_OFN523_n_21282;
wire FE_OFN524_n_21282;
wire FE_OFN529_n_16938;
wire FE_OFN530_n_16938;
wire FE_OFN531_n_12317;
wire FE_OFN532_n_12317;
wire FE_OFN533_n_13775;
wire FE_OFN534_n_13775;
wire FE_OFN535_n_17798;
wire FE_OFN536_n_17798;
wire FE_OFN537_n_10328;
wire FE_OFN538_n_10328;
wire FE_OFN539_n_17809;
wire FE_OFN540_n_17809;
wire FE_OFN541_n_23570;
wire FE_OFN542_n_23570;
wire FE_OFN543_n_9030;
wire FE_OFN544_n_9030;
wire FE_OFN545_n_9036;
wire FE_OFN546_n_9036;
wire FE_OFN547_n_10452;
wire FE_OFN548_n_10452;
wire FE_OFN549_n_6072;
wire FE_OFN54_n_27012;
wire FE_OFN550_n_6072;
wire FE_OFN551_n_9482;
wire FE_OFN552_n_9482;
wire FE_OFN553_n_9468;
wire FE_OFN554_n_9468;
wire FE_OFN555_n_23580;
wire FE_OFN556_n_23580;
wire FE_OFN557_n_26546;
wire FE_OFN558_n_26546;
wire FE_OFN56_n_27012;
wire FE_OFN571_n_12800;
wire FE_OFN572_n_12800;
wire FE_OFN573_n_10137;
wire FE_OFN574_n_10137;
wire FE_OFN575_n_10136;
wire FE_OFN576_n_10136;
wire FE_OFN577_n_6424;
wire FE_OFN578_n_6424;
wire FE_OFN579_n_19119;
wire FE_OFN57_n_27012;
wire FE_OFN580_n_19119;
wire FE_OFN583_n_18103;
wire FE_OFN584_n_18103;
wire FE_OFN585_n_19447;
wire FE_OFN586_n_19447;
wire FE_OFN589_n_20904;
wire FE_OFN58_n_27012;
wire FE_OFN590_n_20904;
wire FE_OFN595_n_16896;
wire FE_OFN596_n_16896;
wire FE_OFN597_n_17615;
wire FE_OFN598_n_17615;
wire FE_OFN599_n_16000;
wire FE_OFN5_n_28597;
wire FE_OFN600_n_16000;
wire FE_OFN601_n_17761;
wire FE_OFN602_n_17761;
wire FE_OFN603_n_21535;
wire FE_OFN604_n_21535;
wire FE_OFN605_n_25225;
wire FE_OFN606_n_25225;
wire FE_OFN60_n_27012;
wire FE_OFN611_n_5698;
wire FE_OFN612_n_5698;
wire FE_OFN613_n_20110;
wire FE_OFN614_n_20110;
wire FE_OFN61_n_27012;
wire FE_OFN623_n_17378;
wire FE_OFN624_n_17378;
wire FE_OFN625_n_26697;
wire FE_OFN626_n_26697;
wire FE_OFN627_n_15605;
wire FE_OFN628_n_15605;
wire FE_OFN629_n_19358;
wire FE_OFN62_n_27012;
wire FE_OFN630_n_19358;
wire FE_OFN631_n_21154;
wire FE_OFN632_n_21154;
wire FE_OFN633_n_27731;
wire FE_OFN634_n_27731;
wire FE_OFN635_n_26260;
wire FE_OFN636_n_26260;
wire FE_OFN63_n_27012;
wire FE_OFN641_n_12432;
wire FE_OFN642_n_12432;
wire FE_OFN645_n_6732;
wire FE_OFN646_n_6732;
wire FE_OFN647_n_22008;
wire FE_OFN648_n_22008;
wire FE_OFN649_n_23576;
wire FE_OFN64_n_27012;
wire FE_OFN650_n_23576;
wire FE_OFN655_n_10503;
wire FE_OFN656_n_10503;
wire FE_OFN657_n_10424;
wire FE_OFN658_n_10424;
wire FE_OFN659_n_19445;
wire FE_OFN65_n_27012;
wire FE_OFN660_n_19445;
wire FE_OFN661_n_27899;
wire FE_OFN662_n_27899;
wire FE_OFN663_n_22027;
wire FE_OFN664_n_22027;
wire FE_OFN665_n_26759;
wire FE_OFN666_n_26759;
wire FE_OFN671_n_17494;
wire FE_OFN672_n_17494;
wire FE_OFN673_n_6720;
wire FE_OFN674_n_6720;
wire FE_OFN675_n_6824;
wire FE_OFN676_n_6824;
wire FE_OFN679_n_9691;
wire FE_OFN680_n_9691;
wire FE_OFN681_n_18155;
wire FE_OFN682_n_18155;
wire FE_OFN683_n_22025;
wire FE_OFN684_n_22025;
wire FE_OFN685_n_22968;
wire FE_OFN686_n_22968;
wire FE_OFN687_n_20109;
wire FE_OFN688_n_20109;
wire FE_OFN689_n_16216;
wire FE_OFN68_n_27012;
wire FE_OFN690_n_16216;
wire FE_OFN691_n_6708;
wire FE_OFN692_n_6708;
wire FE_OFN695_n_19853;
wire FE_OFN696_n_19853;
wire FE_OFN697_n_22333;
wire FE_OFN698_n_22333;
wire FE_OFN69_n_27012;
wire FE_OFN6_n_28597;
wire FE_OFN703_n_10462;
wire FE_OFN704_n_10462;
wire FE_OFN705_n_6444;
wire FE_OFN706_n_6444;
wire FE_OFN707_n_8059;
wire FE_OFN708_n_8059;
wire FE_OFN709_n_20192;
wire FE_OFN710_n_20192;
wire FE_OFN715_n_29187;
wire FE_OFN716_n_29187;
wire FE_OFN717_n_18993;
wire FE_OFN718_n_18993;
wire FE_OFN719_n_20807;
wire FE_OFN71_n_27012;
wire FE_OFN720_n_20807;
wire FE_OFN721_n_17438;
wire FE_OFN722_n_17438;
wire FE_OFN723_n_19019;
wire FE_OFN724_n_19019;
wire FE_OFN725_n_5240;
wire FE_OFN726_n_5240;
wire FE_OFN727_n_23636;
wire FE_OFN728_n_23636;
wire FE_OFN729_n_27888;
wire FE_OFN72_n_27012;
wire FE_OFN730_n_27888;
wire FE_OFN733_n_22952;
wire FE_OFN734_n_22952;
wire FE_OFN739_n_20195;
wire FE_OFN740_n_20195;
wire FE_OFN741_n_24025;
wire FE_OFN742_n_24025;
wire FE_OFN743_n_25732;
wire FE_OFN744_n_25732;
wire FE_OFN745_n_26604;
wire FE_OFN746_n_26604;
wire FE_OFN747_n_16529;
wire FE_OFN748_n_16529;
wire FE_OFN749_n_20252;
wire FE_OFN74_n_27012;
wire FE_OFN750_n_20252;
wire FE_OFN751_n_20252;
wire FE_OFN752_n_22913;
wire FE_OFN753_n_22913;
wire FE_OFN75_n_27012;
wire FE_OFN760_n_9661;
wire FE_OFN761_n_9661;
wire FE_OFN762_n_8501;
wire FE_OFN763_n_8501;
wire FE_OFN764_n_5707;
wire FE_OFN765_n_5707;
wire FE_OFN766_n_20476;
wire FE_OFN767_n_20476;
wire FE_OFN768_n_17379;
wire FE_OFN769_n_17379;
wire FE_OFN76_n_27012;
wire FE_OFN770_n_20323;
wire FE_OFN771_n_20323;
wire FE_OFN772_n_26698;
wire FE_OFN773_n_26698;
wire FE_OFN778_n_12158;
wire FE_OFN779_n_12158;
wire FE_OFN77_n_27012;
wire FE_OFN782_n_10771;
wire FE_OFN783_n_10771;
wire FE_OFN784_n_10198;
wire FE_OFN785_n_10198;
wire FE_OFN786_n_8855;
wire FE_OFN787_n_8855;
wire FE_OFN788_n_20913;
wire FE_OFN789_n_20913;
wire FE_OFN78_n_27012;
wire FE_OFN790_n_28272;
wire FE_OFN791_n_28272;
wire FE_OFN7_n_28597;
wire FE_OFN800_n_6782;
wire FE_OFN801_n_6782;
wire FE_OFN802_n_6771;
wire FE_OFN803_n_6771;
wire FE_OFN806_n_23617;
wire FE_OFN807_n_23617;
wire FE_OFN808_n_24927;
wire FE_OFN809_n_24927;
wire FE_OFN80_n_27012;
wire FE_OFN810_n_12878;
wire FE_OFN811_n_12878;
wire FE_OFN812_n_15982;
wire FE_OFN813_n_15982;
wire FE_OFN814_n_12310;
wire FE_OFN815_n_12310;
wire FE_OFN816_n_13135;
wire FE_OFN817_n_13135;
wire FE_OFN818_n_20821;
wire FE_OFN819_n_20821;
wire FE_OFN81_n_6529;
wire FE_OFN820_n_24644;
wire FE_OFN821_n_24644;
wire FE_OFN826_n_3772;
wire FE_OFN827_n_3772;
wire FE_OFN828_n_8424;
wire FE_OFN829_n_8424;
wire FE_OFN82_n_6529;
wire FE_OFN830_n_14863;
wire FE_OFN831_n_14863;
wire FE_OFN834_n_16760;
wire FE_OFN835_n_16760;
wire FE_OFN83_n_11673;
wire FE_OFN842_n_10412;
wire FE_OFN843_n_10412;
wire FE_OFN844_n_7616;
wire FE_OFN845_n_7616;
wire FE_OFN846_n_22340;
wire FE_OFN847_n_22340;
wire FE_OFN848_n_23567;
wire FE_OFN849_n_23567;
wire FE_OFN84_n_11673;
wire FE_OFN850_n_27728;
wire FE_OFN851_n_27728;
wire FE_OFN852_n_27880;
wire FE_OFN853_n_27880;
wire FE_OFN856_n_12565;
wire FE_OFN857_n_12565;
wire FE_OFN858_n_14125;
wire FE_OFN859_n_14125;
wire FE_OFN85_n_14586;
wire FE_OFN860_n_10492;
wire FE_OFN861_n_10492;
wire FE_OFN862_n_10495;
wire FE_OFN863_n_10495;
wire FE_OFN864_n_10501;
wire FE_OFN865_n_10501;
wire FE_OFN866_n_6151;
wire FE_OFN867_n_6151;
wire FE_OFN868_n_10506;
wire FE_OFN869_n_10506;
wire FE_OFN86_n_14586;
wire FE_OFN870_n_6154;
wire FE_OFN871_n_6154;
wire FE_OFN872_n_8070;
wire FE_OFN873_n_8070;
wire FE_OFN874_n_6157;
wire FE_OFN875_n_6157;
wire FE_OFN876_n_22329;
wire FE_OFN877_n_22329;
wire FE_OFN878_n_28229;
wire FE_OFN879_n_28229;
wire FE_OFN87_n_27449;
wire FE_OFN884_n_28405;
wire FE_OFN885_n_28405;
wire FE_OFN888_n_18291;
wire FE_OFN889_n_18291;
wire FE_OFN88_n_27449;
wire FE_OFN890_n_22165;
wire FE_OFN891_n_22165;
wire FE_OFN892_n_20806;
wire FE_OFN893_n_20806;
wire FE_OFN894_n_15923;
wire FE_OFN895_n_15923;
wire FE_OFN896_n_15930;
wire FE_OFN897_n_15930;
wire FE_OFN898_n_19332;
wire FE_OFN899_n_19332;
wire FE_OFN89_n_27449;
wire FE_OFN8_n_11667;
wire FE_OFN900_n_26098;
wire FE_OFN901_n_26098;
wire FE_OFN902_n_20903;
wire FE_OFN903_n_20903;
wire FE_OFN904_n_24967;
wire FE_OFN905_n_24967;
wire FE_OFN90_n_27449;
wire FE_OFN910_n_19850;
wire FE_OFN911_n_19850;
wire FE_OFN912_n_28409;
wire FE_OFN913_n_28409;
wire FE_OFN916_n_19297;
wire FE_OFN917_n_19297;
wire FE_OFN918_n_19575;
wire FE_OFN919_n_19575;
wire FE_OFN91_n_27449;
wire FE_OFN920_n_22498;
wire FE_OFN921_n_22498;
wire FE_OFN922_n_24430;
wire FE_OFN923_n_24430;
wire FE_OFN92_n_27449;
wire FE_OFN930_n_4898;
wire FE_OFN931_n_4898;
wire FE_OFN932_n_4950;
wire FE_OFN933_n_4950;
wire FE_OFN934_n_22317;
wire FE_OFN935_n_22317;
wire FE_OFN936_n_27359;
wire FE_OFN937_n_27359;
wire FE_OFN938_n_21084;
wire FE_OFN939_n_21084;
wire FE_OFN93_n_27449;
wire FE_OFN940_n_23815;
wire FE_OFN941_n_23815;
wire FE_OFN942_n_24127;
wire FE_OFN943_n_24127;
wire FE_OFN944_n_27398;
wire FE_OFN945_n_27398;
wire FE_OFN94_n_27449;
wire FE_OFN952_n_13421;
wire FE_OFN953_n_13421;
wire FE_OFN956_n_13438;
wire FE_OFN957_n_13438;
wire FE_OFN95_n_27449;
wire FE_OFN962_n_9280;
wire FE_OFN963_n_9280;
wire FE_OFN964_n_9283;
wire FE_OFN965_n_9283;
wire FE_OFN966_n_9286;
wire FE_OFN967_n_9286;
wire FE_OFN96_n_27449;
wire FE_OFN970_n_6854;
wire FE_OFN971_n_6854;
wire FE_OFN972_n_6822;
wire FE_OFN973_n_6822;
wire FE_OFN978_n_12566;
wire FE_OFN979_n_12566;
wire FE_OFN980_n_16353;
wire FE_OFN981_n_16353;
wire FE_OFN986_n_12804;
wire FE_OFN987_n_12804;
wire FE_OFN988_n_13374;
wire FE_OFN989_n_13374;
wire FE_OFN98_n_27449;
wire FE_OFN990_n_5720;
wire FE_OFN991_n_5720;
wire FE_OFN992_n_16934;
wire FE_OFN993_n_16934;
wire FE_OFN994_n_22325;
wire FE_OFN995_n_22325;
wire FE_OFN996_n_23622;
wire FE_OFN997_n_23622;
wire FE_OFN998_n_28782;
wire FE_OFN99_n_27449;
wire FE_OFN9_n_11667;
wire ispd_clk;
wire n_0;
wire n_1;
wire n_10;
wire n_100;
wire n_1000;
wire n_10000;
wire n_10001;
wire n_10002;
wire n_10003;
wire n_10004;
wire n_10005;
wire n_10006;
wire n_10007;
wire n_10008;
wire n_10009;
wire n_1001;
wire n_10010;
wire n_10011;
wire n_10012;
wire n_10013;
wire n_10014;
wire n_10015;
wire n_10016;
wire n_10017;
wire n_10018;
wire n_10019;
wire n_1002;
wire n_10020;
wire n_10021;
wire n_10022;
wire n_10023;
wire n_10024;
wire n_10025;
wire n_10026;
wire n_10027;
wire n_10028;
wire n_10029;
wire n_1003;
wire n_10030;
wire n_10031;
wire n_10032;
wire n_10033;
wire n_10034;
wire n_10035;
wire n_10036;
wire n_10037;
wire n_10038;
wire n_10039;
wire n_1004;
wire n_10040;
wire n_10041;
wire n_10042;
wire n_10043;
wire n_10044;
wire n_10045;
wire n_10046;
wire n_10047;
wire n_10048;
wire n_10049;
wire n_1005;
wire n_10050;
wire n_10051;
wire n_10052;
wire n_10053;
wire n_10054;
wire n_10055;
wire n_10056;
wire n_10057;
wire n_10058;
wire n_10059;
wire n_1006;
wire n_10060;
wire n_10061;
wire n_10062;
wire n_10063;
wire n_10064;
wire n_10065;
wire n_10066;
wire n_10067;
wire n_10068;
wire n_10069;
wire n_1007;
wire n_10070;
wire n_10071;
wire n_10072;
wire n_10073;
wire n_10074;
wire n_10075;
wire n_10076;
wire n_10077;
wire n_10078;
wire n_10079;
wire n_1008;
wire n_10080;
wire n_10081;
wire n_10082;
wire n_10083;
wire n_10084;
wire n_10085;
wire n_10086;
wire n_10087;
wire n_10088;
wire n_10089;
wire n_1009;
wire n_10090;
wire n_10091;
wire n_10092;
wire n_10093;
wire n_10094;
wire n_10095;
wire n_10096;
wire n_10097;
wire n_10098;
wire n_10099;
wire n_101;
wire n_1010;
wire n_10100;
wire n_10101;
wire n_10102;
wire n_10103;
wire n_10104;
wire n_10105;
wire n_10106;
wire n_10107;
wire n_10108;
wire n_10109;
wire n_1011;
wire n_10110;
wire n_10111;
wire n_10112;
wire n_10113;
wire n_10114;
wire n_10115;
wire n_10116;
wire n_10117;
wire n_10118;
wire n_10119;
wire n_1012;
wire n_10120;
wire n_10121;
wire n_10122;
wire n_10123;
wire n_10124;
wire n_10125;
wire n_10126;
wire n_10127;
wire n_10128;
wire n_10129;
wire n_1013;
wire n_10130;
wire n_10131;
wire n_10132;
wire n_10133;
wire n_10134;
wire n_10135;
wire n_10136;
wire n_10137;
wire n_10138;
wire n_10139;
wire n_1014;
wire n_10140;
wire n_10141;
wire n_10142;
wire n_10143;
wire n_10144;
wire n_10145;
wire n_10146;
wire n_10147;
wire n_10148;
wire n_10149;
wire n_1015;
wire n_10150;
wire n_10151;
wire n_10152;
wire n_10153;
wire n_10154;
wire n_10155;
wire n_10156;
wire n_10157;
wire n_10158;
wire n_10159;
wire n_1016;
wire n_10160;
wire n_10161;
wire n_10162;
wire n_10163;
wire n_10164;
wire n_10165;
wire n_10166;
wire n_10167;
wire n_10168;
wire n_10169;
wire n_1017;
wire n_10170;
wire n_10171;
wire n_10172;
wire n_10173;
wire n_10174;
wire n_10175;
wire n_10176;
wire n_10177;
wire n_10178;
wire n_10179;
wire n_1018;
wire n_10180;
wire n_10181;
wire n_10182;
wire n_10183;
wire n_10184;
wire n_10185;
wire n_10186;
wire n_10187;
wire n_10188;
wire n_10189;
wire n_1019;
wire n_10190;
wire n_10191;
wire n_10192;
wire n_10193;
wire n_10194;
wire n_10195;
wire n_10196;
wire n_10197;
wire n_10198;
wire n_10199;
wire n_102;
wire n_1020;
wire n_10200;
wire n_10201;
wire n_10202;
wire n_10203;
wire n_10204;
wire n_10205;
wire n_10206;
wire n_10207;
wire n_10208;
wire n_10209;
wire n_1021;
wire n_10210;
wire n_10211;
wire n_10212;
wire n_10213;
wire n_10214;
wire n_10215;
wire n_10216;
wire n_10217;
wire n_10218;
wire n_10219;
wire n_1022;
wire n_10220;
wire n_10221;
wire n_10222;
wire n_10223;
wire n_10224;
wire n_10225;
wire n_10226;
wire n_10227;
wire n_10228;
wire n_10229;
wire n_1023;
wire n_10230;
wire n_10231;
wire n_10232;
wire n_10233;
wire n_10234;
wire n_10235;
wire n_10236;
wire n_10237;
wire n_10238;
wire n_10239;
wire n_1024;
wire n_10240;
wire n_10241;
wire n_10242;
wire n_10243;
wire n_10244;
wire n_10245;
wire n_10246;
wire n_10247;
wire n_10248;
wire n_10249;
wire n_1025;
wire n_10250;
wire n_10251;
wire n_10252;
wire n_10253;
wire n_10254;
wire n_10255;
wire n_10256;
wire n_10257;
wire n_10258;
wire n_10259;
wire n_1026;
wire n_10260;
wire n_10261;
wire n_10262;
wire n_10263;
wire n_10264;
wire n_10265;
wire n_10266;
wire n_10267;
wire n_10268;
wire n_10269;
wire n_1027;
wire n_10270;
wire n_10271;
wire n_10272;
wire n_10273;
wire n_10274;
wire n_10275;
wire n_10276;
wire n_10277;
wire n_10278;
wire n_10279;
wire n_1028;
wire n_10280;
wire n_10281;
wire n_10282;
wire n_10283;
wire n_10284;
wire n_10285;
wire n_10286;
wire n_10287;
wire n_10288;
wire n_10289;
wire n_1029;
wire n_10290;
wire n_10291;
wire n_10292;
wire n_10293;
wire n_10294;
wire n_10295;
wire n_10296;
wire n_10297;
wire n_10298;
wire n_10299;
wire n_103;
wire n_1030;
wire n_10300;
wire n_10301;
wire n_10302;
wire n_10303;
wire n_10304;
wire n_10305;
wire n_10306;
wire n_10307;
wire n_10308;
wire n_10309;
wire n_1031;
wire n_10310;
wire n_10311;
wire n_10312;
wire n_10313;
wire n_10314;
wire n_10315;
wire n_10316;
wire n_10317;
wire n_10318;
wire n_10319;
wire n_1032;
wire n_10320;
wire n_10321;
wire n_10322;
wire n_10323;
wire n_10324;
wire n_10325;
wire n_10326;
wire n_10327;
wire n_10328;
wire n_10329;
wire n_1033;
wire n_10330;
wire n_10331;
wire n_10332;
wire n_10333;
wire n_10334;
wire n_10335;
wire n_10336;
wire n_10337;
wire n_10338;
wire n_10339;
wire n_1034;
wire n_10340;
wire n_10341;
wire n_10342;
wire n_10343;
wire n_10344;
wire n_10345;
wire n_10346;
wire n_10347;
wire n_10348;
wire n_10349;
wire n_1035;
wire n_10350;
wire n_10351;
wire n_10352;
wire n_10353;
wire n_10354;
wire n_10355;
wire n_10356;
wire n_10357;
wire n_10358;
wire n_10359;
wire n_1036;
wire n_10360;
wire n_10361;
wire n_10362;
wire n_10363;
wire n_10364;
wire n_10365;
wire n_10366;
wire n_10367;
wire n_10368;
wire n_10369;
wire n_1037;
wire n_10370;
wire n_10371;
wire n_10372;
wire n_10373;
wire n_10374;
wire n_10375;
wire n_10376;
wire n_10377;
wire n_10378;
wire n_10379;
wire n_1038;
wire n_10380;
wire n_10381;
wire n_10382;
wire n_10383;
wire n_10384;
wire n_10385;
wire n_10386;
wire n_10387;
wire n_10388;
wire n_10389;
wire n_1039;
wire n_10390;
wire n_10391;
wire n_10392;
wire n_10393;
wire n_10394;
wire n_10395;
wire n_10396;
wire n_10397;
wire n_10398;
wire n_10399;
wire n_104;
wire n_1040;
wire n_10400;
wire n_10401;
wire n_10402;
wire n_10403;
wire n_10404;
wire n_10405;
wire n_10406;
wire n_10407;
wire n_10408;
wire n_10409;
wire n_1041;
wire n_10410;
wire n_10411;
wire n_10412;
wire n_10413;
wire n_10414;
wire n_10415;
wire n_10416;
wire n_10417;
wire n_10418;
wire n_10419;
wire n_1042;
wire n_10420;
wire n_10421;
wire n_10422;
wire n_10423;
wire n_10424;
wire n_10425;
wire n_10426;
wire n_10427;
wire n_10428;
wire n_10429;
wire n_1043;
wire n_10430;
wire n_10431;
wire n_10432;
wire n_10433;
wire n_10434;
wire n_10435;
wire n_10436;
wire n_10437;
wire n_10438;
wire n_10439;
wire n_1044;
wire n_10440;
wire n_10441;
wire n_10442;
wire n_10443;
wire n_10444;
wire n_10445;
wire n_10446;
wire n_10447;
wire n_10448;
wire n_10449;
wire n_1045;
wire n_10450;
wire n_10451;
wire n_10452;
wire n_10453;
wire n_10454;
wire n_10455;
wire n_10456;
wire n_10457;
wire n_10458;
wire n_10459;
wire n_1046;
wire n_10460;
wire n_10461;
wire n_10462;
wire n_10463;
wire n_10464;
wire n_10465;
wire n_10466;
wire n_10467;
wire n_10468;
wire n_10469;
wire n_1047;
wire n_10470;
wire n_10471;
wire n_10472;
wire n_10473;
wire n_10474;
wire n_10475;
wire n_10476;
wire n_10477;
wire n_10478;
wire n_10479;
wire n_1048;
wire n_10480;
wire n_10481;
wire n_10482;
wire n_10483;
wire n_10484;
wire n_10485;
wire n_10486;
wire n_10487;
wire n_10488;
wire n_10489;
wire n_1049;
wire n_10490;
wire n_10491;
wire n_10492;
wire n_10493;
wire n_10494;
wire n_10495;
wire n_10496;
wire n_10497;
wire n_10498;
wire n_10499;
wire n_105;
wire n_1050;
wire n_10500;
wire n_10501;
wire n_10502;
wire n_10503;
wire n_10504;
wire n_10505;
wire n_10506;
wire n_10507;
wire n_10508;
wire n_10509;
wire n_1051;
wire n_10510;
wire n_10511;
wire n_10512;
wire n_10513;
wire n_10514;
wire n_10515;
wire n_10516;
wire n_10517;
wire n_10518;
wire n_10519;
wire n_1052;
wire n_10520;
wire n_10521;
wire n_10522;
wire n_10523;
wire n_10524;
wire n_10525;
wire n_10526;
wire n_10527;
wire n_10528;
wire n_10529;
wire n_1053;
wire n_10530;
wire n_10531;
wire n_10532;
wire n_10533;
wire n_10534;
wire n_10535;
wire n_10536;
wire n_10537;
wire n_10538;
wire n_10539;
wire n_1054;
wire n_10540;
wire n_10541;
wire n_10542;
wire n_10543;
wire n_10544;
wire n_10545;
wire n_10546;
wire n_10547;
wire n_10548;
wire n_10549;
wire n_1055;
wire n_10550;
wire n_10551;
wire n_10552;
wire n_10553;
wire n_10554;
wire n_10555;
wire n_10556;
wire n_10557;
wire n_10558;
wire n_10559;
wire n_1056;
wire n_10560;
wire n_10561;
wire n_10562;
wire n_10563;
wire n_10564;
wire n_10565;
wire n_10566;
wire n_10567;
wire n_10568;
wire n_10569;
wire n_1057;
wire n_10570;
wire n_10571;
wire n_10572;
wire n_10573;
wire n_10574;
wire n_10575;
wire n_10576;
wire n_10577;
wire n_10578;
wire n_10579;
wire n_1058;
wire n_10580;
wire n_10581;
wire n_10582;
wire n_10583;
wire n_10584;
wire n_10585;
wire n_10586;
wire n_10587;
wire n_10588;
wire n_10589;
wire n_1059;
wire n_10590;
wire n_10591;
wire n_10592;
wire n_10593;
wire n_10594;
wire n_10595;
wire n_10596;
wire n_10597;
wire n_10598;
wire n_10599;
wire n_106;
wire n_1060;
wire n_10600;
wire n_10601;
wire n_10602;
wire n_10603;
wire n_10604;
wire n_10605;
wire n_10606;
wire n_10607;
wire n_10608;
wire n_1061;
wire n_10610;
wire n_10611;
wire n_10612;
wire n_10613;
wire n_10614;
wire n_10615;
wire n_10616;
wire n_10617;
wire n_10618;
wire n_10619;
wire n_1062;
wire n_10620;
wire n_10621;
wire n_10622;
wire n_10623;
wire n_10624;
wire n_10625;
wire n_10626;
wire n_10627;
wire n_10628;
wire n_10629;
wire n_1063;
wire n_10630;
wire n_10631;
wire n_10632;
wire n_10633;
wire n_10634;
wire n_10635;
wire n_10636;
wire n_10637;
wire n_10638;
wire n_10639;
wire n_1064;
wire n_10640;
wire n_10641;
wire n_10642;
wire n_10643;
wire n_10644;
wire n_10645;
wire n_10646;
wire n_10647;
wire n_10648;
wire n_10649;
wire n_1065;
wire n_10650;
wire n_10651;
wire n_10652;
wire n_10653;
wire n_10654;
wire n_10655;
wire n_10656;
wire n_10657;
wire n_10658;
wire n_10659;
wire n_1066;
wire n_10660;
wire n_10661;
wire n_10662;
wire n_10663;
wire n_10664;
wire n_10665;
wire n_10666;
wire n_10667;
wire n_10668;
wire n_10669;
wire n_1067;
wire n_10670;
wire n_10671;
wire n_10672;
wire n_10673;
wire n_10674;
wire n_10675;
wire n_10676;
wire n_10677;
wire n_10678;
wire n_10679;
wire n_1068;
wire n_10680;
wire n_10681;
wire n_10682;
wire n_10683;
wire n_10684;
wire n_10685;
wire n_10686;
wire n_10687;
wire n_10688;
wire n_10689;
wire n_1069;
wire n_10690;
wire n_10691;
wire n_10692;
wire n_10693;
wire n_10694;
wire n_10695;
wire n_10696;
wire n_10697;
wire n_10698;
wire n_10699;
wire n_107;
wire n_1070;
wire n_10700;
wire n_10701;
wire n_10702;
wire n_10703;
wire n_10704;
wire n_10705;
wire n_10706;
wire n_10707;
wire n_10708;
wire n_10709;
wire n_1071;
wire n_10710;
wire n_10711;
wire n_10712;
wire n_10713;
wire n_10714;
wire n_10715;
wire n_10716;
wire n_10717;
wire n_10718;
wire n_10719;
wire n_1072;
wire n_10720;
wire n_10721;
wire n_10722;
wire n_10723;
wire n_10724;
wire n_10725;
wire n_10726;
wire n_10727;
wire n_10728;
wire n_10729;
wire n_1073;
wire n_10730;
wire n_10731;
wire n_10732;
wire n_10733;
wire n_10734;
wire n_10735;
wire n_10736;
wire n_10737;
wire n_10738;
wire n_10739;
wire n_1074;
wire n_10740;
wire n_10741;
wire n_10742;
wire n_10743;
wire n_10744;
wire n_10745;
wire n_10746;
wire n_10747;
wire n_10748;
wire n_10749;
wire n_1075;
wire n_10750;
wire n_10751;
wire n_10752;
wire n_10753;
wire n_10754;
wire n_10755;
wire n_10756;
wire n_10757;
wire n_10758;
wire n_10759;
wire n_1076;
wire n_10760;
wire n_10761;
wire n_10762;
wire n_10763;
wire n_10764;
wire n_10765;
wire n_10766;
wire n_10767;
wire n_10768;
wire n_10769;
wire n_1077;
wire n_10770;
wire n_10771;
wire n_10772;
wire n_10773;
wire n_10774;
wire n_10775;
wire n_10776;
wire n_10777;
wire n_10778;
wire n_10779;
wire n_1078;
wire n_10780;
wire n_10781;
wire n_10782;
wire n_10783;
wire n_10784;
wire n_10785;
wire n_10786;
wire n_10787;
wire n_10788;
wire n_10789;
wire n_1079;
wire n_10790;
wire n_10791;
wire n_10792;
wire n_10793;
wire n_10794;
wire n_10795;
wire n_10796;
wire n_10797;
wire n_10798;
wire n_10799;
wire n_108;
wire n_1080;
wire n_10800;
wire n_10801;
wire n_10802;
wire n_10803;
wire n_10804;
wire n_10805;
wire n_10806;
wire n_10807;
wire n_10808;
wire n_10809;
wire n_1081;
wire n_10810;
wire n_10811;
wire n_10812;
wire n_10813;
wire n_10814;
wire n_10815;
wire n_10816;
wire n_10817;
wire n_10818;
wire n_10819;
wire n_1082;
wire n_10820;
wire n_10821;
wire n_10822;
wire n_10823;
wire n_10824;
wire n_10825;
wire n_10826;
wire n_10827;
wire n_10828;
wire n_10829;
wire n_1083;
wire n_10830;
wire n_10831;
wire n_10832;
wire n_10833;
wire n_10834;
wire n_10835;
wire n_10836;
wire n_10837;
wire n_10838;
wire n_10839;
wire n_1084;
wire n_10840;
wire n_10841;
wire n_10842;
wire n_10843;
wire n_10844;
wire n_10845;
wire n_10846;
wire n_10847;
wire n_10848;
wire n_10849;
wire n_1085;
wire n_10850;
wire n_10851;
wire n_10852;
wire n_10853;
wire n_10854;
wire n_10855;
wire n_10856;
wire n_10857;
wire n_10858;
wire n_10859;
wire n_1086;
wire n_10860;
wire n_10861;
wire n_10862;
wire n_10863;
wire n_10864;
wire n_10865;
wire n_10866;
wire n_10867;
wire n_10868;
wire n_10869;
wire n_1087;
wire n_10870;
wire n_10871;
wire n_10872;
wire n_10873;
wire n_10874;
wire n_10875;
wire n_10876;
wire n_10877;
wire n_10878;
wire n_10879;
wire n_1088;
wire n_10880;
wire n_10881;
wire n_10882;
wire n_10883;
wire n_10884;
wire n_10885;
wire n_10886;
wire n_10887;
wire n_10888;
wire n_10889;
wire n_1089;
wire n_10890;
wire n_10891;
wire n_10892;
wire n_10893;
wire n_10894;
wire n_10895;
wire n_10896;
wire n_10897;
wire n_10898;
wire n_10899;
wire n_109;
wire n_1090;
wire n_10900;
wire n_10901;
wire n_10902;
wire n_10903;
wire n_10904;
wire n_10905;
wire n_10906;
wire n_10907;
wire n_10908;
wire n_10909;
wire n_1091;
wire n_10910;
wire n_10911;
wire n_10912;
wire n_10913;
wire n_10914;
wire n_10915;
wire n_10916;
wire n_10917;
wire n_10918;
wire n_10919;
wire n_1092;
wire n_10920;
wire n_10921;
wire n_10922;
wire n_10923;
wire n_10924;
wire n_10925;
wire n_10926;
wire n_10927;
wire n_10928;
wire n_10929;
wire n_1093;
wire n_10930;
wire n_10931;
wire n_10932;
wire n_10933;
wire n_10934;
wire n_10935;
wire n_10936;
wire n_10937;
wire n_10938;
wire n_10939;
wire n_1094;
wire n_10940;
wire n_10941;
wire n_10942;
wire n_10943;
wire n_10944;
wire n_10945;
wire n_10946;
wire n_10947;
wire n_10948;
wire n_10949;
wire n_1095;
wire n_10950;
wire n_10951;
wire n_10952;
wire n_10953;
wire n_10954;
wire n_10955;
wire n_10956;
wire n_10957;
wire n_10958;
wire n_10959;
wire n_1096;
wire n_10960;
wire n_10961;
wire n_10962;
wire n_10963;
wire n_10964;
wire n_10965;
wire n_10966;
wire n_10967;
wire n_10968;
wire n_10969;
wire n_1097;
wire n_10970;
wire n_10971;
wire n_10972;
wire n_10973;
wire n_10974;
wire n_10975;
wire n_10976;
wire n_10977;
wire n_10978;
wire n_10979;
wire n_1098;
wire n_10980;
wire n_10981;
wire n_10982;
wire n_10983;
wire n_10984;
wire n_10985;
wire n_10986;
wire n_10987;
wire n_10988;
wire n_10989;
wire n_1099;
wire n_10990;
wire n_10991;
wire n_10992;
wire n_10993;
wire n_10994;
wire n_10995;
wire n_10996;
wire n_10997;
wire n_10998;
wire n_10999;
wire n_11;
wire n_110;
wire n_1100;
wire n_11000;
wire n_11001;
wire n_11002;
wire n_11003;
wire n_11004;
wire n_11005;
wire n_11006;
wire n_11007;
wire n_11008;
wire n_11009;
wire n_1101;
wire n_11010;
wire n_11011;
wire n_11012;
wire n_11013;
wire n_11014;
wire n_11015;
wire n_11016;
wire n_11017;
wire n_11018;
wire n_11019;
wire n_1102;
wire n_11020;
wire n_11021;
wire n_11022;
wire n_11023;
wire n_11024;
wire n_11025;
wire n_11026;
wire n_11027;
wire n_11028;
wire n_11029;
wire n_1103;
wire n_11030;
wire n_11031;
wire n_11032;
wire n_11033;
wire n_11034;
wire n_11035;
wire n_11036;
wire n_11037;
wire n_11038;
wire n_11039;
wire n_1104;
wire n_11040;
wire n_11041;
wire n_11042;
wire n_11043;
wire n_11044;
wire n_11045;
wire n_11046;
wire n_11047;
wire n_11048;
wire n_11049;
wire n_1105;
wire n_11050;
wire n_11051;
wire n_11052;
wire n_11053;
wire n_11054;
wire n_11055;
wire n_11056;
wire n_11057;
wire n_11058;
wire n_11059;
wire n_1106;
wire n_11060;
wire n_11061;
wire n_11062;
wire n_11063;
wire n_11064;
wire n_11065;
wire n_11066;
wire n_11067;
wire n_11068;
wire n_11069;
wire n_1107;
wire n_11070;
wire n_11071;
wire n_11072;
wire n_11073;
wire n_11074;
wire n_11075;
wire n_11076;
wire n_11077;
wire n_11078;
wire n_11079;
wire n_1108;
wire n_11080;
wire n_11081;
wire n_11082;
wire n_11083;
wire n_11084;
wire n_11085;
wire n_11086;
wire n_11087;
wire n_11088;
wire n_11089;
wire n_1109;
wire n_11090;
wire n_11091;
wire n_11092;
wire n_11093;
wire n_11094;
wire n_11095;
wire n_11096;
wire n_11097;
wire n_11098;
wire n_11099;
wire n_111;
wire n_1110;
wire n_11100;
wire n_11101;
wire n_11102;
wire n_11103;
wire n_11104;
wire n_11105;
wire n_11106;
wire n_11107;
wire n_11108;
wire n_11109;
wire n_1111;
wire n_11110;
wire n_11111;
wire n_11112;
wire n_11113;
wire n_11114;
wire n_11115;
wire n_11116;
wire n_11117;
wire n_11118;
wire n_11119;
wire n_1112;
wire n_11120;
wire n_11121;
wire n_11122;
wire n_11123;
wire n_11124;
wire n_11125;
wire n_11126;
wire n_11127;
wire n_11128;
wire n_11129;
wire n_1113;
wire n_11130;
wire n_11131;
wire n_11132;
wire n_11133;
wire n_11134;
wire n_11135;
wire n_11136;
wire n_11137;
wire n_11138;
wire n_11139;
wire n_1114;
wire n_11140;
wire n_11141;
wire n_11142;
wire n_11143;
wire n_11144;
wire n_11145;
wire n_11146;
wire n_11147;
wire n_11148;
wire n_11149;
wire n_1115;
wire n_11150;
wire n_11151;
wire n_11152;
wire n_11153;
wire n_11154;
wire n_11155;
wire n_11156;
wire n_11157;
wire n_11158;
wire n_11159;
wire n_1116;
wire n_11160;
wire n_11161;
wire n_11162;
wire n_11163;
wire n_11164;
wire n_11165;
wire n_11166;
wire n_11167;
wire n_11168;
wire n_11169;
wire n_1117;
wire n_11170;
wire n_11171;
wire n_11172;
wire n_11173;
wire n_11174;
wire n_11175;
wire n_11176;
wire n_11177;
wire n_11178;
wire n_11179;
wire n_1118;
wire n_11180;
wire n_11181;
wire n_11182;
wire n_11183;
wire n_11184;
wire n_11185;
wire n_11186;
wire n_11187;
wire n_11188;
wire n_11189;
wire n_1119;
wire n_11190;
wire n_11191;
wire n_11192;
wire n_11193;
wire n_11194;
wire n_11195;
wire n_11196;
wire n_11197;
wire n_11198;
wire n_11199;
wire n_112;
wire n_1120;
wire n_11200;
wire n_11201;
wire n_11202;
wire n_11203;
wire n_11204;
wire n_11205;
wire n_11206;
wire n_11207;
wire n_11208;
wire n_11209;
wire n_1121;
wire n_11210;
wire n_11211;
wire n_11212;
wire n_11213;
wire n_11214;
wire n_11215;
wire n_11216;
wire n_11217;
wire n_11218;
wire n_11219;
wire n_1122;
wire n_11220;
wire n_11221;
wire n_11222;
wire n_11223;
wire n_11224;
wire n_11225;
wire n_11226;
wire n_11227;
wire n_11228;
wire n_11229;
wire n_1123;
wire n_11230;
wire n_11231;
wire n_11232;
wire n_11233;
wire n_11234;
wire n_11235;
wire n_11236;
wire n_11237;
wire n_11238;
wire n_11239;
wire n_1124;
wire n_11240;
wire n_11241;
wire n_11242;
wire n_11243;
wire n_11244;
wire n_11245;
wire n_11246;
wire n_11247;
wire n_11248;
wire n_11249;
wire n_1125;
wire n_11250;
wire n_11251;
wire n_11252;
wire n_11253;
wire n_11254;
wire n_11255;
wire n_11256;
wire n_11257;
wire n_11258;
wire n_11259;
wire n_1126;
wire n_11260;
wire n_11261;
wire n_11262;
wire n_11263;
wire n_11264;
wire n_11265;
wire n_11266;
wire n_11267;
wire n_11268;
wire n_11269;
wire n_1127;
wire n_11270;
wire n_11271;
wire n_11272;
wire n_11273;
wire n_11274;
wire n_11275;
wire n_11276;
wire n_11277;
wire n_11278;
wire n_11279;
wire n_1128;
wire n_11280;
wire n_11281;
wire n_11282;
wire n_11283;
wire n_11284;
wire n_11285;
wire n_11286;
wire n_11287;
wire n_11288;
wire n_11289;
wire n_1129;
wire n_11290;
wire n_11291;
wire n_11292;
wire n_11293;
wire n_11294;
wire n_11295;
wire n_11296;
wire n_11297;
wire n_11298;
wire n_11299;
wire n_113;
wire n_1130;
wire n_11300;
wire n_11301;
wire n_11302;
wire n_11303;
wire n_11304;
wire n_11305;
wire n_11306;
wire n_11307;
wire n_11308;
wire n_11309;
wire n_1131;
wire n_11310;
wire n_11311;
wire n_11312;
wire n_11313;
wire n_11314;
wire n_11315;
wire n_11316;
wire n_11317;
wire n_11318;
wire n_11319;
wire n_1132;
wire n_11320;
wire n_11321;
wire n_11322;
wire n_11323;
wire n_11324;
wire n_11325;
wire n_11326;
wire n_11327;
wire n_11328;
wire n_11329;
wire n_1133;
wire n_11330;
wire n_11331;
wire n_11332;
wire n_11333;
wire n_11334;
wire n_11335;
wire n_11336;
wire n_11337;
wire n_11338;
wire n_11339;
wire n_1134;
wire n_11340;
wire n_11341;
wire n_11342;
wire n_11343;
wire n_11344;
wire n_11345;
wire n_11346;
wire n_11347;
wire n_11348;
wire n_11349;
wire n_1135;
wire n_11350;
wire n_11351;
wire n_11352;
wire n_11353;
wire n_11354;
wire n_11355;
wire n_11356;
wire n_11357;
wire n_11358;
wire n_11359;
wire n_1136;
wire n_11360;
wire n_11361;
wire n_11362;
wire n_11363;
wire n_11364;
wire n_11365;
wire n_11366;
wire n_11367;
wire n_11368;
wire n_11369;
wire n_1137;
wire n_11370;
wire n_11371;
wire n_11372;
wire n_11373;
wire n_11374;
wire n_11375;
wire n_11376;
wire n_11377;
wire n_11378;
wire n_11379;
wire n_1138;
wire n_11380;
wire n_11381;
wire n_11382;
wire n_11383;
wire n_11384;
wire n_11385;
wire n_11386;
wire n_11387;
wire n_11388;
wire n_11389;
wire n_1139;
wire n_11390;
wire n_11391;
wire n_11392;
wire n_11393;
wire n_11394;
wire n_11395;
wire n_11396;
wire n_11397;
wire n_11398;
wire n_11399;
wire n_114;
wire n_1140;
wire n_11400;
wire n_11401;
wire n_11402;
wire n_11403;
wire n_11404;
wire n_11405;
wire n_11406;
wire n_11407;
wire n_11408;
wire n_11409;
wire n_1141;
wire n_11410;
wire n_11411;
wire n_11412;
wire n_11413;
wire n_11414;
wire n_11415;
wire n_11416;
wire n_11417;
wire n_11418;
wire n_11419;
wire n_1142;
wire n_11420;
wire n_11421;
wire n_11422;
wire n_11423;
wire n_11424;
wire n_11425;
wire n_11426;
wire n_11427;
wire n_11428;
wire n_11429;
wire n_1143;
wire n_11430;
wire n_11431;
wire n_11432;
wire n_11433;
wire n_11434;
wire n_11435;
wire n_11436;
wire n_11437;
wire n_11438;
wire n_11439;
wire n_1144;
wire n_11440;
wire n_11441;
wire n_11442;
wire n_11443;
wire n_11444;
wire n_11445;
wire n_11446;
wire n_11447;
wire n_11448;
wire n_11449;
wire n_1145;
wire n_11450;
wire n_11451;
wire n_11452;
wire n_11453;
wire n_11454;
wire n_11455;
wire n_11456;
wire n_11457;
wire n_11458;
wire n_11459;
wire n_1146;
wire n_11460;
wire n_11461;
wire n_11462;
wire n_11463;
wire n_11464;
wire n_11465;
wire n_11466;
wire n_11467;
wire n_11468;
wire n_11469;
wire n_1147;
wire n_11470;
wire n_11471;
wire n_11472;
wire n_11473;
wire n_11474;
wire n_11475;
wire n_11476;
wire n_11477;
wire n_11478;
wire n_11479;
wire n_1148;
wire n_11480;
wire n_11481;
wire n_11482;
wire n_11483;
wire n_11484;
wire n_11485;
wire n_11486;
wire n_11487;
wire n_11488;
wire n_11489;
wire n_1149;
wire n_11490;
wire n_11491;
wire n_11492;
wire n_11493;
wire n_11494;
wire n_11495;
wire n_11496;
wire n_11497;
wire n_11498;
wire n_11499;
wire n_115;
wire n_1150;
wire n_11500;
wire n_11501;
wire n_11502;
wire n_11503;
wire n_11504;
wire n_11505;
wire n_11506;
wire n_11507;
wire n_11508;
wire n_11509;
wire n_1151;
wire n_11510;
wire n_11511;
wire n_11512;
wire n_11513;
wire n_11514;
wire n_11515;
wire n_11516;
wire n_11517;
wire n_11518;
wire n_11519;
wire n_1152;
wire n_11520;
wire n_11521;
wire n_11522;
wire n_11523;
wire n_11524;
wire n_11525;
wire n_11526;
wire n_11527;
wire n_11528;
wire n_11529;
wire n_1153;
wire n_11530;
wire n_11531;
wire n_11532;
wire n_11533;
wire n_11534;
wire n_11535;
wire n_11536;
wire n_11537;
wire n_11538;
wire n_11539;
wire n_1154;
wire n_11540;
wire n_11541;
wire n_11542;
wire n_11543;
wire n_11544;
wire n_11545;
wire n_11546;
wire n_11547;
wire n_11548;
wire n_11549;
wire n_1155;
wire n_11550;
wire n_11551;
wire n_11552;
wire n_11553;
wire n_11554;
wire n_11555;
wire n_11556;
wire n_11557;
wire n_11558;
wire n_11559;
wire n_1156;
wire n_11560;
wire n_11561;
wire n_11562;
wire n_11563;
wire n_11564;
wire n_11565;
wire n_11566;
wire n_11567;
wire n_11568;
wire n_11569;
wire n_1157;
wire n_11570;
wire n_11571;
wire n_11572;
wire n_11573;
wire n_11574;
wire n_11575;
wire n_11576;
wire n_11577;
wire n_11578;
wire n_11579;
wire n_1158;
wire n_11580;
wire n_11581;
wire n_11582;
wire n_11583;
wire n_11584;
wire n_11585;
wire n_11586;
wire n_11587;
wire n_11588;
wire n_11589;
wire n_1159;
wire n_11590;
wire n_11591;
wire n_11592;
wire n_11593;
wire n_11594;
wire n_11595;
wire n_11596;
wire n_11597;
wire n_11598;
wire n_11599;
wire n_116;
wire n_1160;
wire n_11600;
wire n_11601;
wire n_11602;
wire n_11603;
wire n_11604;
wire n_11605;
wire n_11606;
wire n_11607;
wire n_11608;
wire n_11609;
wire n_1161;
wire n_11610;
wire n_11611;
wire n_11612;
wire n_11613;
wire n_11614;
wire n_11615;
wire n_11616;
wire n_11617;
wire n_11618;
wire n_11619;
wire n_1162;
wire n_11620;
wire n_11621;
wire n_11622;
wire n_11623;
wire n_11624;
wire n_11625;
wire n_11626;
wire n_11627;
wire n_11628;
wire n_11629;
wire n_1163;
wire n_11630;
wire n_11631;
wire n_11632;
wire n_11633;
wire n_11634;
wire n_11635;
wire n_11636;
wire n_11637;
wire n_11638;
wire n_11639;
wire n_1164;
wire n_11640;
wire n_11641;
wire n_11642;
wire n_11643;
wire n_11644;
wire n_11645;
wire n_11646;
wire n_11647;
wire n_11648;
wire n_11649;
wire n_1165;
wire n_11650;
wire n_11651;
wire n_11652;
wire n_11653;
wire n_11654;
wire n_11655;
wire n_11656;
wire n_11657;
wire n_11658;
wire n_11659;
wire n_1166;
wire n_11660;
wire n_11661;
wire n_11662;
wire n_11663;
wire n_11664;
wire n_11665;
wire n_11666;
wire n_11667;
wire n_11668;
wire n_11669;
wire n_1167;
wire n_11670;
wire n_11671;
wire n_11672;
wire n_11673;
wire n_11674;
wire n_11675;
wire n_11676;
wire n_11677;
wire n_11678;
wire n_11679;
wire n_1168;
wire n_11680;
wire n_11681;
wire n_11682;
wire n_11683;
wire n_11684;
wire n_11685;
wire n_11686;
wire n_11687;
wire n_11688;
wire n_11689;
wire n_1169;
wire n_11690;
wire n_11691;
wire n_11692;
wire n_11693;
wire n_11694;
wire n_11695;
wire n_11696;
wire n_11697;
wire n_11698;
wire n_11699;
wire n_117;
wire n_1170;
wire n_11700;
wire n_11701;
wire n_11702;
wire n_11703;
wire n_11704;
wire n_11705;
wire n_11706;
wire n_11707;
wire n_11708;
wire n_11709;
wire n_1171;
wire n_11710;
wire n_11711;
wire n_11712;
wire n_11713;
wire n_11714;
wire n_11715;
wire n_11716;
wire n_11717;
wire n_11718;
wire n_11719;
wire n_1172;
wire n_11720;
wire n_11721;
wire n_11722;
wire n_11723;
wire n_11724;
wire n_11725;
wire n_11726;
wire n_11727;
wire n_11728;
wire n_11729;
wire n_1173;
wire n_11730;
wire n_11731;
wire n_11732;
wire n_11733;
wire n_11734;
wire n_11735;
wire n_11736;
wire n_11737;
wire n_11738;
wire n_11739;
wire n_1174;
wire n_11740;
wire n_11741;
wire n_11742;
wire n_11743;
wire n_11744;
wire n_11745;
wire n_11746;
wire n_11747;
wire n_11748;
wire n_11749;
wire n_1175;
wire n_11750;
wire n_11751;
wire n_11752;
wire n_11753;
wire n_11754;
wire n_11755;
wire n_11756;
wire n_11757;
wire n_11758;
wire n_11759;
wire n_1176;
wire n_11760;
wire n_11761;
wire n_11762;
wire n_11763;
wire n_11764;
wire n_11765;
wire n_11766;
wire n_11767;
wire n_11768;
wire n_11769;
wire n_1177;
wire n_11770;
wire n_11771;
wire n_11772;
wire n_11773;
wire n_11774;
wire n_11775;
wire n_11776;
wire n_11777;
wire n_11778;
wire n_11779;
wire n_1178;
wire n_11780;
wire n_11781;
wire n_11782;
wire n_11783;
wire n_11784;
wire n_11785;
wire n_11786;
wire n_11787;
wire n_11788;
wire n_11789;
wire n_1179;
wire n_11790;
wire n_11791;
wire n_11792;
wire n_11793;
wire n_11794;
wire n_11795;
wire n_11796;
wire n_11797;
wire n_11798;
wire n_11799;
wire n_118;
wire n_1180;
wire n_11800;
wire n_11801;
wire n_11802;
wire n_11803;
wire n_11804;
wire n_11805;
wire n_11806;
wire n_11807;
wire n_11808;
wire n_11809;
wire n_1181;
wire n_11810;
wire n_11811;
wire n_11812;
wire n_11813;
wire n_11814;
wire n_11815;
wire n_11816;
wire n_11817;
wire n_11818;
wire n_11819;
wire n_1182;
wire n_11820;
wire n_11821;
wire n_11822;
wire n_11823;
wire n_11824;
wire n_11825;
wire n_11826;
wire n_11827;
wire n_11828;
wire n_11829;
wire n_1183;
wire n_11830;
wire n_11831;
wire n_11832;
wire n_11833;
wire n_11834;
wire n_11835;
wire n_11836;
wire n_11837;
wire n_11838;
wire n_11839;
wire n_1184;
wire n_11840;
wire n_11841;
wire n_11842;
wire n_11843;
wire n_11844;
wire n_11845;
wire n_11846;
wire n_11847;
wire n_11848;
wire n_11849;
wire n_1185;
wire n_11850;
wire n_11851;
wire n_11852;
wire n_11853;
wire n_11854;
wire n_11855;
wire n_11856;
wire n_11857;
wire n_11858;
wire n_11859;
wire n_1186;
wire n_11860;
wire n_11861;
wire n_11862;
wire n_11863;
wire n_11864;
wire n_11865;
wire n_11866;
wire n_11867;
wire n_11868;
wire n_11869;
wire n_1187;
wire n_11870;
wire n_11871;
wire n_11872;
wire n_11873;
wire n_11874;
wire n_11875;
wire n_11876;
wire n_11877;
wire n_11878;
wire n_11879;
wire n_1188;
wire n_11880;
wire n_11881;
wire n_11882;
wire n_11883;
wire n_11884;
wire n_11885;
wire n_11886;
wire n_11887;
wire n_11888;
wire n_11889;
wire n_1189;
wire n_11890;
wire n_11891;
wire n_11892;
wire n_11893;
wire n_11894;
wire n_11895;
wire n_11896;
wire n_11897;
wire n_11898;
wire n_11899;
wire n_119;
wire n_1190;
wire n_11900;
wire n_11901;
wire n_11902;
wire n_11903;
wire n_11904;
wire n_11905;
wire n_11906;
wire n_11907;
wire n_11908;
wire n_11909;
wire n_1191;
wire n_11910;
wire n_11911;
wire n_11912;
wire n_11913;
wire n_11914;
wire n_11915;
wire n_11916;
wire n_11917;
wire n_11918;
wire n_11919;
wire n_1192;
wire n_11920;
wire n_11921;
wire n_11922;
wire n_11923;
wire n_11924;
wire n_11925;
wire n_11926;
wire n_11927;
wire n_11928;
wire n_11929;
wire n_1193;
wire n_11930;
wire n_11931;
wire n_11932;
wire n_11933;
wire n_11934;
wire n_11935;
wire n_11936;
wire n_11937;
wire n_11938;
wire n_11939;
wire n_1194;
wire n_11940;
wire n_11941;
wire n_11942;
wire n_11943;
wire n_11944;
wire n_11945;
wire n_11946;
wire n_11947;
wire n_11948;
wire n_11949;
wire n_1195;
wire n_11950;
wire n_11951;
wire n_11952;
wire n_11953;
wire n_11954;
wire n_11955;
wire n_11956;
wire n_11957;
wire n_11958;
wire n_11959;
wire n_1196;
wire n_11960;
wire n_11961;
wire n_11962;
wire n_11963;
wire n_11964;
wire n_11965;
wire n_11966;
wire n_11967;
wire n_11968;
wire n_11969;
wire n_1197;
wire n_11970;
wire n_11971;
wire n_11972;
wire n_11973;
wire n_11974;
wire n_11975;
wire n_11976;
wire n_11977;
wire n_11978;
wire n_11979;
wire n_1198;
wire n_11980;
wire n_11981;
wire n_11982;
wire n_11983;
wire n_11984;
wire n_11985;
wire n_11986;
wire n_11987;
wire n_11988;
wire n_11989;
wire n_1199;
wire n_11990;
wire n_11991;
wire n_11992;
wire n_11993;
wire n_11994;
wire n_11995;
wire n_11996;
wire n_11997;
wire n_11998;
wire n_11999;
wire n_12;
wire n_120;
wire n_1200;
wire n_12000;
wire n_12001;
wire n_12002;
wire n_12003;
wire n_12004;
wire n_12005;
wire n_12006;
wire n_12007;
wire n_12008;
wire n_12009;
wire n_1201;
wire n_12010;
wire n_12011;
wire n_12012;
wire n_12013;
wire n_12014;
wire n_12015;
wire n_12016;
wire n_12017;
wire n_12018;
wire n_12019;
wire n_1202;
wire n_12020;
wire n_12021;
wire n_12022;
wire n_12023;
wire n_12024;
wire n_12025;
wire n_12026;
wire n_12027;
wire n_12028;
wire n_12029;
wire n_1203;
wire n_12030;
wire n_12031;
wire n_12032;
wire n_12033;
wire n_12034;
wire n_12035;
wire n_12036;
wire n_12037;
wire n_12038;
wire n_12039;
wire n_1204;
wire n_12040;
wire n_12041;
wire n_12042;
wire n_12043;
wire n_12044;
wire n_12045;
wire n_12046;
wire n_12047;
wire n_12048;
wire n_12049;
wire n_1205;
wire n_12050;
wire n_12051;
wire n_12052;
wire n_12053;
wire n_12054;
wire n_12055;
wire n_12056;
wire n_12057;
wire n_12058;
wire n_12059;
wire n_1206;
wire n_12060;
wire n_12061;
wire n_12062;
wire n_12063;
wire n_12064;
wire n_12065;
wire n_12066;
wire n_12067;
wire n_12068;
wire n_12069;
wire n_1207;
wire n_12070;
wire n_12071;
wire n_12072;
wire n_12073;
wire n_12074;
wire n_12075;
wire n_12076;
wire n_12077;
wire n_12078;
wire n_12079;
wire n_1208;
wire n_12080;
wire n_12081;
wire n_12082;
wire n_12083;
wire n_12084;
wire n_12085;
wire n_12086;
wire n_12087;
wire n_12088;
wire n_12089;
wire n_1209;
wire n_12090;
wire n_12091;
wire n_12092;
wire n_12093;
wire n_12094;
wire n_12095;
wire n_12096;
wire n_12097;
wire n_12098;
wire n_12099;
wire n_121;
wire n_1210;
wire n_12100;
wire n_12101;
wire n_12102;
wire n_12103;
wire n_12104;
wire n_12105;
wire n_12106;
wire n_12107;
wire n_12108;
wire n_12109;
wire n_1211;
wire n_12110;
wire n_12111;
wire n_12112;
wire n_12113;
wire n_12114;
wire n_12115;
wire n_12116;
wire n_12117;
wire n_12118;
wire n_12119;
wire n_1212;
wire n_12120;
wire n_12121;
wire n_12122;
wire n_12123;
wire n_12124;
wire n_12125;
wire n_12126;
wire n_12127;
wire n_12128;
wire n_12129;
wire n_1213;
wire n_12130;
wire n_12131;
wire n_12132;
wire n_12133;
wire n_12134;
wire n_12135;
wire n_12136;
wire n_12137;
wire n_12138;
wire n_12139;
wire n_1214;
wire n_12140;
wire n_12141;
wire n_12142;
wire n_12143;
wire n_12144;
wire n_12145;
wire n_12146;
wire n_12147;
wire n_12148;
wire n_12149;
wire n_1215;
wire n_12150;
wire n_12151;
wire n_12152;
wire n_12153;
wire n_12154;
wire n_12155;
wire n_12156;
wire n_12157;
wire n_12158;
wire n_12159;
wire n_1216;
wire n_12160;
wire n_12161;
wire n_12162;
wire n_12163;
wire n_12164;
wire n_12165;
wire n_12166;
wire n_12167;
wire n_12168;
wire n_12169;
wire n_1217;
wire n_12170;
wire n_12171;
wire n_12172;
wire n_12173;
wire n_12174;
wire n_12175;
wire n_12176;
wire n_12177;
wire n_12178;
wire n_12179;
wire n_1218;
wire n_12180;
wire n_12181;
wire n_12182;
wire n_12183;
wire n_12184;
wire n_12185;
wire n_12186;
wire n_12187;
wire n_12188;
wire n_12189;
wire n_1219;
wire n_12190;
wire n_12191;
wire n_12192;
wire n_12193;
wire n_12194;
wire n_12195;
wire n_12196;
wire n_12197;
wire n_12198;
wire n_12199;
wire n_122;
wire n_1220;
wire n_12200;
wire n_12201;
wire n_12202;
wire n_12203;
wire n_12204;
wire n_12205;
wire n_12206;
wire n_12207;
wire n_12208;
wire n_12209;
wire n_1221;
wire n_12210;
wire n_12211;
wire n_12212;
wire n_12213;
wire n_12214;
wire n_12215;
wire n_12216;
wire n_12217;
wire n_12218;
wire n_12219;
wire n_1222;
wire n_12220;
wire n_12221;
wire n_12222;
wire n_12223;
wire n_12224;
wire n_12225;
wire n_12226;
wire n_12227;
wire n_12228;
wire n_12229;
wire n_1223;
wire n_12230;
wire n_12231;
wire n_12232;
wire n_12233;
wire n_12234;
wire n_12235;
wire n_12236;
wire n_12237;
wire n_12238;
wire n_12239;
wire n_1224;
wire n_12240;
wire n_12241;
wire n_12242;
wire n_12243;
wire n_12244;
wire n_12245;
wire n_12246;
wire n_12247;
wire n_12248;
wire n_12249;
wire n_1225;
wire n_12250;
wire n_12251;
wire n_12252;
wire n_12253;
wire n_12254;
wire n_12255;
wire n_12256;
wire n_12257;
wire n_12258;
wire n_12259;
wire n_1226;
wire n_12260;
wire n_12261;
wire n_12262;
wire n_12263;
wire n_12264;
wire n_12265;
wire n_12266;
wire n_12267;
wire n_12268;
wire n_12269;
wire n_1227;
wire n_12270;
wire n_12271;
wire n_12272;
wire n_12273;
wire n_12274;
wire n_12275;
wire n_12276;
wire n_12277;
wire n_12278;
wire n_12279;
wire n_1228;
wire n_12280;
wire n_12281;
wire n_12282;
wire n_12283;
wire n_12284;
wire n_12285;
wire n_12286;
wire n_12287;
wire n_12288;
wire n_12289;
wire n_1229;
wire n_12290;
wire n_12291;
wire n_12292;
wire n_12293;
wire n_12294;
wire n_12295;
wire n_12296;
wire n_12297;
wire n_12298;
wire n_12299;
wire n_123;
wire n_1230;
wire n_12300;
wire n_12301;
wire n_12302;
wire n_12303;
wire n_12304;
wire n_12305;
wire n_12306;
wire n_12307;
wire n_12308;
wire n_12309;
wire n_1231;
wire n_12310;
wire n_12311;
wire n_12312;
wire n_12313;
wire n_12314;
wire n_12315;
wire n_12316;
wire n_12317;
wire n_12318;
wire n_12319;
wire n_1232;
wire n_12320;
wire n_12321;
wire n_12322;
wire n_12323;
wire n_12324;
wire n_12325;
wire n_12326;
wire n_12327;
wire n_12328;
wire n_12329;
wire n_1233;
wire n_12330;
wire n_12331;
wire n_12332;
wire n_12333;
wire n_12334;
wire n_12335;
wire n_12336;
wire n_12337;
wire n_12338;
wire n_12339;
wire n_1234;
wire n_12340;
wire n_12341;
wire n_12342;
wire n_12343;
wire n_12344;
wire n_12345;
wire n_12346;
wire n_12347;
wire n_12348;
wire n_12349;
wire n_1235;
wire n_12350;
wire n_12351;
wire n_12352;
wire n_12353;
wire n_12354;
wire n_12355;
wire n_12356;
wire n_12357;
wire n_12358;
wire n_12359;
wire n_1236;
wire n_12360;
wire n_12361;
wire n_12362;
wire n_12363;
wire n_12364;
wire n_12365;
wire n_12366;
wire n_12367;
wire n_12368;
wire n_12369;
wire n_1237;
wire n_12370;
wire n_12371;
wire n_12372;
wire n_12373;
wire n_12374;
wire n_12375;
wire n_12376;
wire n_12377;
wire n_12378;
wire n_12379;
wire n_1238;
wire n_12380;
wire n_12381;
wire n_12382;
wire n_12383;
wire n_12384;
wire n_12385;
wire n_12386;
wire n_12387;
wire n_12388;
wire n_12389;
wire n_1239;
wire n_12390;
wire n_12391;
wire n_12392;
wire n_12393;
wire n_12394;
wire n_12395;
wire n_12396;
wire n_12397;
wire n_12398;
wire n_12399;
wire n_124;
wire n_1240;
wire n_12400;
wire n_12401;
wire n_12402;
wire n_12403;
wire n_12404;
wire n_12405;
wire n_12406;
wire n_12407;
wire n_12408;
wire n_12409;
wire n_1241;
wire n_12410;
wire n_12411;
wire n_12412;
wire n_12413;
wire n_12414;
wire n_12415;
wire n_12416;
wire n_12417;
wire n_12418;
wire n_12419;
wire n_1242;
wire n_12420;
wire n_12421;
wire n_12422;
wire n_12423;
wire n_12424;
wire n_12425;
wire n_12426;
wire n_12427;
wire n_12428;
wire n_12429;
wire n_1243;
wire n_12430;
wire n_12431;
wire n_12432;
wire n_12433;
wire n_12434;
wire n_12435;
wire n_12436;
wire n_12437;
wire n_12438;
wire n_12439;
wire n_1244;
wire n_12440;
wire n_12441;
wire n_12442;
wire n_12443;
wire n_12444;
wire n_12445;
wire n_12446;
wire n_12447;
wire n_12448;
wire n_12449;
wire n_1245;
wire n_12450;
wire n_12451;
wire n_12452;
wire n_12453;
wire n_12454;
wire n_12455;
wire n_12456;
wire n_12457;
wire n_12458;
wire n_12459;
wire n_1246;
wire n_12460;
wire n_12461;
wire n_12462;
wire n_12463;
wire n_12464;
wire n_12465;
wire n_12466;
wire n_12467;
wire n_12468;
wire n_12469;
wire n_1247;
wire n_12470;
wire n_12471;
wire n_12472;
wire n_12473;
wire n_12474;
wire n_12475;
wire n_12476;
wire n_12477;
wire n_12478;
wire n_12479;
wire n_1248;
wire n_12480;
wire n_12481;
wire n_12482;
wire n_12483;
wire n_12484;
wire n_12485;
wire n_12486;
wire n_12487;
wire n_12488;
wire n_12489;
wire n_1249;
wire n_12490;
wire n_12491;
wire n_12492;
wire n_12493;
wire n_12494;
wire n_12495;
wire n_12496;
wire n_12497;
wire n_12498;
wire n_12499;
wire n_125;
wire n_1250;
wire n_12500;
wire n_12501;
wire n_12502;
wire n_12503;
wire n_12504;
wire n_12505;
wire n_12506;
wire n_12507;
wire n_12508;
wire n_12509;
wire n_1251;
wire n_12510;
wire n_12511;
wire n_12512;
wire n_12513;
wire n_12514;
wire n_12515;
wire n_12516;
wire n_12517;
wire n_12518;
wire n_12519;
wire n_1252;
wire n_12520;
wire n_12521;
wire n_12522;
wire n_12523;
wire n_12524;
wire n_12525;
wire n_12526;
wire n_12527;
wire n_12528;
wire n_12529;
wire n_1253;
wire n_12530;
wire n_12531;
wire n_12532;
wire n_12533;
wire n_12534;
wire n_12535;
wire n_12536;
wire n_12537;
wire n_12538;
wire n_12539;
wire n_1254;
wire n_12540;
wire n_12541;
wire n_12542;
wire n_12543;
wire n_12544;
wire n_12545;
wire n_12546;
wire n_12547;
wire n_12548;
wire n_12549;
wire n_1255;
wire n_12550;
wire n_12551;
wire n_12552;
wire n_12553;
wire n_12554;
wire n_12555;
wire n_12556;
wire n_12557;
wire n_12558;
wire n_12559;
wire n_1256;
wire n_12560;
wire n_12561;
wire n_12562;
wire n_12563;
wire n_12564;
wire n_12565;
wire n_12566;
wire n_12567;
wire n_12568;
wire n_12569;
wire n_1257;
wire n_12570;
wire n_12571;
wire n_12572;
wire n_12573;
wire n_12574;
wire n_12575;
wire n_12576;
wire n_12577;
wire n_12578;
wire n_12579;
wire n_1258;
wire n_12580;
wire n_12581;
wire n_12582;
wire n_12583;
wire n_12584;
wire n_12585;
wire n_12586;
wire n_12587;
wire n_12588;
wire n_12589;
wire n_1259;
wire n_12590;
wire n_12591;
wire n_12592;
wire n_12593;
wire n_12594;
wire n_12595;
wire n_12596;
wire n_12597;
wire n_12598;
wire n_12599;
wire n_126;
wire n_1260;
wire n_12600;
wire n_12601;
wire n_12602;
wire n_12603;
wire n_12604;
wire n_12605;
wire n_12606;
wire n_12607;
wire n_12608;
wire n_12609;
wire n_1261;
wire n_12610;
wire n_12611;
wire n_12612;
wire n_12613;
wire n_12614;
wire n_12615;
wire n_12616;
wire n_12617;
wire n_12618;
wire n_12619;
wire n_1262;
wire n_12620;
wire n_12621;
wire n_12622;
wire n_12623;
wire n_12624;
wire n_12625;
wire n_12626;
wire n_12627;
wire n_12628;
wire n_12629;
wire n_1263;
wire n_12630;
wire n_12631;
wire n_12632;
wire n_12633;
wire n_12634;
wire n_12635;
wire n_12636;
wire n_12637;
wire n_12638;
wire n_12639;
wire n_1264;
wire n_12640;
wire n_12641;
wire n_12642;
wire n_12643;
wire n_12644;
wire n_12645;
wire n_12646;
wire n_12647;
wire n_12648;
wire n_12649;
wire n_1265;
wire n_12650;
wire n_12651;
wire n_12652;
wire n_12653;
wire n_12654;
wire n_12655;
wire n_12656;
wire n_12657;
wire n_12658;
wire n_12659;
wire n_1266;
wire n_12660;
wire n_12661;
wire n_12662;
wire n_12663;
wire n_12664;
wire n_12665;
wire n_12666;
wire n_12667;
wire n_12668;
wire n_12669;
wire n_1267;
wire n_12670;
wire n_12671;
wire n_12672;
wire n_12673;
wire n_12674;
wire n_12675;
wire n_12676;
wire n_12677;
wire n_12678;
wire n_12679;
wire n_1268;
wire n_12680;
wire n_12681;
wire n_12682;
wire n_12683;
wire n_12684;
wire n_12685;
wire n_12686;
wire n_12687;
wire n_12688;
wire n_12689;
wire n_1269;
wire n_12690;
wire n_12691;
wire n_12692;
wire n_12693;
wire n_12694;
wire n_12695;
wire n_12696;
wire n_12697;
wire n_12698;
wire n_12699;
wire n_127;
wire n_1270;
wire n_12700;
wire n_12701;
wire n_12702;
wire n_12703;
wire n_12704;
wire n_12705;
wire n_12706;
wire n_12707;
wire n_12708;
wire n_12709;
wire n_1271;
wire n_12710;
wire n_12711;
wire n_12712;
wire n_12713;
wire n_12714;
wire n_12715;
wire n_12716;
wire n_12717;
wire n_12718;
wire n_12719;
wire n_1272;
wire n_12720;
wire n_12721;
wire n_12722;
wire n_12723;
wire n_12724;
wire n_12725;
wire n_12726;
wire n_12727;
wire n_12728;
wire n_12729;
wire n_1273;
wire n_12730;
wire n_12731;
wire n_12732;
wire n_12733;
wire n_12734;
wire n_12735;
wire n_12736;
wire n_12737;
wire n_12738;
wire n_12739;
wire n_1274;
wire n_12740;
wire n_12741;
wire n_12742;
wire n_12743;
wire n_12744;
wire n_12745;
wire n_12746;
wire n_12747;
wire n_12748;
wire n_12749;
wire n_1275;
wire n_12750;
wire n_12751;
wire n_12752;
wire n_12753;
wire n_12754;
wire n_12755;
wire n_12756;
wire n_12757;
wire n_12758;
wire n_12759;
wire n_1276;
wire n_12760;
wire n_12761;
wire n_12762;
wire n_12763;
wire n_12764;
wire n_12765;
wire n_12766;
wire n_12767;
wire n_12768;
wire n_12769;
wire n_1277;
wire n_12770;
wire n_12771;
wire n_12772;
wire n_12773;
wire n_12774;
wire n_12775;
wire n_12776;
wire n_12777;
wire n_12778;
wire n_12779;
wire n_1278;
wire n_12780;
wire n_12781;
wire n_12782;
wire n_12783;
wire n_12784;
wire n_12785;
wire n_12786;
wire n_12787;
wire n_12788;
wire n_12789;
wire n_1279;
wire n_12790;
wire n_12791;
wire n_12792;
wire n_12793;
wire n_12794;
wire n_12795;
wire n_12796;
wire n_12797;
wire n_12798;
wire n_12799;
wire n_128;
wire n_1280;
wire n_12800;
wire n_12801;
wire n_12802;
wire n_12803;
wire n_12804;
wire n_12805;
wire n_12806;
wire n_12807;
wire n_12808;
wire n_12809;
wire n_1281;
wire n_12810;
wire n_12811;
wire n_12812;
wire n_12813;
wire n_12814;
wire n_12815;
wire n_12816;
wire n_12817;
wire n_12818;
wire n_12819;
wire n_1282;
wire n_12820;
wire n_12821;
wire n_12822;
wire n_12823;
wire n_12824;
wire n_12825;
wire n_12826;
wire n_12827;
wire n_12828;
wire n_12829;
wire n_1283;
wire n_12830;
wire n_12831;
wire n_12832;
wire n_12833;
wire n_12834;
wire n_12835;
wire n_12836;
wire n_12837;
wire n_12838;
wire n_12839;
wire n_1284;
wire n_12840;
wire n_12841;
wire n_12842;
wire n_12843;
wire n_12844;
wire n_12845;
wire n_12846;
wire n_12847;
wire n_12848;
wire n_12849;
wire n_1285;
wire n_12850;
wire n_12851;
wire n_12852;
wire n_12853;
wire n_12854;
wire n_12855;
wire n_12856;
wire n_12857;
wire n_12858;
wire n_12859;
wire n_1286;
wire n_12860;
wire n_12861;
wire n_12862;
wire n_12863;
wire n_12864;
wire n_12865;
wire n_12866;
wire n_12867;
wire n_12868;
wire n_12869;
wire n_1287;
wire n_12870;
wire n_12871;
wire n_12872;
wire n_12873;
wire n_12874;
wire n_12875;
wire n_12876;
wire n_12877;
wire n_12878;
wire n_12879;
wire n_1288;
wire n_12880;
wire n_12881;
wire n_12882;
wire n_12883;
wire n_12884;
wire n_12885;
wire n_12886;
wire n_12887;
wire n_12888;
wire n_12889;
wire n_1289;
wire n_12890;
wire n_12891;
wire n_12892;
wire n_12893;
wire n_12894;
wire n_12895;
wire n_12896;
wire n_12897;
wire n_12898;
wire n_12899;
wire n_129;
wire n_1290;
wire n_12900;
wire n_12901;
wire n_12902;
wire n_12903;
wire n_12904;
wire n_12905;
wire n_12906;
wire n_12907;
wire n_12908;
wire n_12909;
wire n_1291;
wire n_12910;
wire n_12911;
wire n_12912;
wire n_12913;
wire n_12914;
wire n_12915;
wire n_12916;
wire n_12917;
wire n_12918;
wire n_12919;
wire n_1292;
wire n_12920;
wire n_12921;
wire n_12922;
wire n_12923;
wire n_12924;
wire n_12925;
wire n_12926;
wire n_12927;
wire n_12928;
wire n_12929;
wire n_1293;
wire n_12930;
wire n_12931;
wire n_12932;
wire n_12933;
wire n_12934;
wire n_12935;
wire n_12936;
wire n_12937;
wire n_12938;
wire n_12939;
wire n_1294;
wire n_12940;
wire n_12941;
wire n_12942;
wire n_12943;
wire n_12944;
wire n_12945;
wire n_12946;
wire n_12947;
wire n_12948;
wire n_12949;
wire n_1295;
wire n_12950;
wire n_12951;
wire n_12952;
wire n_12953;
wire n_12954;
wire n_12955;
wire n_12956;
wire n_12957;
wire n_12958;
wire n_12959;
wire n_1296;
wire n_12960;
wire n_12961;
wire n_12962;
wire n_12963;
wire n_12964;
wire n_12965;
wire n_12966;
wire n_12967;
wire n_12968;
wire n_12969;
wire n_1297;
wire n_12970;
wire n_12971;
wire n_12972;
wire n_12973;
wire n_12974;
wire n_12975;
wire n_12976;
wire n_12977;
wire n_12978;
wire n_12979;
wire n_1298;
wire n_12980;
wire n_12981;
wire n_12982;
wire n_12983;
wire n_12984;
wire n_12985;
wire n_12986;
wire n_12987;
wire n_12988;
wire n_12989;
wire n_1299;
wire n_12990;
wire n_12991;
wire n_12992;
wire n_12993;
wire n_12994;
wire n_12995;
wire n_12996;
wire n_12997;
wire n_12998;
wire n_12999;
wire n_13;
wire n_130;
wire n_1300;
wire n_13000;
wire n_13001;
wire n_13002;
wire n_13003;
wire n_13004;
wire n_13005;
wire n_13006;
wire n_13007;
wire n_13008;
wire n_13009;
wire n_1301;
wire n_13010;
wire n_13011;
wire n_13012;
wire n_13013;
wire n_13014;
wire n_13015;
wire n_13016;
wire n_13017;
wire n_13018;
wire n_13019;
wire n_1302;
wire n_13020;
wire n_13021;
wire n_13022;
wire n_13023;
wire n_13024;
wire n_13025;
wire n_13026;
wire n_13027;
wire n_13028;
wire n_13029;
wire n_1303;
wire n_13030;
wire n_13031;
wire n_13032;
wire n_13033;
wire n_13034;
wire n_13035;
wire n_13036;
wire n_13037;
wire n_13038;
wire n_13039;
wire n_1304;
wire n_13040;
wire n_13041;
wire n_13042;
wire n_13043;
wire n_13044;
wire n_13045;
wire n_13046;
wire n_13047;
wire n_13048;
wire n_13049;
wire n_1305;
wire n_13050;
wire n_13051;
wire n_13052;
wire n_13053;
wire n_13054;
wire n_13055;
wire n_13056;
wire n_13057;
wire n_13058;
wire n_13059;
wire n_1306;
wire n_13060;
wire n_13061;
wire n_13062;
wire n_13063;
wire n_13064;
wire n_13065;
wire n_13066;
wire n_13067;
wire n_13068;
wire n_13069;
wire n_1307;
wire n_13070;
wire n_13071;
wire n_13072;
wire n_13073;
wire n_13074;
wire n_13075;
wire n_13076;
wire n_13077;
wire n_13078;
wire n_13079;
wire n_1308;
wire n_13080;
wire n_13081;
wire n_13082;
wire n_13083;
wire n_13084;
wire n_13085;
wire n_13086;
wire n_13087;
wire n_13088;
wire n_13089;
wire n_1309;
wire n_13090;
wire n_13091;
wire n_13092;
wire n_13093;
wire n_13094;
wire n_13095;
wire n_13096;
wire n_13097;
wire n_13098;
wire n_13099;
wire n_131;
wire n_1310;
wire n_13100;
wire n_13101;
wire n_13102;
wire n_13103;
wire n_13104;
wire n_13105;
wire n_13106;
wire n_13107;
wire n_13108;
wire n_13109;
wire n_1311;
wire n_13110;
wire n_13111;
wire n_13112;
wire n_13113;
wire n_13114;
wire n_13115;
wire n_13116;
wire n_13117;
wire n_13118;
wire n_13119;
wire n_1312;
wire n_13120;
wire n_13121;
wire n_13122;
wire n_13123;
wire n_13124;
wire n_13125;
wire n_13126;
wire n_13127;
wire n_13128;
wire n_13129;
wire n_1313;
wire n_13130;
wire n_13131;
wire n_13132;
wire n_13133;
wire n_13134;
wire n_13135;
wire n_13136;
wire n_13137;
wire n_13138;
wire n_13139;
wire n_1314;
wire n_13140;
wire n_13141;
wire n_13142;
wire n_13143;
wire n_13144;
wire n_13145;
wire n_13146;
wire n_13147;
wire n_13148;
wire n_13149;
wire n_1315;
wire n_13150;
wire n_13151;
wire n_13152;
wire n_13153;
wire n_13154;
wire n_13155;
wire n_13156;
wire n_13157;
wire n_13158;
wire n_13159;
wire n_1316;
wire n_13160;
wire n_13161;
wire n_13162;
wire n_13163;
wire n_13164;
wire n_13165;
wire n_13166;
wire n_13167;
wire n_13168;
wire n_13169;
wire n_1317;
wire n_13170;
wire n_13171;
wire n_13172;
wire n_13173;
wire n_13174;
wire n_13175;
wire n_13176;
wire n_13177;
wire n_13178;
wire n_13179;
wire n_1318;
wire n_13180;
wire n_13181;
wire n_13182;
wire n_13183;
wire n_13184;
wire n_13185;
wire n_13186;
wire n_13187;
wire n_13188;
wire n_13189;
wire n_1319;
wire n_13190;
wire n_13191;
wire n_13192;
wire n_13193;
wire n_13194;
wire n_13195;
wire n_13196;
wire n_13197;
wire n_13198;
wire n_13199;
wire n_132;
wire n_1320;
wire n_13200;
wire n_13201;
wire n_13202;
wire n_13203;
wire n_13204;
wire n_13205;
wire n_13206;
wire n_13207;
wire n_13208;
wire n_13209;
wire n_1321;
wire n_13210;
wire n_13211;
wire n_13212;
wire n_13213;
wire n_13214;
wire n_13215;
wire n_13216;
wire n_13217;
wire n_13218;
wire n_13219;
wire n_1322;
wire n_13220;
wire n_13221;
wire n_13222;
wire n_13223;
wire n_13224;
wire n_13225;
wire n_13226;
wire n_13227;
wire n_13228;
wire n_13229;
wire n_1323;
wire n_13230;
wire n_13231;
wire n_13232;
wire n_13233;
wire n_13234;
wire n_13235;
wire n_13236;
wire n_13237;
wire n_13238;
wire n_13239;
wire n_1324;
wire n_13240;
wire n_13241;
wire n_13242;
wire n_13243;
wire n_13244;
wire n_13245;
wire n_13246;
wire n_13247;
wire n_13248;
wire n_13249;
wire n_1325;
wire n_13250;
wire n_13251;
wire n_13252;
wire n_13253;
wire n_13254;
wire n_13255;
wire n_13256;
wire n_13257;
wire n_13258;
wire n_13259;
wire n_1326;
wire n_13260;
wire n_13261;
wire n_13262;
wire n_13263;
wire n_13264;
wire n_13265;
wire n_13266;
wire n_13267;
wire n_13268;
wire n_13269;
wire n_1327;
wire n_13270;
wire n_13271;
wire n_13272;
wire n_13273;
wire n_13274;
wire n_13275;
wire n_13276;
wire n_13277;
wire n_13278;
wire n_13279;
wire n_1328;
wire n_13280;
wire n_13281;
wire n_13282;
wire n_13283;
wire n_13284;
wire n_13285;
wire n_13286;
wire n_13287;
wire n_13288;
wire n_13289;
wire n_1329;
wire n_13290;
wire n_13291;
wire n_13292;
wire n_13293;
wire n_13294;
wire n_13295;
wire n_13296;
wire n_13297;
wire n_13298;
wire n_13299;
wire n_133;
wire n_1330;
wire n_13300;
wire n_13301;
wire n_13302;
wire n_13303;
wire n_13304;
wire n_13305;
wire n_13306;
wire n_13307;
wire n_13308;
wire n_13309;
wire n_1331;
wire n_13310;
wire n_13311;
wire n_13312;
wire n_13313;
wire n_13314;
wire n_13315;
wire n_13316;
wire n_13317;
wire n_13318;
wire n_13319;
wire n_1332;
wire n_13320;
wire n_13321;
wire n_13322;
wire n_13323;
wire n_13324;
wire n_13325;
wire n_13326;
wire n_13327;
wire n_13328;
wire n_13329;
wire n_1333;
wire n_13330;
wire n_13331;
wire n_13332;
wire n_13333;
wire n_13334;
wire n_13335;
wire n_13336;
wire n_13337;
wire n_13338;
wire n_13339;
wire n_1334;
wire n_13340;
wire n_13341;
wire n_13342;
wire n_13343;
wire n_13344;
wire n_13345;
wire n_13346;
wire n_13347;
wire n_13348;
wire n_13349;
wire n_1335;
wire n_13350;
wire n_13351;
wire n_13352;
wire n_13353;
wire n_13354;
wire n_13355;
wire n_13356;
wire n_13357;
wire n_13358;
wire n_13359;
wire n_1336;
wire n_13360;
wire n_13361;
wire n_13362;
wire n_13363;
wire n_13364;
wire n_13365;
wire n_13366;
wire n_13367;
wire n_13368;
wire n_13369;
wire n_1337;
wire n_13370;
wire n_13371;
wire n_13372;
wire n_13373;
wire n_13374;
wire n_13375;
wire n_13376;
wire n_13377;
wire n_13378;
wire n_13379;
wire n_1338;
wire n_13380;
wire n_13381;
wire n_13382;
wire n_13383;
wire n_13384;
wire n_13385;
wire n_13386;
wire n_13387;
wire n_13388;
wire n_13389;
wire n_1339;
wire n_13390;
wire n_13391;
wire n_13392;
wire n_13393;
wire n_13394;
wire n_13395;
wire n_13396;
wire n_13397;
wire n_13398;
wire n_13399;
wire n_134;
wire n_1340;
wire n_13400;
wire n_13401;
wire n_13402;
wire n_13403;
wire n_13404;
wire n_13405;
wire n_13406;
wire n_13407;
wire n_13408;
wire n_13409;
wire n_1341;
wire n_13410;
wire n_13411;
wire n_13412;
wire n_13413;
wire n_13414;
wire n_13415;
wire n_13416;
wire n_13417;
wire n_13418;
wire n_13419;
wire n_1342;
wire n_13420;
wire n_13421;
wire n_13422;
wire n_13423;
wire n_13424;
wire n_13425;
wire n_13426;
wire n_13427;
wire n_13428;
wire n_13429;
wire n_1343;
wire n_13430;
wire n_13431;
wire n_13432;
wire n_13433;
wire n_13434;
wire n_13435;
wire n_13436;
wire n_13437;
wire n_13438;
wire n_13439;
wire n_1344;
wire n_13440;
wire n_13441;
wire n_13442;
wire n_13443;
wire n_13444;
wire n_13445;
wire n_13446;
wire n_13447;
wire n_13448;
wire n_13449;
wire n_1345;
wire n_13450;
wire n_13451;
wire n_13452;
wire n_13453;
wire n_13454;
wire n_13455;
wire n_13456;
wire n_13457;
wire n_13458;
wire n_13459;
wire n_1346;
wire n_13460;
wire n_13461;
wire n_13462;
wire n_13463;
wire n_13464;
wire n_13465;
wire n_13466;
wire n_13467;
wire n_13468;
wire n_13469;
wire n_1347;
wire n_13470;
wire n_13471;
wire n_13472;
wire n_13473;
wire n_13474;
wire n_13475;
wire n_13476;
wire n_13477;
wire n_13478;
wire n_13479;
wire n_1348;
wire n_13480;
wire n_13481;
wire n_13482;
wire n_13483;
wire n_13484;
wire n_13485;
wire n_13486;
wire n_13487;
wire n_13488;
wire n_13489;
wire n_1349;
wire n_13490;
wire n_13491;
wire n_13492;
wire n_13493;
wire n_13494;
wire n_13495;
wire n_13496;
wire n_13497;
wire n_13498;
wire n_13499;
wire n_135;
wire n_1350;
wire n_13500;
wire n_13501;
wire n_13502;
wire n_13503;
wire n_13504;
wire n_13505;
wire n_13506;
wire n_13507;
wire n_13508;
wire n_13509;
wire n_1351;
wire n_13510;
wire n_13511;
wire n_13512;
wire n_13513;
wire n_13514;
wire n_13515;
wire n_13516;
wire n_13517;
wire n_13518;
wire n_13519;
wire n_1352;
wire n_13520;
wire n_13521;
wire n_13522;
wire n_13523;
wire n_13524;
wire n_13525;
wire n_13526;
wire n_13527;
wire n_13528;
wire n_13529;
wire n_1353;
wire n_13530;
wire n_13531;
wire n_13532;
wire n_13533;
wire n_13534;
wire n_13535;
wire n_13536;
wire n_13537;
wire n_13538;
wire n_13539;
wire n_1354;
wire n_13540;
wire n_13541;
wire n_13542;
wire n_13543;
wire n_13544;
wire n_13545;
wire n_13546;
wire n_13547;
wire n_13548;
wire n_13549;
wire n_1355;
wire n_13550;
wire n_13551;
wire n_13552;
wire n_13553;
wire n_13554;
wire n_13555;
wire n_13556;
wire n_13557;
wire n_13558;
wire n_13559;
wire n_1356;
wire n_13560;
wire n_13561;
wire n_13562;
wire n_13563;
wire n_13564;
wire n_13565;
wire n_13566;
wire n_13567;
wire n_13568;
wire n_13569;
wire n_1357;
wire n_13570;
wire n_13571;
wire n_13572;
wire n_13573;
wire n_13574;
wire n_13575;
wire n_13576;
wire n_13577;
wire n_13578;
wire n_13579;
wire n_1358;
wire n_13580;
wire n_13581;
wire n_13582;
wire n_13583;
wire n_13584;
wire n_13585;
wire n_13586;
wire n_13587;
wire n_13588;
wire n_13589;
wire n_1359;
wire n_13590;
wire n_13591;
wire n_13592;
wire n_13593;
wire n_13594;
wire n_13595;
wire n_13596;
wire n_13597;
wire n_13598;
wire n_13599;
wire n_136;
wire n_1360;
wire n_13600;
wire n_13601;
wire n_13602;
wire n_13603;
wire n_13604;
wire n_13605;
wire n_13606;
wire n_13607;
wire n_13608;
wire n_13609;
wire n_1361;
wire n_13610;
wire n_13611;
wire n_13612;
wire n_13613;
wire n_13614;
wire n_13615;
wire n_13616;
wire n_13617;
wire n_13618;
wire n_13619;
wire n_1362;
wire n_13620;
wire n_13621;
wire n_13622;
wire n_13623;
wire n_13624;
wire n_13625;
wire n_13626;
wire n_13627;
wire n_13628;
wire n_13629;
wire n_1363;
wire n_13630;
wire n_13631;
wire n_13632;
wire n_13633;
wire n_13634;
wire n_13635;
wire n_13636;
wire n_13637;
wire n_13638;
wire n_13639;
wire n_1364;
wire n_13640;
wire n_13641;
wire n_13642;
wire n_13643;
wire n_13644;
wire n_13645;
wire n_13646;
wire n_13647;
wire n_13648;
wire n_13649;
wire n_1365;
wire n_13650;
wire n_13651;
wire n_13652;
wire n_13653;
wire n_13654;
wire n_13655;
wire n_13656;
wire n_13657;
wire n_13658;
wire n_13659;
wire n_1366;
wire n_13660;
wire n_13661;
wire n_13662;
wire n_13663;
wire n_13664;
wire n_13665;
wire n_13666;
wire n_13667;
wire n_13668;
wire n_13669;
wire n_1367;
wire n_13670;
wire n_13671;
wire n_13672;
wire n_13673;
wire n_13674;
wire n_13675;
wire n_13676;
wire n_13677;
wire n_13678;
wire n_13679;
wire n_1368;
wire n_13680;
wire n_13681;
wire n_13682;
wire n_13683;
wire n_13684;
wire n_13685;
wire n_13686;
wire n_13687;
wire n_13688;
wire n_13689;
wire n_1369;
wire n_13690;
wire n_13691;
wire n_13692;
wire n_13693;
wire n_13694;
wire n_13695;
wire n_13696;
wire n_13697;
wire n_13698;
wire n_13699;
wire n_137;
wire n_1370;
wire n_13700;
wire n_13701;
wire n_13702;
wire n_13703;
wire n_13704;
wire n_13705;
wire n_13706;
wire n_13707;
wire n_13708;
wire n_13709;
wire n_1371;
wire n_13710;
wire n_13711;
wire n_13712;
wire n_13713;
wire n_13714;
wire n_13715;
wire n_13716;
wire n_13717;
wire n_13718;
wire n_13719;
wire n_1372;
wire n_13720;
wire n_13721;
wire n_13722;
wire n_13723;
wire n_13724;
wire n_13725;
wire n_13726;
wire n_13727;
wire n_13728;
wire n_13729;
wire n_1373;
wire n_13730;
wire n_13731;
wire n_13732;
wire n_13733;
wire n_13734;
wire n_13735;
wire n_13736;
wire n_13737;
wire n_13738;
wire n_13739;
wire n_1374;
wire n_13740;
wire n_13741;
wire n_13742;
wire n_13743;
wire n_13744;
wire n_13745;
wire n_13746;
wire n_13747;
wire n_13748;
wire n_13749;
wire n_1375;
wire n_13750;
wire n_13751;
wire n_13752;
wire n_13753;
wire n_13754;
wire n_13755;
wire n_13756;
wire n_13757;
wire n_13758;
wire n_13759;
wire n_1376;
wire n_13760;
wire n_13761;
wire n_13762;
wire n_13763;
wire n_13764;
wire n_13765;
wire n_13766;
wire n_13767;
wire n_13768;
wire n_13769;
wire n_1377;
wire n_13770;
wire n_13771;
wire n_13772;
wire n_13773;
wire n_13774;
wire n_13775;
wire n_13776;
wire n_13777;
wire n_13778;
wire n_13779;
wire n_1378;
wire n_13780;
wire n_13781;
wire n_13782;
wire n_13783;
wire n_13784;
wire n_13785;
wire n_13786;
wire n_13787;
wire n_13788;
wire n_13789;
wire n_1379;
wire n_13790;
wire n_13791;
wire n_13792;
wire n_13793;
wire n_13794;
wire n_13795;
wire n_13796;
wire n_13797;
wire n_13798;
wire n_13799;
wire n_138;
wire n_1380;
wire n_13800;
wire n_13801;
wire n_13802;
wire n_13803;
wire n_13804;
wire n_13805;
wire n_13806;
wire n_13807;
wire n_13808;
wire n_13809;
wire n_1381;
wire n_13810;
wire n_13811;
wire n_13812;
wire n_13813;
wire n_13814;
wire n_13815;
wire n_13816;
wire n_13817;
wire n_13818;
wire n_13819;
wire n_1382;
wire n_13820;
wire n_13821;
wire n_13822;
wire n_13823;
wire n_13824;
wire n_13825;
wire n_13826;
wire n_13827;
wire n_13828;
wire n_13829;
wire n_1383;
wire n_13830;
wire n_13831;
wire n_13832;
wire n_13833;
wire n_13834;
wire n_13835;
wire n_13836;
wire n_13837;
wire n_13838;
wire n_13839;
wire n_1384;
wire n_13840;
wire n_13841;
wire n_13842;
wire n_13843;
wire n_13844;
wire n_13845;
wire n_13846;
wire n_13847;
wire n_13848;
wire n_13849;
wire n_1385;
wire n_13850;
wire n_13851;
wire n_13852;
wire n_13853;
wire n_13854;
wire n_13855;
wire n_13856;
wire n_13857;
wire n_13858;
wire n_13859;
wire n_1386;
wire n_13860;
wire n_13861;
wire n_13862;
wire n_13863;
wire n_13864;
wire n_13865;
wire n_13866;
wire n_13867;
wire n_13868;
wire n_13869;
wire n_1387;
wire n_13870;
wire n_13871;
wire n_13872;
wire n_13873;
wire n_13874;
wire n_13875;
wire n_13876;
wire n_13877;
wire n_13878;
wire n_13879;
wire n_1388;
wire n_13880;
wire n_13881;
wire n_13882;
wire n_13883;
wire n_13884;
wire n_13885;
wire n_13886;
wire n_13887;
wire n_13888;
wire n_13889;
wire n_1389;
wire n_13890;
wire n_13891;
wire n_13892;
wire n_13893;
wire n_13894;
wire n_13895;
wire n_13896;
wire n_13897;
wire n_13898;
wire n_13899;
wire n_139;
wire n_1390;
wire n_13900;
wire n_13901;
wire n_13902;
wire n_13903;
wire n_13904;
wire n_13905;
wire n_13906;
wire n_13907;
wire n_13908;
wire n_13909;
wire n_1391;
wire n_13910;
wire n_13911;
wire n_13912;
wire n_13913;
wire n_13914;
wire n_13915;
wire n_13916;
wire n_13917;
wire n_13918;
wire n_13919;
wire n_1392;
wire n_13920;
wire n_13921;
wire n_13922;
wire n_13923;
wire n_13924;
wire n_13925;
wire n_13926;
wire n_13927;
wire n_13928;
wire n_13929;
wire n_1393;
wire n_13930;
wire n_13931;
wire n_13932;
wire n_13933;
wire n_13934;
wire n_13935;
wire n_13936;
wire n_13937;
wire n_13938;
wire n_13939;
wire n_1394;
wire n_13940;
wire n_13941;
wire n_13942;
wire n_13943;
wire n_13944;
wire n_13945;
wire n_13946;
wire n_13947;
wire n_13948;
wire n_13949;
wire n_1395;
wire n_13950;
wire n_13951;
wire n_13952;
wire n_13953;
wire n_13954;
wire n_13955;
wire n_13956;
wire n_13957;
wire n_13958;
wire n_13959;
wire n_1396;
wire n_13960;
wire n_13961;
wire n_13962;
wire n_13963;
wire n_13964;
wire n_13965;
wire n_13966;
wire n_13967;
wire n_13968;
wire n_13969;
wire n_1397;
wire n_13970;
wire n_13971;
wire n_13972;
wire n_13973;
wire n_13974;
wire n_13975;
wire n_13976;
wire n_13977;
wire n_13978;
wire n_13979;
wire n_1398;
wire n_13980;
wire n_13981;
wire n_13982;
wire n_13983;
wire n_13984;
wire n_13985;
wire n_13986;
wire n_13987;
wire n_13988;
wire n_13989;
wire n_1399;
wire n_13990;
wire n_13991;
wire n_13992;
wire n_13993;
wire n_13994;
wire n_13995;
wire n_13996;
wire n_13997;
wire n_13998;
wire n_13999;
wire n_14;
wire n_140;
wire n_1400;
wire n_14000;
wire n_14001;
wire n_14002;
wire n_14003;
wire n_14004;
wire n_14005;
wire n_14006;
wire n_14007;
wire n_14008;
wire n_14009;
wire n_1401;
wire n_14010;
wire n_14011;
wire n_14012;
wire n_14013;
wire n_14014;
wire n_14015;
wire n_14016;
wire n_14017;
wire n_14018;
wire n_14019;
wire n_1402;
wire n_14020;
wire n_14021;
wire n_14022;
wire n_14023;
wire n_14024;
wire n_14025;
wire n_14026;
wire n_14027;
wire n_14028;
wire n_14029;
wire n_1403;
wire n_14030;
wire n_14031;
wire n_14032;
wire n_14033;
wire n_14034;
wire n_14035;
wire n_14036;
wire n_14037;
wire n_14038;
wire n_14039;
wire n_1404;
wire n_14040;
wire n_14041;
wire n_14042;
wire n_14043;
wire n_14044;
wire n_14045;
wire n_14046;
wire n_14047;
wire n_14048;
wire n_14049;
wire n_1405;
wire n_14050;
wire n_14051;
wire n_14052;
wire n_14053;
wire n_14054;
wire n_14055;
wire n_14056;
wire n_14057;
wire n_14058;
wire n_14059;
wire n_1406;
wire n_14060;
wire n_14061;
wire n_14062;
wire n_14063;
wire n_14064;
wire n_14065;
wire n_14066;
wire n_14067;
wire n_14068;
wire n_14069;
wire n_1407;
wire n_14070;
wire n_14071;
wire n_14072;
wire n_14073;
wire n_14075;
wire n_14076;
wire n_14077;
wire n_14078;
wire n_14079;
wire n_1408;
wire n_14080;
wire n_14081;
wire n_14082;
wire n_14083;
wire n_14084;
wire n_14085;
wire n_14086;
wire n_14087;
wire n_14088;
wire n_14089;
wire n_1409;
wire n_14090;
wire n_14091;
wire n_14092;
wire n_14093;
wire n_14094;
wire n_14095;
wire n_14096;
wire n_14097;
wire n_14098;
wire n_14099;
wire n_141;
wire n_1410;
wire n_14100;
wire n_14101;
wire n_14102;
wire n_14103;
wire n_14104;
wire n_14105;
wire n_14106;
wire n_14107;
wire n_14108;
wire n_14109;
wire n_1411;
wire n_14110;
wire n_14111;
wire n_14112;
wire n_14113;
wire n_14114;
wire n_14115;
wire n_14116;
wire n_14117;
wire n_14118;
wire n_14119;
wire n_1412;
wire n_14120;
wire n_14121;
wire n_14122;
wire n_14123;
wire n_14124;
wire n_14125;
wire n_14126;
wire n_14127;
wire n_14128;
wire n_14129;
wire n_1413;
wire n_14130;
wire n_14131;
wire n_14132;
wire n_14133;
wire n_14134;
wire n_14135;
wire n_14136;
wire n_14137;
wire n_14138;
wire n_14139;
wire n_1414;
wire n_14140;
wire n_14141;
wire n_14142;
wire n_14143;
wire n_14144;
wire n_14145;
wire n_14146;
wire n_14147;
wire n_14148;
wire n_14149;
wire n_1415;
wire n_14150;
wire n_14151;
wire n_14152;
wire n_14153;
wire n_14154;
wire n_14155;
wire n_14156;
wire n_14157;
wire n_14158;
wire n_14159;
wire n_1416;
wire n_14160;
wire n_14161;
wire n_14162;
wire n_14163;
wire n_14164;
wire n_14165;
wire n_14166;
wire n_14167;
wire n_14168;
wire n_14169;
wire n_1417;
wire n_14170;
wire n_14171;
wire n_14172;
wire n_14173;
wire n_14174;
wire n_14175;
wire n_14176;
wire n_14177;
wire n_14178;
wire n_14179;
wire n_1418;
wire n_14180;
wire n_14181;
wire n_14182;
wire n_14183;
wire n_14184;
wire n_14185;
wire n_14186;
wire n_14187;
wire n_14188;
wire n_14189;
wire n_1419;
wire n_14190;
wire n_14191;
wire n_14192;
wire n_14193;
wire n_14194;
wire n_14195;
wire n_14196;
wire n_14197;
wire n_14198;
wire n_14199;
wire n_142;
wire n_1420;
wire n_14200;
wire n_14201;
wire n_14202;
wire n_14203;
wire n_14204;
wire n_14205;
wire n_14206;
wire n_14207;
wire n_14208;
wire n_14209;
wire n_1421;
wire n_14210;
wire n_14211;
wire n_14212;
wire n_14213;
wire n_14214;
wire n_14215;
wire n_14216;
wire n_14217;
wire n_14218;
wire n_14219;
wire n_1422;
wire n_14220;
wire n_14221;
wire n_14222;
wire n_14223;
wire n_14224;
wire n_14225;
wire n_14226;
wire n_14227;
wire n_14228;
wire n_14229;
wire n_1423;
wire n_14230;
wire n_14231;
wire n_14232;
wire n_14233;
wire n_14234;
wire n_14235;
wire n_14236;
wire n_14237;
wire n_14238;
wire n_14239;
wire n_1424;
wire n_14240;
wire n_14241;
wire n_14242;
wire n_14243;
wire n_14244;
wire n_14245;
wire n_14246;
wire n_14247;
wire n_14248;
wire n_14249;
wire n_1425;
wire n_14250;
wire n_14251;
wire n_14252;
wire n_14253;
wire n_14254;
wire n_14255;
wire n_14256;
wire n_14257;
wire n_14258;
wire n_14259;
wire n_1426;
wire n_14260;
wire n_14261;
wire n_14262;
wire n_14263;
wire n_14264;
wire n_14265;
wire n_14266;
wire n_14267;
wire n_14268;
wire n_14269;
wire n_1427;
wire n_14270;
wire n_14271;
wire n_14272;
wire n_14273;
wire n_14274;
wire n_14275;
wire n_14276;
wire n_14277;
wire n_14278;
wire n_14279;
wire n_1428;
wire n_14280;
wire n_14281;
wire n_14282;
wire n_14283;
wire n_14284;
wire n_14285;
wire n_14286;
wire n_14287;
wire n_14288;
wire n_14289;
wire n_1429;
wire n_14290;
wire n_14291;
wire n_14292;
wire n_14293;
wire n_14294;
wire n_14295;
wire n_14296;
wire n_14297;
wire n_14298;
wire n_14299;
wire n_143;
wire n_1430;
wire n_14300;
wire n_14301;
wire n_14302;
wire n_14303;
wire n_14304;
wire n_14305;
wire n_14306;
wire n_14307;
wire n_14308;
wire n_14309;
wire n_1431;
wire n_14310;
wire n_14311;
wire n_14312;
wire n_14313;
wire n_14314;
wire n_14315;
wire n_14316;
wire n_14317;
wire n_14318;
wire n_14319;
wire n_1432;
wire n_14320;
wire n_14321;
wire n_14322;
wire n_14323;
wire n_14324;
wire n_14325;
wire n_14326;
wire n_14327;
wire n_14328;
wire n_14329;
wire n_1433;
wire n_14330;
wire n_14331;
wire n_14332;
wire n_14333;
wire n_14334;
wire n_14335;
wire n_14336;
wire n_14337;
wire n_14338;
wire n_14339;
wire n_1434;
wire n_14340;
wire n_14341;
wire n_14342;
wire n_14343;
wire n_14344;
wire n_14345;
wire n_14346;
wire n_14347;
wire n_14348;
wire n_14349;
wire n_1435;
wire n_14350;
wire n_14351;
wire n_14352;
wire n_14353;
wire n_14354;
wire n_14355;
wire n_14356;
wire n_14357;
wire n_14358;
wire n_14359;
wire n_1436;
wire n_14360;
wire n_14361;
wire n_14362;
wire n_14363;
wire n_14364;
wire n_14365;
wire n_14366;
wire n_14367;
wire n_14368;
wire n_14369;
wire n_1437;
wire n_14370;
wire n_14371;
wire n_14372;
wire n_14373;
wire n_14374;
wire n_14375;
wire n_14376;
wire n_14377;
wire n_14378;
wire n_14379;
wire n_1438;
wire n_14380;
wire n_14381;
wire n_14382;
wire n_14383;
wire n_14384;
wire n_14385;
wire n_14386;
wire n_14387;
wire n_14388;
wire n_14389;
wire n_1439;
wire n_14390;
wire n_14391;
wire n_14392;
wire n_14393;
wire n_14394;
wire n_14395;
wire n_14396;
wire n_14397;
wire n_14398;
wire n_14399;
wire n_144;
wire n_1440;
wire n_14400;
wire n_14401;
wire n_14402;
wire n_14403;
wire n_14404;
wire n_14405;
wire n_14406;
wire n_14407;
wire n_14408;
wire n_14409;
wire n_1441;
wire n_14410;
wire n_14411;
wire n_14412;
wire n_14413;
wire n_14414;
wire n_14415;
wire n_14416;
wire n_14417;
wire n_14418;
wire n_14419;
wire n_1442;
wire n_14420;
wire n_14421;
wire n_14422;
wire n_14423;
wire n_14424;
wire n_14425;
wire n_14426;
wire n_14427;
wire n_14428;
wire n_14429;
wire n_1443;
wire n_14430;
wire n_14431;
wire n_14432;
wire n_14433;
wire n_14434;
wire n_14435;
wire n_14436;
wire n_14437;
wire n_14438;
wire n_14439;
wire n_1444;
wire n_14440;
wire n_14441;
wire n_14442;
wire n_14443;
wire n_14444;
wire n_14445;
wire n_14446;
wire n_14447;
wire n_14448;
wire n_14449;
wire n_1445;
wire n_14450;
wire n_14451;
wire n_14452;
wire n_14453;
wire n_14454;
wire n_14455;
wire n_14456;
wire n_14457;
wire n_14458;
wire n_14459;
wire n_1446;
wire n_14460;
wire n_14461;
wire n_14462;
wire n_14463;
wire n_14464;
wire n_14465;
wire n_14466;
wire n_14467;
wire n_14468;
wire n_14469;
wire n_1447;
wire n_14470;
wire n_14471;
wire n_14472;
wire n_14473;
wire n_14474;
wire n_14475;
wire n_14476;
wire n_14477;
wire n_14478;
wire n_14479;
wire n_1448;
wire n_14480;
wire n_14481;
wire n_14482;
wire n_14483;
wire n_14484;
wire n_14485;
wire n_14486;
wire n_14487;
wire n_14488;
wire n_14489;
wire n_1449;
wire n_14490;
wire n_14491;
wire n_14492;
wire n_14493;
wire n_14494;
wire n_14495;
wire n_14496;
wire n_14497;
wire n_14498;
wire n_14499;
wire n_145;
wire n_1450;
wire n_14500;
wire n_14501;
wire n_14502;
wire n_14503;
wire n_14504;
wire n_14505;
wire n_14506;
wire n_14507;
wire n_14508;
wire n_14509;
wire n_1451;
wire n_14510;
wire n_14511;
wire n_14512;
wire n_14513;
wire n_14514;
wire n_14515;
wire n_14516;
wire n_14517;
wire n_14518;
wire n_14519;
wire n_1452;
wire n_14520;
wire n_14521;
wire n_14522;
wire n_14523;
wire n_14524;
wire n_14525;
wire n_14526;
wire n_14527;
wire n_14528;
wire n_14529;
wire n_1453;
wire n_14530;
wire n_14531;
wire n_14532;
wire n_14533;
wire n_14534;
wire n_14535;
wire n_14536;
wire n_14537;
wire n_14538;
wire n_14539;
wire n_1454;
wire n_14540;
wire n_14541;
wire n_14542;
wire n_14543;
wire n_14544;
wire n_14545;
wire n_14546;
wire n_14547;
wire n_14548;
wire n_14549;
wire n_1455;
wire n_14550;
wire n_14551;
wire n_14552;
wire n_14553;
wire n_14554;
wire n_14555;
wire n_14556;
wire n_14557;
wire n_14558;
wire n_14559;
wire n_1456;
wire n_14560;
wire n_14561;
wire n_14562;
wire n_14563;
wire n_14564;
wire n_14565;
wire n_14566;
wire n_14567;
wire n_14568;
wire n_14569;
wire n_1457;
wire n_14570;
wire n_14571;
wire n_14572;
wire n_14573;
wire n_14574;
wire n_14575;
wire n_14576;
wire n_14577;
wire n_14578;
wire n_14579;
wire n_1458;
wire n_14580;
wire n_14581;
wire n_14582;
wire n_14583;
wire n_14584;
wire n_14585;
wire n_14587;
wire n_14588;
wire n_14589;
wire n_1459;
wire n_14590;
wire n_14591;
wire n_14592;
wire n_14593;
wire n_14594;
wire n_14595;
wire n_14596;
wire n_14597;
wire n_14598;
wire n_14599;
wire n_146;
wire n_1460;
wire n_14600;
wire n_14601;
wire n_14602;
wire n_14603;
wire n_14604;
wire n_14605;
wire n_14606;
wire n_14607;
wire n_14608;
wire n_14609;
wire n_1461;
wire n_14610;
wire n_14611;
wire n_14612;
wire n_14613;
wire n_14614;
wire n_14615;
wire n_14616;
wire n_14617;
wire n_14618;
wire n_14619;
wire n_1462;
wire n_14620;
wire n_14621;
wire n_14622;
wire n_14623;
wire n_14624;
wire n_14625;
wire n_14626;
wire n_14627;
wire n_14628;
wire n_14629;
wire n_1463;
wire n_14630;
wire n_14631;
wire n_14632;
wire n_14633;
wire n_14634;
wire n_14635;
wire n_14636;
wire n_14637;
wire n_14638;
wire n_14639;
wire n_1464;
wire n_14640;
wire n_14641;
wire n_14642;
wire n_14643;
wire n_14644;
wire n_14645;
wire n_14646;
wire n_14647;
wire n_14648;
wire n_14649;
wire n_1465;
wire n_14650;
wire n_14651;
wire n_14652;
wire n_14653;
wire n_14654;
wire n_14655;
wire n_14656;
wire n_14657;
wire n_14658;
wire n_14659;
wire n_1466;
wire n_14660;
wire n_14661;
wire n_14662;
wire n_14663;
wire n_14664;
wire n_14665;
wire n_14666;
wire n_14667;
wire n_14668;
wire n_14669;
wire n_1467;
wire n_14670;
wire n_14671;
wire n_14672;
wire n_14673;
wire n_14674;
wire n_14675;
wire n_14676;
wire n_14677;
wire n_14678;
wire n_14679;
wire n_1468;
wire n_14680;
wire n_14681;
wire n_14682;
wire n_14683;
wire n_14684;
wire n_14685;
wire n_14686;
wire n_14687;
wire n_14688;
wire n_14689;
wire n_1469;
wire n_14690;
wire n_14691;
wire n_14692;
wire n_14693;
wire n_14694;
wire n_14695;
wire n_14696;
wire n_14697;
wire n_14698;
wire n_14699;
wire n_147;
wire n_1470;
wire n_14700;
wire n_14701;
wire n_14702;
wire n_14703;
wire n_14704;
wire n_14705;
wire n_14706;
wire n_14707;
wire n_14708;
wire n_14709;
wire n_1471;
wire n_14710;
wire n_14711;
wire n_14712;
wire n_14713;
wire n_14714;
wire n_14715;
wire n_14716;
wire n_14717;
wire n_14718;
wire n_14719;
wire n_1472;
wire n_14720;
wire n_14721;
wire n_14722;
wire n_14723;
wire n_14724;
wire n_14725;
wire n_14726;
wire n_14727;
wire n_14728;
wire n_14729;
wire n_1473;
wire n_14730;
wire n_14731;
wire n_14732;
wire n_14733;
wire n_14734;
wire n_14735;
wire n_14736;
wire n_14737;
wire n_14738;
wire n_14739;
wire n_1474;
wire n_14740;
wire n_14741;
wire n_14742;
wire n_14743;
wire n_14744;
wire n_14745;
wire n_14746;
wire n_14747;
wire n_14748;
wire n_14749;
wire n_1475;
wire n_14750;
wire n_14751;
wire n_14752;
wire n_14753;
wire n_14754;
wire n_14755;
wire n_14756;
wire n_14757;
wire n_14758;
wire n_14759;
wire n_1476;
wire n_14760;
wire n_14761;
wire n_14762;
wire n_14763;
wire n_14764;
wire n_14765;
wire n_14766;
wire n_14767;
wire n_14768;
wire n_14769;
wire n_1477;
wire n_14770;
wire n_14771;
wire n_14772;
wire n_14773;
wire n_14774;
wire n_14775;
wire n_14776;
wire n_14777;
wire n_14778;
wire n_14779;
wire n_1478;
wire n_14780;
wire n_14781;
wire n_14782;
wire n_14783;
wire n_14784;
wire n_14785;
wire n_14786;
wire n_14787;
wire n_14788;
wire n_14789;
wire n_1479;
wire n_14790;
wire n_14791;
wire n_14792;
wire n_14793;
wire n_14794;
wire n_14795;
wire n_14796;
wire n_14797;
wire n_14798;
wire n_14799;
wire n_148;
wire n_1480;
wire n_14800;
wire n_14801;
wire n_14802;
wire n_14803;
wire n_14804;
wire n_14805;
wire n_14806;
wire n_14807;
wire n_14808;
wire n_14809;
wire n_1481;
wire n_14810;
wire n_14811;
wire n_14812;
wire n_14813;
wire n_14814;
wire n_14815;
wire n_14816;
wire n_14817;
wire n_14818;
wire n_14819;
wire n_1482;
wire n_14820;
wire n_14821;
wire n_14822;
wire n_14823;
wire n_14824;
wire n_14825;
wire n_14826;
wire n_14827;
wire n_14828;
wire n_14829;
wire n_1483;
wire n_14830;
wire n_14831;
wire n_14832;
wire n_14833;
wire n_14834;
wire n_14835;
wire n_14836;
wire n_14837;
wire n_14838;
wire n_14839;
wire n_1484;
wire n_14840;
wire n_14841;
wire n_14842;
wire n_14843;
wire n_14844;
wire n_14845;
wire n_14846;
wire n_14847;
wire n_14848;
wire n_14849;
wire n_1485;
wire n_14850;
wire n_14851;
wire n_14852;
wire n_14853;
wire n_14854;
wire n_14855;
wire n_14856;
wire n_14857;
wire n_14858;
wire n_14859;
wire n_1486;
wire n_14860;
wire n_14861;
wire n_14862;
wire n_14863;
wire n_14864;
wire n_14865;
wire n_14866;
wire n_14867;
wire n_14868;
wire n_14869;
wire n_1487;
wire n_14870;
wire n_14871;
wire n_14872;
wire n_14873;
wire n_14874;
wire n_14875;
wire n_14876;
wire n_14877;
wire n_14878;
wire n_14879;
wire n_1488;
wire n_14880;
wire n_14881;
wire n_14882;
wire n_14883;
wire n_14884;
wire n_14885;
wire n_14886;
wire n_14887;
wire n_14888;
wire n_14889;
wire n_1489;
wire n_14890;
wire n_14891;
wire n_14892;
wire n_14893;
wire n_14894;
wire n_14895;
wire n_14896;
wire n_14897;
wire n_14898;
wire n_14899;
wire n_149;
wire n_1490;
wire n_14900;
wire n_14901;
wire n_14902;
wire n_14903;
wire n_14904;
wire n_14905;
wire n_14906;
wire n_14907;
wire n_14908;
wire n_14909;
wire n_1491;
wire n_14910;
wire n_14911;
wire n_14912;
wire n_14913;
wire n_14914;
wire n_14915;
wire n_14916;
wire n_14917;
wire n_14918;
wire n_14919;
wire n_1492;
wire n_14920;
wire n_14921;
wire n_14922;
wire n_14923;
wire n_14924;
wire n_14925;
wire n_14926;
wire n_14927;
wire n_14928;
wire n_14929;
wire n_1493;
wire n_14930;
wire n_14931;
wire n_14932;
wire n_14933;
wire n_14934;
wire n_14935;
wire n_14936;
wire n_14937;
wire n_14938;
wire n_14939;
wire n_1494;
wire n_14940;
wire n_14941;
wire n_14942;
wire n_14943;
wire n_14944;
wire n_14945;
wire n_14946;
wire n_14947;
wire n_14948;
wire n_14949;
wire n_1495;
wire n_14950;
wire n_14951;
wire n_14952;
wire n_14953;
wire n_14954;
wire n_14955;
wire n_14956;
wire n_14957;
wire n_14958;
wire n_14959;
wire n_1496;
wire n_14960;
wire n_14961;
wire n_14962;
wire n_14963;
wire n_14964;
wire n_14965;
wire n_14966;
wire n_14967;
wire n_14968;
wire n_14969;
wire n_1497;
wire n_14970;
wire n_14971;
wire n_14972;
wire n_14973;
wire n_14974;
wire n_14975;
wire n_14976;
wire n_14977;
wire n_14978;
wire n_14979;
wire n_1498;
wire n_14980;
wire n_14981;
wire n_14982;
wire n_14983;
wire n_14984;
wire n_14985;
wire n_14986;
wire n_14987;
wire n_14988;
wire n_14989;
wire n_1499;
wire n_14990;
wire n_14991;
wire n_14992;
wire n_14993;
wire n_14994;
wire n_14995;
wire n_14996;
wire n_14997;
wire n_14998;
wire n_14999;
wire n_15;
wire n_150;
wire n_1500;
wire n_15000;
wire n_15001;
wire n_15002;
wire n_15003;
wire n_15004;
wire n_15005;
wire n_15006;
wire n_15007;
wire n_15008;
wire n_15009;
wire n_1501;
wire n_15010;
wire n_15011;
wire n_15012;
wire n_15013;
wire n_15014;
wire n_15015;
wire n_15016;
wire n_15017;
wire n_15018;
wire n_15019;
wire n_1502;
wire n_15020;
wire n_15021;
wire n_15022;
wire n_15023;
wire n_15024;
wire n_15025;
wire n_15026;
wire n_15027;
wire n_15028;
wire n_15029;
wire n_1503;
wire n_15030;
wire n_15031;
wire n_15032;
wire n_15033;
wire n_15034;
wire n_15035;
wire n_15036;
wire n_15037;
wire n_15038;
wire n_15039;
wire n_1504;
wire n_15040;
wire n_15041;
wire n_15042;
wire n_15043;
wire n_15044;
wire n_15045;
wire n_15046;
wire n_15047;
wire n_15048;
wire n_15049;
wire n_1505;
wire n_15050;
wire n_15051;
wire n_15052;
wire n_15053;
wire n_15054;
wire n_15055;
wire n_15056;
wire n_15057;
wire n_15058;
wire n_15059;
wire n_1506;
wire n_15060;
wire n_15061;
wire n_15062;
wire n_15063;
wire n_15064;
wire n_15065;
wire n_15066;
wire n_15067;
wire n_15068;
wire n_15069;
wire n_1507;
wire n_15070;
wire n_15071;
wire n_15072;
wire n_15073;
wire n_15074;
wire n_15075;
wire n_15076;
wire n_15077;
wire n_15078;
wire n_15079;
wire n_1508;
wire n_15080;
wire n_15081;
wire n_15082;
wire n_15083;
wire n_15084;
wire n_15085;
wire n_15086;
wire n_15087;
wire n_15088;
wire n_15089;
wire n_1509;
wire n_15090;
wire n_15091;
wire n_15092;
wire n_15093;
wire n_15094;
wire n_15095;
wire n_15096;
wire n_15097;
wire n_15098;
wire n_15099;
wire n_151;
wire n_1510;
wire n_15100;
wire n_15101;
wire n_15102;
wire n_15103;
wire n_15104;
wire n_15105;
wire n_15106;
wire n_15107;
wire n_15108;
wire n_15109;
wire n_1511;
wire n_15110;
wire n_15111;
wire n_15112;
wire n_15113;
wire n_15114;
wire n_15115;
wire n_15116;
wire n_15117;
wire n_15118;
wire n_15119;
wire n_1512;
wire n_15120;
wire n_15121;
wire n_15122;
wire n_15123;
wire n_15124;
wire n_15125;
wire n_15126;
wire n_15127;
wire n_15128;
wire n_15129;
wire n_1513;
wire n_15130;
wire n_15131;
wire n_15132;
wire n_15133;
wire n_15134;
wire n_15135;
wire n_15136;
wire n_15137;
wire n_15138;
wire n_15139;
wire n_1514;
wire n_15140;
wire n_15141;
wire n_15142;
wire n_15143;
wire n_15144;
wire n_15145;
wire n_15146;
wire n_15147;
wire n_15148;
wire n_15149;
wire n_1515;
wire n_15150;
wire n_15151;
wire n_15152;
wire n_15153;
wire n_15154;
wire n_15155;
wire n_15156;
wire n_15157;
wire n_15158;
wire n_15159;
wire n_1516;
wire n_15160;
wire n_15161;
wire n_15162;
wire n_15163;
wire n_15164;
wire n_15165;
wire n_15166;
wire n_15167;
wire n_15168;
wire n_15169;
wire n_1517;
wire n_15170;
wire n_15171;
wire n_15172;
wire n_15173;
wire n_15174;
wire n_15175;
wire n_15176;
wire n_15177;
wire n_15178;
wire n_15179;
wire n_1518;
wire n_15180;
wire n_15181;
wire n_15182;
wire n_15183;
wire n_15184;
wire n_15185;
wire n_15186;
wire n_15187;
wire n_15188;
wire n_15189;
wire n_1519;
wire n_15190;
wire n_15191;
wire n_15192;
wire n_15193;
wire n_15194;
wire n_15195;
wire n_15196;
wire n_15197;
wire n_15198;
wire n_15199;
wire n_152;
wire n_1520;
wire n_15200;
wire n_15201;
wire n_15202;
wire n_15203;
wire n_15204;
wire n_15205;
wire n_15206;
wire n_15207;
wire n_15208;
wire n_15209;
wire n_1521;
wire n_15210;
wire n_15211;
wire n_15212;
wire n_15213;
wire n_15214;
wire n_15215;
wire n_15216;
wire n_15217;
wire n_15218;
wire n_15219;
wire n_1522;
wire n_15220;
wire n_15221;
wire n_15222;
wire n_15223;
wire n_15224;
wire n_15225;
wire n_15226;
wire n_15227;
wire n_15228;
wire n_15229;
wire n_1523;
wire n_15230;
wire n_15231;
wire n_15232;
wire n_15233;
wire n_15234;
wire n_15235;
wire n_15236;
wire n_15237;
wire n_15238;
wire n_15239;
wire n_1524;
wire n_15240;
wire n_15241;
wire n_15242;
wire n_15243;
wire n_15244;
wire n_15245;
wire n_15246;
wire n_15247;
wire n_15248;
wire n_15249;
wire n_1525;
wire n_15250;
wire n_15251;
wire n_15252;
wire n_15253;
wire n_15254;
wire n_15255;
wire n_15256;
wire n_15257;
wire n_15258;
wire n_15259;
wire n_1526;
wire n_15261;
wire n_15262;
wire n_15263;
wire n_15264;
wire n_15265;
wire n_15266;
wire n_15267;
wire n_15268;
wire n_15269;
wire n_1527;
wire n_15270;
wire n_15271;
wire n_15272;
wire n_15273;
wire n_15274;
wire n_15275;
wire n_15276;
wire n_15277;
wire n_15278;
wire n_15279;
wire n_1528;
wire n_15280;
wire n_15281;
wire n_15282;
wire n_15283;
wire n_15284;
wire n_15285;
wire n_15286;
wire n_15287;
wire n_15288;
wire n_15289;
wire n_1529;
wire n_15290;
wire n_15291;
wire n_15292;
wire n_15293;
wire n_15294;
wire n_15295;
wire n_15296;
wire n_15297;
wire n_15298;
wire n_15299;
wire n_153;
wire n_1530;
wire n_15300;
wire n_15301;
wire n_15302;
wire n_15303;
wire n_15304;
wire n_15305;
wire n_15306;
wire n_15307;
wire n_15308;
wire n_15309;
wire n_1531;
wire n_15310;
wire n_15311;
wire n_15312;
wire n_15313;
wire n_15314;
wire n_15315;
wire n_15316;
wire n_15317;
wire n_15318;
wire n_15319;
wire n_1532;
wire n_15320;
wire n_15321;
wire n_15322;
wire n_15323;
wire n_15324;
wire n_15325;
wire n_15326;
wire n_15327;
wire n_15328;
wire n_15329;
wire n_1533;
wire n_15330;
wire n_15331;
wire n_15332;
wire n_15333;
wire n_15334;
wire n_15335;
wire n_15336;
wire n_15337;
wire n_15338;
wire n_15339;
wire n_1534;
wire n_15340;
wire n_15341;
wire n_15342;
wire n_15343;
wire n_15344;
wire n_15345;
wire n_15346;
wire n_15347;
wire n_15348;
wire n_15349;
wire n_1535;
wire n_15350;
wire n_15351;
wire n_15352;
wire n_15353;
wire n_15354;
wire n_15355;
wire n_15356;
wire n_15357;
wire n_15358;
wire n_15359;
wire n_1536;
wire n_15360;
wire n_15361;
wire n_15362;
wire n_15363;
wire n_15364;
wire n_15365;
wire n_15366;
wire n_15367;
wire n_15368;
wire n_15369;
wire n_1537;
wire n_15370;
wire n_15371;
wire n_15372;
wire n_15373;
wire n_15374;
wire n_15375;
wire n_15376;
wire n_15377;
wire n_15378;
wire n_15379;
wire n_1538;
wire n_15380;
wire n_15381;
wire n_15382;
wire n_15383;
wire n_15384;
wire n_15385;
wire n_15386;
wire n_15387;
wire n_15388;
wire n_15389;
wire n_1539;
wire n_15390;
wire n_15391;
wire n_15392;
wire n_15393;
wire n_15394;
wire n_15395;
wire n_15396;
wire n_15397;
wire n_15398;
wire n_15399;
wire n_154;
wire n_1540;
wire n_15400;
wire n_15401;
wire n_15402;
wire n_15403;
wire n_15404;
wire n_15405;
wire n_15406;
wire n_15407;
wire n_15408;
wire n_15409;
wire n_1541;
wire n_15410;
wire n_15411;
wire n_15412;
wire n_15413;
wire n_15414;
wire n_15415;
wire n_15416;
wire n_15417;
wire n_15418;
wire n_15419;
wire n_1542;
wire n_15420;
wire n_15421;
wire n_15422;
wire n_15423;
wire n_15424;
wire n_15425;
wire n_15426;
wire n_15427;
wire n_15428;
wire n_15429;
wire n_1543;
wire n_15430;
wire n_15431;
wire n_15432;
wire n_15433;
wire n_15434;
wire n_15435;
wire n_15436;
wire n_15437;
wire n_15438;
wire n_15439;
wire n_1544;
wire n_15440;
wire n_15441;
wire n_15442;
wire n_15443;
wire n_15444;
wire n_15445;
wire n_15446;
wire n_15447;
wire n_15448;
wire n_15449;
wire n_1545;
wire n_15450;
wire n_15451;
wire n_15452;
wire n_15453;
wire n_15454;
wire n_15455;
wire n_15456;
wire n_15457;
wire n_15458;
wire n_15459;
wire n_1546;
wire n_15460;
wire n_15461;
wire n_15462;
wire n_15463;
wire n_15464;
wire n_15465;
wire n_15466;
wire n_15467;
wire n_15468;
wire n_15469;
wire n_1547;
wire n_15470;
wire n_15471;
wire n_15472;
wire n_15473;
wire n_15474;
wire n_15475;
wire n_15476;
wire n_15477;
wire n_15478;
wire n_15479;
wire n_1548;
wire n_15480;
wire n_15481;
wire n_15482;
wire n_15483;
wire n_15484;
wire n_15485;
wire n_15486;
wire n_15487;
wire n_15488;
wire n_15489;
wire n_1549;
wire n_15490;
wire n_15491;
wire n_15492;
wire n_15493;
wire n_15494;
wire n_15495;
wire n_15496;
wire n_15497;
wire n_15498;
wire n_15499;
wire n_155;
wire n_1550;
wire n_15500;
wire n_15501;
wire n_15502;
wire n_15503;
wire n_15504;
wire n_15505;
wire n_15506;
wire n_15507;
wire n_15508;
wire n_15509;
wire n_1551;
wire n_15510;
wire n_15511;
wire n_15512;
wire n_15513;
wire n_15514;
wire n_15515;
wire n_15516;
wire n_15517;
wire n_15518;
wire n_15519;
wire n_1552;
wire n_15520;
wire n_15521;
wire n_15522;
wire n_15523;
wire n_15524;
wire n_15525;
wire n_15526;
wire n_15527;
wire n_15528;
wire n_15529;
wire n_1553;
wire n_15530;
wire n_15531;
wire n_15532;
wire n_15533;
wire n_15534;
wire n_15535;
wire n_15536;
wire n_15537;
wire n_15538;
wire n_15539;
wire n_1554;
wire n_15540;
wire n_15541;
wire n_15542;
wire n_15543;
wire n_15544;
wire n_15545;
wire n_15546;
wire n_15547;
wire n_15548;
wire n_15549;
wire n_1555;
wire n_15550;
wire n_15551;
wire n_15552;
wire n_15553;
wire n_15554;
wire n_15555;
wire n_15556;
wire n_15557;
wire n_15558;
wire n_15559;
wire n_1556;
wire n_15560;
wire n_15561;
wire n_15562;
wire n_15563;
wire n_15564;
wire n_15565;
wire n_15566;
wire n_15567;
wire n_15568;
wire n_15569;
wire n_1557;
wire n_15570;
wire n_15571;
wire n_15572;
wire n_15573;
wire n_15574;
wire n_15575;
wire n_15576;
wire n_15577;
wire n_15578;
wire n_15579;
wire n_1558;
wire n_15580;
wire n_15581;
wire n_15582;
wire n_15583;
wire n_15584;
wire n_15585;
wire n_15586;
wire n_15587;
wire n_15588;
wire n_15589;
wire n_1559;
wire n_15590;
wire n_15591;
wire n_15592;
wire n_15593;
wire n_15594;
wire n_15595;
wire n_15596;
wire n_15597;
wire n_15598;
wire n_15599;
wire n_156;
wire n_1560;
wire n_15600;
wire n_15601;
wire n_15602;
wire n_15603;
wire n_15604;
wire n_15605;
wire n_15606;
wire n_15607;
wire n_15608;
wire n_15609;
wire n_1561;
wire n_15610;
wire n_15611;
wire n_15612;
wire n_15613;
wire n_15614;
wire n_15615;
wire n_15616;
wire n_15617;
wire n_15618;
wire n_15619;
wire n_1562;
wire n_15620;
wire n_15621;
wire n_15622;
wire n_15623;
wire n_15624;
wire n_15625;
wire n_15626;
wire n_15627;
wire n_15628;
wire n_15629;
wire n_1563;
wire n_15630;
wire n_15631;
wire n_15632;
wire n_15633;
wire n_15634;
wire n_15635;
wire n_15636;
wire n_15637;
wire n_15638;
wire n_15639;
wire n_1564;
wire n_15640;
wire n_15641;
wire n_15642;
wire n_15643;
wire n_15644;
wire n_15645;
wire n_15646;
wire n_15647;
wire n_15648;
wire n_15649;
wire n_1565;
wire n_15650;
wire n_15651;
wire n_15652;
wire n_15653;
wire n_15654;
wire n_15655;
wire n_15656;
wire n_15657;
wire n_15658;
wire n_15659;
wire n_1566;
wire n_15660;
wire n_15661;
wire n_15662;
wire n_15663;
wire n_15664;
wire n_15665;
wire n_15666;
wire n_15667;
wire n_15668;
wire n_15669;
wire n_1567;
wire n_15670;
wire n_15671;
wire n_15672;
wire n_15673;
wire n_15674;
wire n_15675;
wire n_15676;
wire n_15677;
wire n_15678;
wire n_15679;
wire n_1568;
wire n_15680;
wire n_15681;
wire n_15682;
wire n_15683;
wire n_15684;
wire n_15685;
wire n_15686;
wire n_15687;
wire n_15688;
wire n_15689;
wire n_1569;
wire n_15690;
wire n_15691;
wire n_15692;
wire n_15693;
wire n_15694;
wire n_15695;
wire n_15696;
wire n_15697;
wire n_15698;
wire n_15699;
wire n_157;
wire n_1570;
wire n_15700;
wire n_15701;
wire n_15702;
wire n_15703;
wire n_15704;
wire n_15705;
wire n_15706;
wire n_15707;
wire n_15708;
wire n_15709;
wire n_1571;
wire n_15710;
wire n_15711;
wire n_15712;
wire n_15713;
wire n_15714;
wire n_15715;
wire n_15716;
wire n_15717;
wire n_15718;
wire n_15719;
wire n_1572;
wire n_15720;
wire n_15721;
wire n_15722;
wire n_15723;
wire n_15724;
wire n_15725;
wire n_15726;
wire n_15727;
wire n_15728;
wire n_15729;
wire n_1573;
wire n_15730;
wire n_15731;
wire n_15732;
wire n_15733;
wire n_15734;
wire n_15735;
wire n_15736;
wire n_15737;
wire n_15738;
wire n_15739;
wire n_1574;
wire n_15740;
wire n_15741;
wire n_15742;
wire n_15743;
wire n_15744;
wire n_15745;
wire n_15746;
wire n_15747;
wire n_15748;
wire n_15749;
wire n_1575;
wire n_15750;
wire n_15751;
wire n_15752;
wire n_15753;
wire n_15754;
wire n_15755;
wire n_15756;
wire n_15757;
wire n_15758;
wire n_15759;
wire n_1576;
wire n_15760;
wire n_15761;
wire n_15762;
wire n_15763;
wire n_15764;
wire n_15765;
wire n_15766;
wire n_15767;
wire n_15768;
wire n_15769;
wire n_1577;
wire n_15770;
wire n_15771;
wire n_15772;
wire n_15773;
wire n_15774;
wire n_15775;
wire n_15776;
wire n_15777;
wire n_15778;
wire n_15779;
wire n_1578;
wire n_15780;
wire n_15781;
wire n_15782;
wire n_15783;
wire n_15784;
wire n_15785;
wire n_15786;
wire n_15787;
wire n_15788;
wire n_15789;
wire n_1579;
wire n_15790;
wire n_15791;
wire n_15792;
wire n_15793;
wire n_15794;
wire n_15795;
wire n_15796;
wire n_15797;
wire n_15798;
wire n_15799;
wire n_158;
wire n_1580;
wire n_15800;
wire n_15801;
wire n_15802;
wire n_15803;
wire n_15804;
wire n_15805;
wire n_15806;
wire n_15807;
wire n_15808;
wire n_15809;
wire n_1581;
wire n_15810;
wire n_15811;
wire n_15812;
wire n_15813;
wire n_15814;
wire n_15815;
wire n_15816;
wire n_15817;
wire n_15818;
wire n_15819;
wire n_1582;
wire n_15820;
wire n_15821;
wire n_15822;
wire n_15823;
wire n_15824;
wire n_15825;
wire n_15826;
wire n_15827;
wire n_15828;
wire n_15829;
wire n_1583;
wire n_15830;
wire n_15831;
wire n_15832;
wire n_15833;
wire n_15834;
wire n_15835;
wire n_15836;
wire n_15837;
wire n_15838;
wire n_15839;
wire n_1584;
wire n_15840;
wire n_15841;
wire n_15842;
wire n_15843;
wire n_15844;
wire n_15845;
wire n_15846;
wire n_15847;
wire n_15848;
wire n_15849;
wire n_1585;
wire n_15850;
wire n_15851;
wire n_15852;
wire n_15853;
wire n_15854;
wire n_15855;
wire n_15856;
wire n_15857;
wire n_15858;
wire n_15859;
wire n_1586;
wire n_15860;
wire n_15861;
wire n_15862;
wire n_15863;
wire n_15864;
wire n_15865;
wire n_15866;
wire n_15867;
wire n_15868;
wire n_15869;
wire n_1587;
wire n_15870;
wire n_15871;
wire n_15872;
wire n_15873;
wire n_15874;
wire n_15875;
wire n_15876;
wire n_15877;
wire n_15878;
wire n_15879;
wire n_1588;
wire n_15880;
wire n_15881;
wire n_15882;
wire n_15883;
wire n_15884;
wire n_15885;
wire n_15886;
wire n_15887;
wire n_15888;
wire n_15889;
wire n_1589;
wire n_15890;
wire n_15891;
wire n_15892;
wire n_15893;
wire n_15894;
wire n_15895;
wire n_15896;
wire n_15897;
wire n_15898;
wire n_15899;
wire n_159;
wire n_1590;
wire n_15900;
wire n_15901;
wire n_15902;
wire n_15903;
wire n_15904;
wire n_15905;
wire n_15906;
wire n_15907;
wire n_15908;
wire n_15909;
wire n_1591;
wire n_15910;
wire n_15911;
wire n_15912;
wire n_15913;
wire n_15914;
wire n_15915;
wire n_15916;
wire n_15917;
wire n_15918;
wire n_15919;
wire n_1592;
wire n_15920;
wire n_15921;
wire n_15922;
wire n_15923;
wire n_15924;
wire n_15925;
wire n_15926;
wire n_15927;
wire n_15928;
wire n_15929;
wire n_1593;
wire n_15930;
wire n_15931;
wire n_15932;
wire n_15933;
wire n_15934;
wire n_15935;
wire n_15936;
wire n_15937;
wire n_15938;
wire n_15939;
wire n_1594;
wire n_15940;
wire n_15941;
wire n_15942;
wire n_15943;
wire n_15944;
wire n_15945;
wire n_15946;
wire n_15947;
wire n_15948;
wire n_15949;
wire n_1595;
wire n_15950;
wire n_15951;
wire n_15952;
wire n_15953;
wire n_15954;
wire n_15955;
wire n_15956;
wire n_15957;
wire n_15958;
wire n_15959;
wire n_1596;
wire n_15960;
wire n_15961;
wire n_15962;
wire n_15963;
wire n_15964;
wire n_15965;
wire n_15966;
wire n_15967;
wire n_15968;
wire n_15969;
wire n_1597;
wire n_15970;
wire n_15971;
wire n_15972;
wire n_15973;
wire n_15974;
wire n_15975;
wire n_15976;
wire n_15977;
wire n_15978;
wire n_15979;
wire n_1598;
wire n_15980;
wire n_15981;
wire n_15982;
wire n_15983;
wire n_15984;
wire n_15985;
wire n_15986;
wire n_15987;
wire n_15988;
wire n_15989;
wire n_1599;
wire n_15990;
wire n_15991;
wire n_15992;
wire n_15993;
wire n_15994;
wire n_15995;
wire n_15996;
wire n_15997;
wire n_15998;
wire n_15999;
wire n_16;
wire n_160;
wire n_1600;
wire n_16000;
wire n_16001;
wire n_16002;
wire n_16003;
wire n_16004;
wire n_16005;
wire n_16006;
wire n_16007;
wire n_16008;
wire n_16009;
wire n_1601;
wire n_16010;
wire n_16011;
wire n_16012;
wire n_16013;
wire n_16014;
wire n_16015;
wire n_16016;
wire n_16017;
wire n_16018;
wire n_16019;
wire n_1602;
wire n_16020;
wire n_16021;
wire n_16022;
wire n_16023;
wire n_16024;
wire n_16025;
wire n_16026;
wire n_16027;
wire n_16028;
wire n_16029;
wire n_1603;
wire n_16030;
wire n_16031;
wire n_16032;
wire n_16033;
wire n_16034;
wire n_16035;
wire n_16036;
wire n_16037;
wire n_16038;
wire n_16039;
wire n_1604;
wire n_16040;
wire n_16041;
wire n_16042;
wire n_16043;
wire n_16044;
wire n_16045;
wire n_16046;
wire n_16047;
wire n_16048;
wire n_16049;
wire n_1605;
wire n_16050;
wire n_16051;
wire n_16052;
wire n_16053;
wire n_16054;
wire n_16055;
wire n_16056;
wire n_16057;
wire n_16058;
wire n_16059;
wire n_1606;
wire n_16060;
wire n_16061;
wire n_16062;
wire n_16063;
wire n_16064;
wire n_16065;
wire n_16066;
wire n_16067;
wire n_16068;
wire n_16069;
wire n_1607;
wire n_16070;
wire n_16071;
wire n_16072;
wire n_16073;
wire n_16074;
wire n_16075;
wire n_16076;
wire n_16077;
wire n_16078;
wire n_16079;
wire n_1608;
wire n_16080;
wire n_16081;
wire n_16082;
wire n_16083;
wire n_16084;
wire n_16085;
wire n_16086;
wire n_16087;
wire n_16088;
wire n_16089;
wire n_1609;
wire n_16090;
wire n_16091;
wire n_16092;
wire n_16093;
wire n_16094;
wire n_16095;
wire n_16096;
wire n_16097;
wire n_16098;
wire n_16099;
wire n_161;
wire n_1610;
wire n_16100;
wire n_16101;
wire n_16102;
wire n_16103;
wire n_16104;
wire n_16105;
wire n_16106;
wire n_16107;
wire n_16108;
wire n_16109;
wire n_1611;
wire n_16110;
wire n_16112;
wire n_16113;
wire n_16114;
wire n_16115;
wire n_16116;
wire n_16117;
wire n_16118;
wire n_16119;
wire n_1612;
wire n_16120;
wire n_16121;
wire n_16122;
wire n_16123;
wire n_16124;
wire n_16125;
wire n_16126;
wire n_16127;
wire n_16128;
wire n_16129;
wire n_1613;
wire n_16130;
wire n_16131;
wire n_16132;
wire n_16133;
wire n_16134;
wire n_16135;
wire n_16136;
wire n_16137;
wire n_16138;
wire n_16139;
wire n_1614;
wire n_16140;
wire n_16141;
wire n_16142;
wire n_16143;
wire n_16144;
wire n_16145;
wire n_16146;
wire n_16147;
wire n_16148;
wire n_16149;
wire n_1615;
wire n_16150;
wire n_16151;
wire n_16152;
wire n_16153;
wire n_16154;
wire n_16155;
wire n_16156;
wire n_16157;
wire n_16158;
wire n_16159;
wire n_1616;
wire n_16160;
wire n_16161;
wire n_16162;
wire n_16163;
wire n_16164;
wire n_16165;
wire n_16166;
wire n_16167;
wire n_16168;
wire n_16169;
wire n_1617;
wire n_16170;
wire n_16171;
wire n_16172;
wire n_16173;
wire n_16174;
wire n_16175;
wire n_16176;
wire n_16177;
wire n_16178;
wire n_16179;
wire n_1618;
wire n_16180;
wire n_16181;
wire n_16182;
wire n_16183;
wire n_16184;
wire n_16185;
wire n_16186;
wire n_16187;
wire n_16188;
wire n_16189;
wire n_1619;
wire n_16190;
wire n_16191;
wire n_16192;
wire n_16193;
wire n_16194;
wire n_16195;
wire n_16196;
wire n_16197;
wire n_16198;
wire n_16199;
wire n_162;
wire n_1620;
wire n_16200;
wire n_16201;
wire n_16202;
wire n_16203;
wire n_16204;
wire n_16205;
wire n_16206;
wire n_16207;
wire n_16208;
wire n_16209;
wire n_1621;
wire n_16210;
wire n_16211;
wire n_16212;
wire n_16213;
wire n_16214;
wire n_16215;
wire n_16216;
wire n_16217;
wire n_16218;
wire n_16219;
wire n_1622;
wire n_16220;
wire n_16221;
wire n_16222;
wire n_16223;
wire n_16224;
wire n_16225;
wire n_16226;
wire n_16227;
wire n_16228;
wire n_16229;
wire n_1623;
wire n_16230;
wire n_16231;
wire n_16232;
wire n_16233;
wire n_16234;
wire n_16235;
wire n_16236;
wire n_16237;
wire n_16238;
wire n_16239;
wire n_1624;
wire n_16240;
wire n_16242;
wire n_16243;
wire n_16244;
wire n_16245;
wire n_16246;
wire n_16247;
wire n_16248;
wire n_16249;
wire n_1625;
wire n_16250;
wire n_16251;
wire n_16252;
wire n_16253;
wire n_16254;
wire n_16255;
wire n_16256;
wire n_16257;
wire n_16258;
wire n_16259;
wire n_1626;
wire n_16260;
wire n_16261;
wire n_16262;
wire n_16263;
wire n_16264;
wire n_16265;
wire n_16266;
wire n_16267;
wire n_16268;
wire n_16269;
wire n_1627;
wire n_16270;
wire n_16271;
wire n_16272;
wire n_16273;
wire n_16274;
wire n_16275;
wire n_16276;
wire n_16277;
wire n_16278;
wire n_16279;
wire n_1628;
wire n_16280;
wire n_16281;
wire n_16282;
wire n_16283;
wire n_16284;
wire n_16285;
wire n_16286;
wire n_16287;
wire n_16288;
wire n_16289;
wire n_1629;
wire n_16290;
wire n_16291;
wire n_16292;
wire n_16293;
wire n_16294;
wire n_16295;
wire n_16296;
wire n_16297;
wire n_16298;
wire n_16299;
wire n_163;
wire n_1630;
wire n_16300;
wire n_16301;
wire n_16302;
wire n_16303;
wire n_16304;
wire n_16305;
wire n_16306;
wire n_16307;
wire n_16308;
wire n_16309;
wire n_1631;
wire n_16310;
wire n_16311;
wire n_16312;
wire n_16313;
wire n_16314;
wire n_16315;
wire n_16316;
wire n_16317;
wire n_16318;
wire n_16319;
wire n_1632;
wire n_16320;
wire n_16321;
wire n_16322;
wire n_16323;
wire n_16324;
wire n_16325;
wire n_16326;
wire n_16327;
wire n_16328;
wire n_16329;
wire n_1633;
wire n_16330;
wire n_16331;
wire n_16332;
wire n_16333;
wire n_16334;
wire n_16335;
wire n_16336;
wire n_16337;
wire n_16338;
wire n_16339;
wire n_1634;
wire n_16340;
wire n_16341;
wire n_16342;
wire n_16343;
wire n_16344;
wire n_16345;
wire n_16346;
wire n_16347;
wire n_16348;
wire n_16349;
wire n_1635;
wire n_16350;
wire n_16351;
wire n_16352;
wire n_16353;
wire n_16354;
wire n_16355;
wire n_16356;
wire n_16357;
wire n_16358;
wire n_16359;
wire n_1636;
wire n_16360;
wire n_16361;
wire n_16362;
wire n_16363;
wire n_16364;
wire n_16365;
wire n_16366;
wire n_16367;
wire n_16368;
wire n_16369;
wire n_1637;
wire n_16370;
wire n_16371;
wire n_16372;
wire n_16373;
wire n_16374;
wire n_16375;
wire n_16376;
wire n_16377;
wire n_16378;
wire n_16379;
wire n_1638;
wire n_16380;
wire n_16381;
wire n_16382;
wire n_16383;
wire n_16384;
wire n_16385;
wire n_16386;
wire n_16387;
wire n_16388;
wire n_16389;
wire n_1639;
wire n_16390;
wire n_16391;
wire n_16392;
wire n_16393;
wire n_16394;
wire n_16395;
wire n_16396;
wire n_16397;
wire n_16398;
wire n_16399;
wire n_164;
wire n_1640;
wire n_16400;
wire n_16401;
wire n_16402;
wire n_16403;
wire n_16404;
wire n_16405;
wire n_16406;
wire n_16407;
wire n_16408;
wire n_16409;
wire n_1641;
wire n_16410;
wire n_16411;
wire n_16412;
wire n_16413;
wire n_16414;
wire n_16415;
wire n_16416;
wire n_16417;
wire n_16418;
wire n_16419;
wire n_1642;
wire n_16420;
wire n_16421;
wire n_16422;
wire n_16423;
wire n_16424;
wire n_16425;
wire n_16426;
wire n_16427;
wire n_16428;
wire n_16429;
wire n_1643;
wire n_16430;
wire n_16431;
wire n_16432;
wire n_16433;
wire n_16434;
wire n_16435;
wire n_16436;
wire n_16437;
wire n_16438;
wire n_16439;
wire n_1644;
wire n_16440;
wire n_16441;
wire n_16442;
wire n_16443;
wire n_16444;
wire n_16445;
wire n_16446;
wire n_16447;
wire n_16448;
wire n_16449;
wire n_1645;
wire n_16450;
wire n_16451;
wire n_16452;
wire n_16453;
wire n_16454;
wire n_16455;
wire n_16456;
wire n_16457;
wire n_16458;
wire n_16459;
wire n_1646;
wire n_16460;
wire n_16461;
wire n_16462;
wire n_16463;
wire n_16464;
wire n_16465;
wire n_16466;
wire n_16467;
wire n_16468;
wire n_16469;
wire n_1647;
wire n_16470;
wire n_16471;
wire n_16472;
wire n_16473;
wire n_16474;
wire n_16475;
wire n_16476;
wire n_16477;
wire n_16478;
wire n_16479;
wire n_1648;
wire n_16480;
wire n_16481;
wire n_16482;
wire n_16483;
wire n_16484;
wire n_16485;
wire n_16486;
wire n_16487;
wire n_16488;
wire n_16489;
wire n_1649;
wire n_16490;
wire n_16491;
wire n_16492;
wire n_16493;
wire n_16494;
wire n_16495;
wire n_16496;
wire n_16497;
wire n_16498;
wire n_165;
wire n_1650;
wire n_16500;
wire n_16501;
wire n_16502;
wire n_16503;
wire n_16504;
wire n_16505;
wire n_16506;
wire n_16507;
wire n_16508;
wire n_16509;
wire n_1651;
wire n_16510;
wire n_16511;
wire n_16512;
wire n_16513;
wire n_16514;
wire n_16515;
wire n_16516;
wire n_16517;
wire n_16518;
wire n_16519;
wire n_1652;
wire n_16520;
wire n_16521;
wire n_16522;
wire n_16523;
wire n_16524;
wire n_16525;
wire n_16526;
wire n_16527;
wire n_16528;
wire n_16529;
wire n_1653;
wire n_16530;
wire n_16531;
wire n_16532;
wire n_16533;
wire n_16534;
wire n_16535;
wire n_16536;
wire n_16537;
wire n_16538;
wire n_16539;
wire n_1654;
wire n_16540;
wire n_16541;
wire n_16542;
wire n_16543;
wire n_16544;
wire n_16545;
wire n_16546;
wire n_16547;
wire n_16548;
wire n_16549;
wire n_1655;
wire n_16550;
wire n_16551;
wire n_16552;
wire n_16553;
wire n_16554;
wire n_16555;
wire n_16556;
wire n_16557;
wire n_16558;
wire n_16559;
wire n_1656;
wire n_16560;
wire n_16561;
wire n_16562;
wire n_16563;
wire n_16564;
wire n_16565;
wire n_16566;
wire n_16567;
wire n_16568;
wire n_16569;
wire n_1657;
wire n_16570;
wire n_16571;
wire n_16572;
wire n_16573;
wire n_16574;
wire n_16575;
wire n_16576;
wire n_16577;
wire n_16578;
wire n_16579;
wire n_1658;
wire n_16580;
wire n_16581;
wire n_16582;
wire n_16583;
wire n_16584;
wire n_16585;
wire n_16586;
wire n_16587;
wire n_16588;
wire n_16589;
wire n_1659;
wire n_16590;
wire n_16591;
wire n_16592;
wire n_16593;
wire n_16594;
wire n_16595;
wire n_16596;
wire n_16597;
wire n_16598;
wire n_16599;
wire n_166;
wire n_1660;
wire n_16600;
wire n_16601;
wire n_16602;
wire n_16603;
wire n_16604;
wire n_16605;
wire n_16606;
wire n_16607;
wire n_16608;
wire n_16609;
wire n_1661;
wire n_16610;
wire n_16611;
wire n_16612;
wire n_16613;
wire n_16614;
wire n_16615;
wire n_16616;
wire n_16617;
wire n_16618;
wire n_16619;
wire n_1662;
wire n_16620;
wire n_16621;
wire n_16622;
wire n_16623;
wire n_16624;
wire n_16625;
wire n_16626;
wire n_16627;
wire n_16628;
wire n_16629;
wire n_1663;
wire n_16630;
wire n_16631;
wire n_16632;
wire n_16633;
wire n_16634;
wire n_16635;
wire n_16636;
wire n_16637;
wire n_16638;
wire n_16639;
wire n_1664;
wire n_16640;
wire n_16641;
wire n_16642;
wire n_16643;
wire n_16644;
wire n_16645;
wire n_16646;
wire n_16647;
wire n_16648;
wire n_16649;
wire n_1665;
wire n_16650;
wire n_16651;
wire n_16652;
wire n_16653;
wire n_16654;
wire n_16655;
wire n_16656;
wire n_16657;
wire n_16658;
wire n_16659;
wire n_1666;
wire n_16660;
wire n_16661;
wire n_16662;
wire n_16663;
wire n_16664;
wire n_16665;
wire n_16666;
wire n_16667;
wire n_16668;
wire n_16669;
wire n_1667;
wire n_16670;
wire n_16671;
wire n_16672;
wire n_16673;
wire n_16674;
wire n_16675;
wire n_16676;
wire n_16677;
wire n_16678;
wire n_16679;
wire n_1668;
wire n_16680;
wire n_16681;
wire n_16682;
wire n_16683;
wire n_16684;
wire n_16685;
wire n_16686;
wire n_16687;
wire n_16688;
wire n_16689;
wire n_1669;
wire n_16690;
wire n_16691;
wire n_16692;
wire n_16693;
wire n_16694;
wire n_16695;
wire n_16696;
wire n_16697;
wire n_16698;
wire n_16699;
wire n_167;
wire n_1670;
wire n_16700;
wire n_16701;
wire n_16702;
wire n_16703;
wire n_16704;
wire n_16705;
wire n_16706;
wire n_16707;
wire n_16708;
wire n_16709;
wire n_1671;
wire n_16710;
wire n_16711;
wire n_16712;
wire n_16713;
wire n_16714;
wire n_16715;
wire n_16716;
wire n_16717;
wire n_16718;
wire n_16719;
wire n_1672;
wire n_16720;
wire n_16721;
wire n_16722;
wire n_16723;
wire n_16724;
wire n_16725;
wire n_16726;
wire n_16727;
wire n_16728;
wire n_16729;
wire n_1673;
wire n_16730;
wire n_16731;
wire n_16732;
wire n_16733;
wire n_16734;
wire n_16735;
wire n_16736;
wire n_16737;
wire n_16738;
wire n_16739;
wire n_1674;
wire n_16740;
wire n_16741;
wire n_16742;
wire n_16743;
wire n_16744;
wire n_16745;
wire n_16746;
wire n_16747;
wire n_16748;
wire n_16749;
wire n_1675;
wire n_16750;
wire n_16751;
wire n_16752;
wire n_16753;
wire n_16754;
wire n_16755;
wire n_16756;
wire n_16757;
wire n_16758;
wire n_16759;
wire n_1676;
wire n_16760;
wire n_16761;
wire n_16762;
wire n_16763;
wire n_16764;
wire n_16765;
wire n_16766;
wire n_16767;
wire n_16768;
wire n_16769;
wire n_1677;
wire n_16770;
wire n_16771;
wire n_16772;
wire n_16773;
wire n_16774;
wire n_16775;
wire n_16776;
wire n_16777;
wire n_16778;
wire n_16779;
wire n_1678;
wire n_16780;
wire n_16781;
wire n_16782;
wire n_16783;
wire n_16784;
wire n_16785;
wire n_16786;
wire n_16787;
wire n_16788;
wire n_16789;
wire n_1679;
wire n_16790;
wire n_16791;
wire n_16792;
wire n_16793;
wire n_16794;
wire n_16795;
wire n_16796;
wire n_16797;
wire n_16798;
wire n_16799;
wire n_168;
wire n_1680;
wire n_16800;
wire n_16801;
wire n_16802;
wire n_16803;
wire n_16804;
wire n_16805;
wire n_16806;
wire n_16807;
wire n_16808;
wire n_16809;
wire n_1681;
wire n_16810;
wire n_16811;
wire n_16812;
wire n_16813;
wire n_16814;
wire n_16815;
wire n_16816;
wire n_16817;
wire n_16818;
wire n_16819;
wire n_1682;
wire n_16820;
wire n_16821;
wire n_16822;
wire n_16823;
wire n_16824;
wire n_16825;
wire n_16826;
wire n_16827;
wire n_16828;
wire n_16829;
wire n_1683;
wire n_16830;
wire n_16831;
wire n_16832;
wire n_16833;
wire n_16834;
wire n_16835;
wire n_16836;
wire n_16837;
wire n_16838;
wire n_16839;
wire n_1684;
wire n_16840;
wire n_16841;
wire n_16842;
wire n_16843;
wire n_16844;
wire n_16845;
wire n_16846;
wire n_16847;
wire n_16848;
wire n_16849;
wire n_1685;
wire n_16850;
wire n_16851;
wire n_16852;
wire n_16853;
wire n_16854;
wire n_16855;
wire n_16856;
wire n_16857;
wire n_16858;
wire n_16859;
wire n_1686;
wire n_16860;
wire n_16861;
wire n_16862;
wire n_16863;
wire n_16864;
wire n_16865;
wire n_16866;
wire n_16867;
wire n_16868;
wire n_16869;
wire n_1687;
wire n_16870;
wire n_16871;
wire n_16872;
wire n_16873;
wire n_16874;
wire n_16875;
wire n_16876;
wire n_16877;
wire n_16878;
wire n_16879;
wire n_1688;
wire n_16880;
wire n_16881;
wire n_16882;
wire n_16883;
wire n_16884;
wire n_16885;
wire n_16886;
wire n_16887;
wire n_16888;
wire n_16889;
wire n_1689;
wire n_16890;
wire n_16891;
wire n_16892;
wire n_16893;
wire n_16894;
wire n_16895;
wire n_16896;
wire n_16897;
wire n_16898;
wire n_16899;
wire n_169;
wire n_1690;
wire n_16900;
wire n_16901;
wire n_16902;
wire n_16903;
wire n_16904;
wire n_16905;
wire n_16906;
wire n_16907;
wire n_16908;
wire n_16909;
wire n_1691;
wire n_16910;
wire n_16911;
wire n_16912;
wire n_16913;
wire n_16914;
wire n_16915;
wire n_16916;
wire n_16917;
wire n_16918;
wire n_16919;
wire n_1692;
wire n_16920;
wire n_16921;
wire n_16922;
wire n_16923;
wire n_16924;
wire n_16925;
wire n_16926;
wire n_16927;
wire n_16928;
wire n_16929;
wire n_1693;
wire n_16930;
wire n_16931;
wire n_16932;
wire n_16933;
wire n_16934;
wire n_16935;
wire n_16936;
wire n_16937;
wire n_16938;
wire n_16939;
wire n_1694;
wire n_16940;
wire n_16941;
wire n_16942;
wire n_16943;
wire n_16944;
wire n_16945;
wire n_16946;
wire n_16947;
wire n_16948;
wire n_16949;
wire n_1695;
wire n_16950;
wire n_16951;
wire n_16952;
wire n_16953;
wire n_16954;
wire n_16955;
wire n_16956;
wire n_16957;
wire n_16958;
wire n_16959;
wire n_1696;
wire n_16960;
wire n_16961;
wire n_16962;
wire n_16963;
wire n_16964;
wire n_16965;
wire n_16966;
wire n_16967;
wire n_16968;
wire n_16969;
wire n_1697;
wire n_16970;
wire n_16971;
wire n_16972;
wire n_16973;
wire n_16974;
wire n_16975;
wire n_16976;
wire n_16977;
wire n_16978;
wire n_16979;
wire n_1698;
wire n_16980;
wire n_16981;
wire n_16982;
wire n_16983;
wire n_16984;
wire n_16985;
wire n_16986;
wire n_16987;
wire n_16988;
wire n_16989;
wire n_1699;
wire n_16990;
wire n_16991;
wire n_16992;
wire n_16993;
wire n_16994;
wire n_16995;
wire n_16996;
wire n_16997;
wire n_16998;
wire n_16999;
wire n_17;
wire n_170;
wire n_1700;
wire n_17000;
wire n_17001;
wire n_17002;
wire n_17003;
wire n_17004;
wire n_17005;
wire n_17006;
wire n_17007;
wire n_17008;
wire n_17009;
wire n_1701;
wire n_17010;
wire n_17011;
wire n_17012;
wire n_17013;
wire n_17014;
wire n_17015;
wire n_17016;
wire n_17017;
wire n_17018;
wire n_17019;
wire n_1702;
wire n_17020;
wire n_17021;
wire n_17022;
wire n_17023;
wire n_17024;
wire n_17025;
wire n_17026;
wire n_17027;
wire n_17028;
wire n_17029;
wire n_1703;
wire n_17030;
wire n_17031;
wire n_17032;
wire n_17033;
wire n_17034;
wire n_17035;
wire n_17036;
wire n_17037;
wire n_17038;
wire n_17039;
wire n_1704;
wire n_17040;
wire n_17041;
wire n_17042;
wire n_17043;
wire n_17044;
wire n_17045;
wire n_17046;
wire n_17047;
wire n_17048;
wire n_17049;
wire n_1705;
wire n_17050;
wire n_17051;
wire n_17052;
wire n_17053;
wire n_17054;
wire n_17055;
wire n_17056;
wire n_17057;
wire n_17058;
wire n_17059;
wire n_1706;
wire n_17060;
wire n_17061;
wire n_17062;
wire n_17063;
wire n_17064;
wire n_17065;
wire n_17066;
wire n_17067;
wire n_17068;
wire n_17069;
wire n_1707;
wire n_17070;
wire n_17071;
wire n_17072;
wire n_17073;
wire n_17074;
wire n_17075;
wire n_17076;
wire n_17077;
wire n_17078;
wire n_17079;
wire n_1708;
wire n_17080;
wire n_17081;
wire n_17082;
wire n_17083;
wire n_17084;
wire n_17085;
wire n_17086;
wire n_17087;
wire n_17088;
wire n_17089;
wire n_1709;
wire n_17090;
wire n_17091;
wire n_17092;
wire n_17093;
wire n_17094;
wire n_17095;
wire n_17096;
wire n_17097;
wire n_17098;
wire n_17099;
wire n_171;
wire n_1710;
wire n_17100;
wire n_17101;
wire n_17102;
wire n_17103;
wire n_17104;
wire n_17105;
wire n_17106;
wire n_17107;
wire n_17108;
wire n_17109;
wire n_1711;
wire n_17110;
wire n_17111;
wire n_17112;
wire n_17113;
wire n_17114;
wire n_17115;
wire n_17116;
wire n_17117;
wire n_17118;
wire n_17119;
wire n_1712;
wire n_17120;
wire n_17121;
wire n_17122;
wire n_17123;
wire n_17124;
wire n_17125;
wire n_17126;
wire n_17127;
wire n_17128;
wire n_17129;
wire n_1713;
wire n_17130;
wire n_17131;
wire n_17132;
wire n_17133;
wire n_17134;
wire n_17135;
wire n_17136;
wire n_17137;
wire n_17138;
wire n_17139;
wire n_1714;
wire n_17140;
wire n_17141;
wire n_17142;
wire n_17143;
wire n_17144;
wire n_17145;
wire n_17146;
wire n_17147;
wire n_17148;
wire n_17149;
wire n_1715;
wire n_17150;
wire n_17151;
wire n_17152;
wire n_17153;
wire n_17154;
wire n_17155;
wire n_17156;
wire n_17157;
wire n_17158;
wire n_17159;
wire n_1716;
wire n_17160;
wire n_17161;
wire n_17162;
wire n_17163;
wire n_17164;
wire n_17165;
wire n_17166;
wire n_17167;
wire n_17168;
wire n_17169;
wire n_1717;
wire n_17170;
wire n_17171;
wire n_17172;
wire n_17173;
wire n_17174;
wire n_17175;
wire n_17176;
wire n_17177;
wire n_17178;
wire n_17179;
wire n_1718;
wire n_17180;
wire n_17181;
wire n_17182;
wire n_17183;
wire n_17184;
wire n_17185;
wire n_17187;
wire n_17188;
wire n_17189;
wire n_1719;
wire n_17190;
wire n_17191;
wire n_17192;
wire n_17193;
wire n_17194;
wire n_17195;
wire n_17196;
wire n_17197;
wire n_17198;
wire n_17199;
wire n_172;
wire n_1720;
wire n_17200;
wire n_17201;
wire n_17202;
wire n_17203;
wire n_17204;
wire n_17205;
wire n_17206;
wire n_17207;
wire n_17208;
wire n_17209;
wire n_1721;
wire n_17210;
wire n_17211;
wire n_17212;
wire n_17213;
wire n_17214;
wire n_17215;
wire n_17216;
wire n_17217;
wire n_17218;
wire n_17219;
wire n_1722;
wire n_17220;
wire n_17221;
wire n_17222;
wire n_17223;
wire n_17224;
wire n_17225;
wire n_17226;
wire n_17227;
wire n_17228;
wire n_17229;
wire n_1723;
wire n_17230;
wire n_17231;
wire n_17232;
wire n_17233;
wire n_17234;
wire n_17236;
wire n_17237;
wire n_17238;
wire n_17239;
wire n_1724;
wire n_17240;
wire n_17241;
wire n_17242;
wire n_17243;
wire n_17244;
wire n_17245;
wire n_17246;
wire n_17247;
wire n_17248;
wire n_17249;
wire n_1725;
wire n_17250;
wire n_17251;
wire n_17252;
wire n_17253;
wire n_17254;
wire n_17255;
wire n_17256;
wire n_17257;
wire n_17258;
wire n_17259;
wire n_1726;
wire n_17260;
wire n_17261;
wire n_17262;
wire n_17263;
wire n_17264;
wire n_17265;
wire n_17266;
wire n_17267;
wire n_17268;
wire n_17269;
wire n_1727;
wire n_17270;
wire n_17271;
wire n_17272;
wire n_17273;
wire n_17274;
wire n_17275;
wire n_17276;
wire n_17277;
wire n_17278;
wire n_17279;
wire n_1728;
wire n_17280;
wire n_17281;
wire n_17282;
wire n_17283;
wire n_17284;
wire n_17285;
wire n_17286;
wire n_17287;
wire n_17288;
wire n_17289;
wire n_1729;
wire n_17290;
wire n_17291;
wire n_17292;
wire n_17293;
wire n_17294;
wire n_17295;
wire n_17296;
wire n_17297;
wire n_17298;
wire n_17299;
wire n_173;
wire n_1730;
wire n_17300;
wire n_17301;
wire n_17302;
wire n_17303;
wire n_17304;
wire n_17305;
wire n_17306;
wire n_17307;
wire n_17308;
wire n_17309;
wire n_1731;
wire n_17310;
wire n_17311;
wire n_17312;
wire n_17313;
wire n_17314;
wire n_17315;
wire n_17316;
wire n_17317;
wire n_17318;
wire n_17319;
wire n_1732;
wire n_17320;
wire n_17321;
wire n_17322;
wire n_17323;
wire n_17324;
wire n_17325;
wire n_17326;
wire n_17327;
wire n_17328;
wire n_17329;
wire n_1733;
wire n_17330;
wire n_17331;
wire n_17332;
wire n_17333;
wire n_17334;
wire n_17335;
wire n_17336;
wire n_17337;
wire n_17338;
wire n_17339;
wire n_1734;
wire n_17340;
wire n_17341;
wire n_17342;
wire n_17343;
wire n_17344;
wire n_17345;
wire n_17346;
wire n_17347;
wire n_17348;
wire n_17349;
wire n_1735;
wire n_17350;
wire n_17351;
wire n_17352;
wire n_17353;
wire n_17354;
wire n_17355;
wire n_17356;
wire n_17357;
wire n_17358;
wire n_17359;
wire n_1736;
wire n_17360;
wire n_17361;
wire n_17362;
wire n_17363;
wire n_17364;
wire n_17365;
wire n_17366;
wire n_17367;
wire n_17368;
wire n_17369;
wire n_1737;
wire n_17370;
wire n_17371;
wire n_17372;
wire n_17373;
wire n_17374;
wire n_17375;
wire n_17376;
wire n_17377;
wire n_17378;
wire n_17379;
wire n_1738;
wire n_17380;
wire n_17381;
wire n_17382;
wire n_17383;
wire n_17384;
wire n_17385;
wire n_17386;
wire n_17387;
wire n_17388;
wire n_17389;
wire n_1739;
wire n_17390;
wire n_17391;
wire n_17392;
wire n_17393;
wire n_17394;
wire n_17395;
wire n_17396;
wire n_17397;
wire n_17398;
wire n_17399;
wire n_174;
wire n_1740;
wire n_17400;
wire n_17401;
wire n_17402;
wire n_17403;
wire n_17404;
wire n_17405;
wire n_17406;
wire n_17407;
wire n_17408;
wire n_17409;
wire n_1741;
wire n_17410;
wire n_17411;
wire n_17412;
wire n_17413;
wire n_17414;
wire n_17415;
wire n_17416;
wire n_17417;
wire n_17418;
wire n_17419;
wire n_1742;
wire n_17420;
wire n_17421;
wire n_17422;
wire n_17423;
wire n_17424;
wire n_17425;
wire n_17426;
wire n_17427;
wire n_17428;
wire n_17429;
wire n_1743;
wire n_17430;
wire n_17431;
wire n_17432;
wire n_17433;
wire n_17434;
wire n_17435;
wire n_17436;
wire n_17437;
wire n_17438;
wire n_17439;
wire n_1744;
wire n_17440;
wire n_17441;
wire n_17442;
wire n_17443;
wire n_17444;
wire n_17445;
wire n_17446;
wire n_17447;
wire n_17448;
wire n_17449;
wire n_1745;
wire n_17450;
wire n_17451;
wire n_17452;
wire n_17453;
wire n_17454;
wire n_17455;
wire n_17456;
wire n_17457;
wire n_17458;
wire n_17459;
wire n_1746;
wire n_17460;
wire n_17461;
wire n_17462;
wire n_17463;
wire n_17464;
wire n_17465;
wire n_17466;
wire n_17467;
wire n_17468;
wire n_17469;
wire n_1747;
wire n_17470;
wire n_17471;
wire n_17472;
wire n_17473;
wire n_17474;
wire n_17475;
wire n_17476;
wire n_17477;
wire n_17478;
wire n_17479;
wire n_1748;
wire n_17480;
wire n_17481;
wire n_17482;
wire n_17483;
wire n_17484;
wire n_17485;
wire n_17486;
wire n_17487;
wire n_17488;
wire n_17489;
wire n_1749;
wire n_17490;
wire n_17491;
wire n_17492;
wire n_17493;
wire n_17494;
wire n_17495;
wire n_17496;
wire n_17497;
wire n_17498;
wire n_17499;
wire n_175;
wire n_1750;
wire n_17500;
wire n_17501;
wire n_17502;
wire n_17503;
wire n_17504;
wire n_17505;
wire n_17506;
wire n_17507;
wire n_17508;
wire n_17509;
wire n_1751;
wire n_17510;
wire n_17511;
wire n_17512;
wire n_17513;
wire n_17514;
wire n_17515;
wire n_17516;
wire n_17517;
wire n_17518;
wire n_17519;
wire n_1752;
wire n_17520;
wire n_17521;
wire n_17522;
wire n_17523;
wire n_17524;
wire n_17525;
wire n_17526;
wire n_17527;
wire n_17528;
wire n_17529;
wire n_1753;
wire n_17530;
wire n_17531;
wire n_17532;
wire n_17533;
wire n_17534;
wire n_17535;
wire n_17536;
wire n_17537;
wire n_17538;
wire n_17539;
wire n_1754;
wire n_17540;
wire n_17541;
wire n_17542;
wire n_17543;
wire n_17544;
wire n_17545;
wire n_17546;
wire n_17547;
wire n_17548;
wire n_17549;
wire n_1755;
wire n_17550;
wire n_17551;
wire n_17552;
wire n_17553;
wire n_17554;
wire n_17555;
wire n_17556;
wire n_17557;
wire n_17558;
wire n_17559;
wire n_1756;
wire n_17560;
wire n_17561;
wire n_17562;
wire n_17563;
wire n_17564;
wire n_17565;
wire n_17566;
wire n_17567;
wire n_17568;
wire n_17569;
wire n_1757;
wire n_17570;
wire n_17571;
wire n_17572;
wire n_17573;
wire n_17574;
wire n_17575;
wire n_17576;
wire n_17577;
wire n_17578;
wire n_17579;
wire n_1758;
wire n_17580;
wire n_17581;
wire n_17582;
wire n_17583;
wire n_17584;
wire n_17585;
wire n_17586;
wire n_17587;
wire n_17588;
wire n_17589;
wire n_1759;
wire n_17590;
wire n_17591;
wire n_17592;
wire n_17593;
wire n_17594;
wire n_17595;
wire n_17596;
wire n_17597;
wire n_17598;
wire n_17599;
wire n_176;
wire n_1760;
wire n_17600;
wire n_17601;
wire n_17602;
wire n_17603;
wire n_17604;
wire n_17605;
wire n_17606;
wire n_17607;
wire n_17608;
wire n_17609;
wire n_1761;
wire n_17610;
wire n_17611;
wire n_17612;
wire n_17613;
wire n_17614;
wire n_17615;
wire n_17616;
wire n_17617;
wire n_17618;
wire n_17619;
wire n_1762;
wire n_17620;
wire n_17621;
wire n_17622;
wire n_17623;
wire n_17624;
wire n_17625;
wire n_17626;
wire n_17627;
wire n_17628;
wire n_17629;
wire n_1763;
wire n_17630;
wire n_17631;
wire n_17632;
wire n_17633;
wire n_17634;
wire n_17635;
wire n_17636;
wire n_17637;
wire n_17638;
wire n_17639;
wire n_1764;
wire n_17640;
wire n_17641;
wire n_17642;
wire n_17643;
wire n_17644;
wire n_17645;
wire n_17646;
wire n_17647;
wire n_17648;
wire n_17649;
wire n_1765;
wire n_17650;
wire n_17651;
wire n_17652;
wire n_17653;
wire n_17654;
wire n_17655;
wire n_17656;
wire n_17657;
wire n_17658;
wire n_17659;
wire n_1766;
wire n_17660;
wire n_17661;
wire n_17662;
wire n_17663;
wire n_17664;
wire n_17665;
wire n_17666;
wire n_17667;
wire n_17668;
wire n_17669;
wire n_1767;
wire n_17670;
wire n_17671;
wire n_17672;
wire n_17673;
wire n_17674;
wire n_17675;
wire n_17676;
wire n_17677;
wire n_17678;
wire n_17679;
wire n_1768;
wire n_17680;
wire n_17681;
wire n_17682;
wire n_17683;
wire n_17684;
wire n_17685;
wire n_17686;
wire n_17687;
wire n_17688;
wire n_17689;
wire n_1769;
wire n_17690;
wire n_17691;
wire n_17692;
wire n_17693;
wire n_17694;
wire n_17695;
wire n_17696;
wire n_17697;
wire n_17698;
wire n_17699;
wire n_177;
wire n_1770;
wire n_17700;
wire n_17701;
wire n_17702;
wire n_17703;
wire n_17704;
wire n_17705;
wire n_17706;
wire n_17707;
wire n_17708;
wire n_17709;
wire n_1771;
wire n_17710;
wire n_17711;
wire n_17712;
wire n_17713;
wire n_17714;
wire n_17715;
wire n_17716;
wire n_17717;
wire n_17718;
wire n_17719;
wire n_1772;
wire n_17720;
wire n_17721;
wire n_17722;
wire n_17723;
wire n_17724;
wire n_17725;
wire n_17726;
wire n_17727;
wire n_17728;
wire n_17729;
wire n_1773;
wire n_17730;
wire n_17731;
wire n_17732;
wire n_17733;
wire n_17734;
wire n_17735;
wire n_17736;
wire n_17737;
wire n_17738;
wire n_17739;
wire n_1774;
wire n_17740;
wire n_17741;
wire n_17742;
wire n_17743;
wire n_17744;
wire n_17745;
wire n_17746;
wire n_17747;
wire n_17748;
wire n_17749;
wire n_1775;
wire n_17750;
wire n_17751;
wire n_17752;
wire n_17753;
wire n_17754;
wire n_17755;
wire n_17756;
wire n_17757;
wire n_17758;
wire n_17759;
wire n_1776;
wire n_17760;
wire n_17761;
wire n_17762;
wire n_17763;
wire n_17764;
wire n_17765;
wire n_17766;
wire n_17767;
wire n_17768;
wire n_17769;
wire n_1777;
wire n_17770;
wire n_17771;
wire n_17772;
wire n_17773;
wire n_17774;
wire n_17775;
wire n_17776;
wire n_17777;
wire n_17778;
wire n_17779;
wire n_1778;
wire n_17780;
wire n_17781;
wire n_17782;
wire n_17783;
wire n_17784;
wire n_17785;
wire n_17786;
wire n_17787;
wire n_17788;
wire n_17789;
wire n_1779;
wire n_17790;
wire n_17791;
wire n_17792;
wire n_17793;
wire n_17794;
wire n_17795;
wire n_17796;
wire n_17797;
wire n_17798;
wire n_17799;
wire n_178;
wire n_1780;
wire n_17800;
wire n_17801;
wire n_17802;
wire n_17803;
wire n_17804;
wire n_17805;
wire n_17806;
wire n_17807;
wire n_17808;
wire n_17809;
wire n_1781;
wire n_17810;
wire n_17811;
wire n_17812;
wire n_17813;
wire n_17814;
wire n_17815;
wire n_17816;
wire n_17817;
wire n_17818;
wire n_17819;
wire n_1782;
wire n_17820;
wire n_17821;
wire n_17822;
wire n_17823;
wire n_17824;
wire n_17825;
wire n_17826;
wire n_17827;
wire n_17828;
wire n_17829;
wire n_1783;
wire n_17830;
wire n_17831;
wire n_17832;
wire n_17833;
wire n_17834;
wire n_17835;
wire n_17836;
wire n_17837;
wire n_17838;
wire n_17839;
wire n_1784;
wire n_17840;
wire n_17841;
wire n_17843;
wire n_17844;
wire n_17845;
wire n_17846;
wire n_17847;
wire n_17848;
wire n_17849;
wire n_1785;
wire n_17850;
wire n_17851;
wire n_17852;
wire n_17853;
wire n_17854;
wire n_17855;
wire n_17856;
wire n_17857;
wire n_17858;
wire n_17859;
wire n_1786;
wire n_17860;
wire n_17861;
wire n_17862;
wire n_17863;
wire n_17864;
wire n_17865;
wire n_17866;
wire n_17867;
wire n_17868;
wire n_17869;
wire n_1787;
wire n_17870;
wire n_17871;
wire n_17872;
wire n_17873;
wire n_17874;
wire n_17875;
wire n_17876;
wire n_17877;
wire n_17878;
wire n_17879;
wire n_1788;
wire n_17880;
wire n_17881;
wire n_17882;
wire n_17883;
wire n_17884;
wire n_17885;
wire n_17886;
wire n_17887;
wire n_17888;
wire n_17889;
wire n_1789;
wire n_17890;
wire n_17891;
wire n_17892;
wire n_17893;
wire n_17894;
wire n_17895;
wire n_17896;
wire n_17897;
wire n_17898;
wire n_17899;
wire n_179;
wire n_1790;
wire n_17900;
wire n_17901;
wire n_17902;
wire n_17903;
wire n_17904;
wire n_17905;
wire n_17906;
wire n_17907;
wire n_17908;
wire n_17909;
wire n_1791;
wire n_17910;
wire n_17911;
wire n_17912;
wire n_17913;
wire n_17914;
wire n_17915;
wire n_17916;
wire n_17917;
wire n_17918;
wire n_17919;
wire n_1792;
wire n_17920;
wire n_17921;
wire n_17922;
wire n_17923;
wire n_17924;
wire n_17925;
wire n_17926;
wire n_17927;
wire n_17928;
wire n_17929;
wire n_1793;
wire n_17930;
wire n_17931;
wire n_17932;
wire n_17933;
wire n_17934;
wire n_17935;
wire n_17936;
wire n_17937;
wire n_17938;
wire n_17939;
wire n_1794;
wire n_17940;
wire n_17941;
wire n_17942;
wire n_17943;
wire n_17944;
wire n_17945;
wire n_17946;
wire n_17947;
wire n_17948;
wire n_17949;
wire n_1795;
wire n_17950;
wire n_17951;
wire n_17952;
wire n_17953;
wire n_17954;
wire n_17955;
wire n_17956;
wire n_17957;
wire n_17958;
wire n_17959;
wire n_1796;
wire n_17960;
wire n_17961;
wire n_17962;
wire n_17963;
wire n_17964;
wire n_17965;
wire n_17966;
wire n_17967;
wire n_17968;
wire n_17969;
wire n_1797;
wire n_17970;
wire n_17971;
wire n_17972;
wire n_17973;
wire n_17974;
wire n_17975;
wire n_17976;
wire n_17977;
wire n_17978;
wire n_17979;
wire n_1798;
wire n_17980;
wire n_17981;
wire n_17982;
wire n_17983;
wire n_17984;
wire n_17985;
wire n_17986;
wire n_17987;
wire n_17988;
wire n_17989;
wire n_1799;
wire n_17990;
wire n_17991;
wire n_17992;
wire n_17993;
wire n_17994;
wire n_17995;
wire n_17996;
wire n_17997;
wire n_17998;
wire n_17999;
wire n_18;
wire n_180;
wire n_1800;
wire n_18000;
wire n_18001;
wire n_18002;
wire n_18003;
wire n_18004;
wire n_18005;
wire n_18006;
wire n_18007;
wire n_18008;
wire n_18009;
wire n_1801;
wire n_18010;
wire n_18011;
wire n_18012;
wire n_18013;
wire n_18014;
wire n_18015;
wire n_18016;
wire n_18017;
wire n_18018;
wire n_18019;
wire n_1802;
wire n_18020;
wire n_18021;
wire n_18022;
wire n_18023;
wire n_18024;
wire n_18025;
wire n_18026;
wire n_18027;
wire n_18028;
wire n_18029;
wire n_1803;
wire n_18030;
wire n_18031;
wire n_18032;
wire n_18033;
wire n_18034;
wire n_18035;
wire n_18036;
wire n_18037;
wire n_18038;
wire n_18039;
wire n_1804;
wire n_18040;
wire n_18041;
wire n_18042;
wire n_18043;
wire n_18044;
wire n_18045;
wire n_18046;
wire n_18047;
wire n_18048;
wire n_18049;
wire n_1805;
wire n_18050;
wire n_18051;
wire n_18052;
wire n_18053;
wire n_18054;
wire n_18055;
wire n_18056;
wire n_18057;
wire n_18058;
wire n_18059;
wire n_1806;
wire n_18060;
wire n_18061;
wire n_18062;
wire n_18063;
wire n_18064;
wire n_18065;
wire n_18066;
wire n_18067;
wire n_18068;
wire n_18069;
wire n_1807;
wire n_18070;
wire n_18071;
wire n_18072;
wire n_18073;
wire n_18074;
wire n_18075;
wire n_18076;
wire n_18077;
wire n_18078;
wire n_18079;
wire n_1808;
wire n_18080;
wire n_18081;
wire n_18082;
wire n_18083;
wire n_18084;
wire n_18085;
wire n_18086;
wire n_18087;
wire n_18088;
wire n_18089;
wire n_1809;
wire n_18090;
wire n_18091;
wire n_18092;
wire n_18093;
wire n_18094;
wire n_18095;
wire n_18096;
wire n_18097;
wire n_18098;
wire n_18099;
wire n_181;
wire n_1810;
wire n_18100;
wire n_18101;
wire n_18102;
wire n_18103;
wire n_18104;
wire n_18105;
wire n_18106;
wire n_18107;
wire n_18108;
wire n_18109;
wire n_1811;
wire n_18110;
wire n_18111;
wire n_18112;
wire n_18113;
wire n_18114;
wire n_18115;
wire n_18116;
wire n_18117;
wire n_18118;
wire n_18119;
wire n_1812;
wire n_18120;
wire n_18121;
wire n_18122;
wire n_18123;
wire n_18124;
wire n_18125;
wire n_18126;
wire n_18127;
wire n_18128;
wire n_18129;
wire n_1813;
wire n_18130;
wire n_18131;
wire n_18132;
wire n_18133;
wire n_18134;
wire n_18135;
wire n_18136;
wire n_18137;
wire n_18138;
wire n_18139;
wire n_1814;
wire n_18140;
wire n_18141;
wire n_18142;
wire n_18143;
wire n_18144;
wire n_18145;
wire n_18146;
wire n_18147;
wire n_18148;
wire n_18149;
wire n_1815;
wire n_18150;
wire n_18151;
wire n_18152;
wire n_18153;
wire n_18154;
wire n_18155;
wire n_18156;
wire n_18157;
wire n_18158;
wire n_18159;
wire n_1816;
wire n_18160;
wire n_18161;
wire n_18162;
wire n_18163;
wire n_18164;
wire n_18165;
wire n_18166;
wire n_18167;
wire n_18168;
wire n_18169;
wire n_1817;
wire n_18170;
wire n_18171;
wire n_18172;
wire n_18173;
wire n_18174;
wire n_18175;
wire n_18176;
wire n_18177;
wire n_18178;
wire n_18179;
wire n_1818;
wire n_18180;
wire n_18181;
wire n_18182;
wire n_18183;
wire n_18184;
wire n_18185;
wire n_18186;
wire n_18187;
wire n_18188;
wire n_18189;
wire n_1819;
wire n_18190;
wire n_18191;
wire n_18192;
wire n_18193;
wire n_18194;
wire n_18195;
wire n_18196;
wire n_18197;
wire n_18198;
wire n_18199;
wire n_182;
wire n_1820;
wire n_18200;
wire n_18201;
wire n_18202;
wire n_18203;
wire n_18204;
wire n_18205;
wire n_18206;
wire n_18207;
wire n_18208;
wire n_18209;
wire n_1821;
wire n_18210;
wire n_18211;
wire n_18212;
wire n_18213;
wire n_18214;
wire n_18215;
wire n_18216;
wire n_18217;
wire n_18218;
wire n_18219;
wire n_1822;
wire n_18220;
wire n_18221;
wire n_18222;
wire n_18223;
wire n_18224;
wire n_18225;
wire n_18226;
wire n_18227;
wire n_18228;
wire n_18229;
wire n_1823;
wire n_18230;
wire n_18231;
wire n_18232;
wire n_18233;
wire n_18234;
wire n_18235;
wire n_18236;
wire n_18237;
wire n_18238;
wire n_18239;
wire n_1824;
wire n_18240;
wire n_18241;
wire n_18242;
wire n_18243;
wire n_18244;
wire n_18245;
wire n_18246;
wire n_18247;
wire n_18248;
wire n_18249;
wire n_1825;
wire n_18250;
wire n_18251;
wire n_18252;
wire n_18253;
wire n_18254;
wire n_18255;
wire n_18256;
wire n_18257;
wire n_18258;
wire n_18259;
wire n_1826;
wire n_18260;
wire n_18261;
wire n_18262;
wire n_18263;
wire n_18264;
wire n_18265;
wire n_18266;
wire n_18267;
wire n_18268;
wire n_18269;
wire n_1827;
wire n_18270;
wire n_18271;
wire n_18272;
wire n_18273;
wire n_18274;
wire n_18275;
wire n_18276;
wire n_18277;
wire n_18278;
wire n_18279;
wire n_1828;
wire n_18280;
wire n_18281;
wire n_18282;
wire n_18283;
wire n_18284;
wire n_18285;
wire n_18286;
wire n_18287;
wire n_18288;
wire n_18289;
wire n_1829;
wire n_18290;
wire n_18291;
wire n_18292;
wire n_18293;
wire n_18294;
wire n_18295;
wire n_18296;
wire n_18297;
wire n_18298;
wire n_18299;
wire n_183;
wire n_1830;
wire n_18300;
wire n_18301;
wire n_18302;
wire n_18303;
wire n_18304;
wire n_18305;
wire n_18306;
wire n_18307;
wire n_18308;
wire n_18309;
wire n_1831;
wire n_18310;
wire n_18311;
wire n_18312;
wire n_18313;
wire n_18314;
wire n_18315;
wire n_18316;
wire n_18317;
wire n_18318;
wire n_18319;
wire n_1832;
wire n_18320;
wire n_18321;
wire n_18322;
wire n_18323;
wire n_18324;
wire n_18325;
wire n_18326;
wire n_18327;
wire n_18328;
wire n_18329;
wire n_1833;
wire n_18330;
wire n_18331;
wire n_18332;
wire n_18333;
wire n_18334;
wire n_18335;
wire n_18336;
wire n_18337;
wire n_18338;
wire n_18339;
wire n_1834;
wire n_18340;
wire n_18341;
wire n_18342;
wire n_18343;
wire n_18344;
wire n_18345;
wire n_18346;
wire n_18347;
wire n_18348;
wire n_18349;
wire n_1835;
wire n_18350;
wire n_18351;
wire n_18352;
wire n_18353;
wire n_18354;
wire n_18355;
wire n_18356;
wire n_18357;
wire n_18358;
wire n_18359;
wire n_1836;
wire n_18360;
wire n_18361;
wire n_18362;
wire n_18363;
wire n_18364;
wire n_18365;
wire n_18366;
wire n_18367;
wire n_18368;
wire n_18369;
wire n_1837;
wire n_18370;
wire n_18371;
wire n_18372;
wire n_18373;
wire n_18374;
wire n_18375;
wire n_18376;
wire n_18377;
wire n_18378;
wire n_18379;
wire n_1838;
wire n_18380;
wire n_18381;
wire n_18382;
wire n_18383;
wire n_18384;
wire n_18385;
wire n_18386;
wire n_18387;
wire n_18388;
wire n_18389;
wire n_1839;
wire n_18390;
wire n_18391;
wire n_18392;
wire n_18393;
wire n_18394;
wire n_18395;
wire n_18396;
wire n_18397;
wire n_18398;
wire n_18399;
wire n_184;
wire n_1840;
wire n_18400;
wire n_18401;
wire n_18402;
wire n_18403;
wire n_18404;
wire n_18405;
wire n_18406;
wire n_18407;
wire n_18408;
wire n_18409;
wire n_1841;
wire n_18410;
wire n_18411;
wire n_18412;
wire n_18413;
wire n_18414;
wire n_18415;
wire n_18416;
wire n_18417;
wire n_18418;
wire n_18419;
wire n_1842;
wire n_18420;
wire n_18421;
wire n_18422;
wire n_18423;
wire n_18424;
wire n_18425;
wire n_18426;
wire n_18427;
wire n_18428;
wire n_18429;
wire n_1843;
wire n_18430;
wire n_18431;
wire n_18432;
wire n_18433;
wire n_18434;
wire n_18435;
wire n_18436;
wire n_18437;
wire n_18438;
wire n_18439;
wire n_1844;
wire n_18440;
wire n_18441;
wire n_18442;
wire n_18443;
wire n_18444;
wire n_18445;
wire n_18446;
wire n_18447;
wire n_18448;
wire n_18449;
wire n_1845;
wire n_18450;
wire n_18451;
wire n_18452;
wire n_18453;
wire n_18454;
wire n_18455;
wire n_18456;
wire n_18457;
wire n_18458;
wire n_18459;
wire n_1846;
wire n_18460;
wire n_18461;
wire n_18462;
wire n_18463;
wire n_18464;
wire n_18465;
wire n_18466;
wire n_18467;
wire n_18468;
wire n_18469;
wire n_1847;
wire n_18470;
wire n_18471;
wire n_18472;
wire n_18473;
wire n_18474;
wire n_18475;
wire n_18476;
wire n_18477;
wire n_18478;
wire n_18479;
wire n_1848;
wire n_18480;
wire n_18481;
wire n_18482;
wire n_18483;
wire n_18484;
wire n_18485;
wire n_18486;
wire n_18487;
wire n_18488;
wire n_18489;
wire n_1849;
wire n_18490;
wire n_18491;
wire n_18492;
wire n_18493;
wire n_18494;
wire n_18495;
wire n_18496;
wire n_18497;
wire n_18498;
wire n_18499;
wire n_185;
wire n_1850;
wire n_18500;
wire n_18501;
wire n_18502;
wire n_18503;
wire n_18504;
wire n_18505;
wire n_18506;
wire n_18507;
wire n_18508;
wire n_18509;
wire n_1851;
wire n_18510;
wire n_18511;
wire n_18512;
wire n_18513;
wire n_18514;
wire n_18515;
wire n_18516;
wire n_18517;
wire n_18518;
wire n_18519;
wire n_1852;
wire n_18520;
wire n_18522;
wire n_18523;
wire n_18524;
wire n_18526;
wire n_18527;
wire n_18528;
wire n_18529;
wire n_1853;
wire n_18530;
wire n_18531;
wire n_18532;
wire n_18533;
wire n_18534;
wire n_18535;
wire n_18536;
wire n_18537;
wire n_18538;
wire n_18539;
wire n_1854;
wire n_18540;
wire n_18541;
wire n_18542;
wire n_18543;
wire n_18544;
wire n_18545;
wire n_18546;
wire n_18547;
wire n_18548;
wire n_18549;
wire n_1855;
wire n_18550;
wire n_18551;
wire n_18552;
wire n_18553;
wire n_18554;
wire n_18555;
wire n_18556;
wire n_18557;
wire n_18558;
wire n_18559;
wire n_1856;
wire n_18560;
wire n_18561;
wire n_18562;
wire n_18563;
wire n_18564;
wire n_18565;
wire n_18566;
wire n_18567;
wire n_18568;
wire n_18569;
wire n_1857;
wire n_18570;
wire n_18571;
wire n_18572;
wire n_18573;
wire n_18574;
wire n_18575;
wire n_18576;
wire n_18577;
wire n_18578;
wire n_18579;
wire n_1858;
wire n_18580;
wire n_18581;
wire n_18582;
wire n_18583;
wire n_18584;
wire n_18585;
wire n_18586;
wire n_18587;
wire n_18588;
wire n_18589;
wire n_1859;
wire n_18590;
wire n_18591;
wire n_18592;
wire n_18593;
wire n_18594;
wire n_18595;
wire n_18596;
wire n_18597;
wire n_18598;
wire n_18599;
wire n_186;
wire n_1860;
wire n_18600;
wire n_18601;
wire n_18602;
wire n_18603;
wire n_18604;
wire n_18605;
wire n_18606;
wire n_18607;
wire n_18608;
wire n_18609;
wire n_1861;
wire n_18610;
wire n_18611;
wire n_18612;
wire n_18613;
wire n_18614;
wire n_18615;
wire n_18616;
wire n_18617;
wire n_18618;
wire n_18619;
wire n_1862;
wire n_18620;
wire n_18621;
wire n_18622;
wire n_18623;
wire n_18624;
wire n_18625;
wire n_18626;
wire n_18627;
wire n_18628;
wire n_18629;
wire n_1863;
wire n_18630;
wire n_18631;
wire n_18632;
wire n_18633;
wire n_18634;
wire n_18635;
wire n_18636;
wire n_18637;
wire n_18638;
wire n_18639;
wire n_1864;
wire n_18640;
wire n_18641;
wire n_18642;
wire n_18643;
wire n_18644;
wire n_18645;
wire n_18646;
wire n_18647;
wire n_18648;
wire n_18649;
wire n_1865;
wire n_18650;
wire n_18651;
wire n_18652;
wire n_18653;
wire n_18654;
wire n_18655;
wire n_18656;
wire n_18657;
wire n_18658;
wire n_18659;
wire n_1866;
wire n_18660;
wire n_18661;
wire n_18662;
wire n_18663;
wire n_18664;
wire n_18665;
wire n_18666;
wire n_18667;
wire n_18668;
wire n_18669;
wire n_1867;
wire n_18670;
wire n_18671;
wire n_18672;
wire n_18673;
wire n_18674;
wire n_18675;
wire n_18676;
wire n_18677;
wire n_18678;
wire n_18679;
wire n_1868;
wire n_18680;
wire n_18681;
wire n_18682;
wire n_18683;
wire n_18684;
wire n_18685;
wire n_18686;
wire n_18687;
wire n_18688;
wire n_18689;
wire n_1869;
wire n_18690;
wire n_18691;
wire n_18692;
wire n_18693;
wire n_18694;
wire n_18695;
wire n_18696;
wire n_18697;
wire n_18698;
wire n_18699;
wire n_187;
wire n_1870;
wire n_18700;
wire n_18701;
wire n_18702;
wire n_18703;
wire n_18704;
wire n_18705;
wire n_18706;
wire n_18707;
wire n_18708;
wire n_18709;
wire n_1871;
wire n_18710;
wire n_18711;
wire n_18712;
wire n_18713;
wire n_18714;
wire n_18715;
wire n_18716;
wire n_18717;
wire n_18718;
wire n_18719;
wire n_1872;
wire n_18720;
wire n_18721;
wire n_18722;
wire n_18723;
wire n_18724;
wire n_18725;
wire n_18726;
wire n_18727;
wire n_18728;
wire n_18729;
wire n_1873;
wire n_18730;
wire n_18731;
wire n_18732;
wire n_18733;
wire n_18734;
wire n_18735;
wire n_18736;
wire n_18737;
wire n_18738;
wire n_18739;
wire n_1874;
wire n_18740;
wire n_18741;
wire n_18742;
wire n_18743;
wire n_18744;
wire n_18745;
wire n_18746;
wire n_18747;
wire n_18748;
wire n_18749;
wire n_1875;
wire n_18750;
wire n_18751;
wire n_18752;
wire n_18753;
wire n_18754;
wire n_18755;
wire n_18756;
wire n_18757;
wire n_18758;
wire n_18759;
wire n_1876;
wire n_18760;
wire n_18761;
wire n_18762;
wire n_18763;
wire n_18764;
wire n_18765;
wire n_18766;
wire n_18767;
wire n_18768;
wire n_18769;
wire n_1877;
wire n_18770;
wire n_18771;
wire n_18772;
wire n_18773;
wire n_18774;
wire n_18775;
wire n_18776;
wire n_18777;
wire n_18778;
wire n_18779;
wire n_1878;
wire n_18780;
wire n_18781;
wire n_18782;
wire n_18783;
wire n_18784;
wire n_18785;
wire n_18786;
wire n_18787;
wire n_18788;
wire n_18789;
wire n_1879;
wire n_18790;
wire n_18791;
wire n_18792;
wire n_18793;
wire n_18794;
wire n_18795;
wire n_18796;
wire n_18797;
wire n_18798;
wire n_18799;
wire n_188;
wire n_1880;
wire n_18800;
wire n_18801;
wire n_18802;
wire n_18803;
wire n_18804;
wire n_18805;
wire n_18806;
wire n_18807;
wire n_18808;
wire n_18809;
wire n_1881;
wire n_18810;
wire n_18811;
wire n_18812;
wire n_18813;
wire n_18814;
wire n_18815;
wire n_18816;
wire n_18817;
wire n_18818;
wire n_18819;
wire n_1882;
wire n_18820;
wire n_18821;
wire n_18822;
wire n_18823;
wire n_18824;
wire n_18825;
wire n_18826;
wire n_18827;
wire n_18828;
wire n_18829;
wire n_1883;
wire n_18830;
wire n_18831;
wire n_18832;
wire n_18833;
wire n_18834;
wire n_18835;
wire n_18836;
wire n_18837;
wire n_18838;
wire n_18839;
wire n_1884;
wire n_18840;
wire n_18841;
wire n_18842;
wire n_18843;
wire n_18844;
wire n_18845;
wire n_18846;
wire n_18847;
wire n_18848;
wire n_18849;
wire n_1885;
wire n_18850;
wire n_18851;
wire n_18852;
wire n_18853;
wire n_18854;
wire n_18855;
wire n_18856;
wire n_18857;
wire n_18858;
wire n_18859;
wire n_1886;
wire n_18860;
wire n_18861;
wire n_18862;
wire n_18863;
wire n_18864;
wire n_18865;
wire n_18866;
wire n_18867;
wire n_18868;
wire n_18869;
wire n_1887;
wire n_18870;
wire n_18871;
wire n_18872;
wire n_18873;
wire n_18874;
wire n_18875;
wire n_18876;
wire n_18877;
wire n_18878;
wire n_18879;
wire n_1888;
wire n_18880;
wire n_18881;
wire n_18882;
wire n_18883;
wire n_18884;
wire n_18885;
wire n_18886;
wire n_18887;
wire n_18888;
wire n_18889;
wire n_1889;
wire n_18890;
wire n_18891;
wire n_18892;
wire n_18893;
wire n_18894;
wire n_18895;
wire n_18896;
wire n_18897;
wire n_18898;
wire n_18899;
wire n_189;
wire n_1890;
wire n_18900;
wire n_18901;
wire n_18902;
wire n_18903;
wire n_18904;
wire n_18905;
wire n_18906;
wire n_18907;
wire n_18908;
wire n_18909;
wire n_1891;
wire n_18910;
wire n_18911;
wire n_18912;
wire n_18913;
wire n_18914;
wire n_18915;
wire n_18916;
wire n_18917;
wire n_18918;
wire n_18919;
wire n_1892;
wire n_18920;
wire n_18921;
wire n_18922;
wire n_18923;
wire n_18924;
wire n_18925;
wire n_18926;
wire n_18927;
wire n_18928;
wire n_18929;
wire n_1893;
wire n_18930;
wire n_18931;
wire n_18932;
wire n_18933;
wire n_18934;
wire n_18935;
wire n_18936;
wire n_18937;
wire n_18938;
wire n_18939;
wire n_1894;
wire n_18940;
wire n_18941;
wire n_18942;
wire n_18943;
wire n_18944;
wire n_18945;
wire n_18946;
wire n_18947;
wire n_18948;
wire n_18949;
wire n_1895;
wire n_18950;
wire n_18951;
wire n_18952;
wire n_18953;
wire n_18954;
wire n_18955;
wire n_18956;
wire n_18957;
wire n_18958;
wire n_18959;
wire n_1896;
wire n_18960;
wire n_18961;
wire n_18962;
wire n_18963;
wire n_18964;
wire n_18965;
wire n_18966;
wire n_18967;
wire n_18968;
wire n_18969;
wire n_1897;
wire n_18970;
wire n_18971;
wire n_18972;
wire n_18973;
wire n_18974;
wire n_18975;
wire n_18976;
wire n_18977;
wire n_18978;
wire n_18979;
wire n_1898;
wire n_18980;
wire n_18981;
wire n_18982;
wire n_18983;
wire n_18984;
wire n_18985;
wire n_18986;
wire n_18987;
wire n_18988;
wire n_18989;
wire n_1899;
wire n_18990;
wire n_18991;
wire n_18992;
wire n_18993;
wire n_18994;
wire n_18995;
wire n_18996;
wire n_18997;
wire n_18998;
wire n_18999;
wire n_19;
wire n_190;
wire n_1900;
wire n_19000;
wire n_19001;
wire n_19002;
wire n_19003;
wire n_19004;
wire n_19005;
wire n_19006;
wire n_19007;
wire n_19008;
wire n_19009;
wire n_1901;
wire n_19010;
wire n_19011;
wire n_19012;
wire n_19013;
wire n_19014;
wire n_19015;
wire n_19016;
wire n_19017;
wire n_19018;
wire n_19019;
wire n_1902;
wire n_19020;
wire n_19021;
wire n_19022;
wire n_19023;
wire n_19024;
wire n_19025;
wire n_19026;
wire n_19027;
wire n_19028;
wire n_19029;
wire n_1903;
wire n_19030;
wire n_19031;
wire n_19032;
wire n_19033;
wire n_19034;
wire n_19035;
wire n_19036;
wire n_19037;
wire n_19038;
wire n_19039;
wire n_1904;
wire n_19040;
wire n_19041;
wire n_19042;
wire n_19043;
wire n_19044;
wire n_19045;
wire n_19046;
wire n_19047;
wire n_19048;
wire n_19049;
wire n_1905;
wire n_19050;
wire n_19051;
wire n_19052;
wire n_19053;
wire n_19054;
wire n_19055;
wire n_19056;
wire n_19057;
wire n_19058;
wire n_19059;
wire n_1906;
wire n_19060;
wire n_19061;
wire n_19062;
wire n_19063;
wire n_19064;
wire n_19065;
wire n_19066;
wire n_19067;
wire n_19068;
wire n_19069;
wire n_1907;
wire n_19070;
wire n_19071;
wire n_19072;
wire n_19073;
wire n_19074;
wire n_19075;
wire n_19076;
wire n_19077;
wire n_19078;
wire n_19079;
wire n_1908;
wire n_19080;
wire n_19081;
wire n_19082;
wire n_19083;
wire n_19084;
wire n_19085;
wire n_19086;
wire n_19087;
wire n_19088;
wire n_19089;
wire n_1909;
wire n_19090;
wire n_19091;
wire n_19092;
wire n_19093;
wire n_19094;
wire n_19095;
wire n_19096;
wire n_19097;
wire n_19098;
wire n_19099;
wire n_191;
wire n_1910;
wire n_19100;
wire n_19101;
wire n_19102;
wire n_19103;
wire n_19104;
wire n_19105;
wire n_19106;
wire n_19107;
wire n_19108;
wire n_19109;
wire n_1911;
wire n_19110;
wire n_19111;
wire n_19112;
wire n_19113;
wire n_19114;
wire n_19115;
wire n_19116;
wire n_19117;
wire n_19118;
wire n_19119;
wire n_1912;
wire n_19120;
wire n_19121;
wire n_19122;
wire n_19123;
wire n_19124;
wire n_19125;
wire n_19126;
wire n_19127;
wire n_19128;
wire n_19129;
wire n_1913;
wire n_19130;
wire n_19131;
wire n_19132;
wire n_19133;
wire n_19134;
wire n_19135;
wire n_19136;
wire n_19137;
wire n_19138;
wire n_19139;
wire n_1914;
wire n_19140;
wire n_19141;
wire n_19142;
wire n_19143;
wire n_19144;
wire n_19145;
wire n_19146;
wire n_19147;
wire n_19148;
wire n_19149;
wire n_1915;
wire n_19150;
wire n_19151;
wire n_19152;
wire n_19153;
wire n_19154;
wire n_19155;
wire n_19156;
wire n_19157;
wire n_19158;
wire n_19159;
wire n_1916;
wire n_19160;
wire n_19161;
wire n_19162;
wire n_19163;
wire n_19164;
wire n_19165;
wire n_19166;
wire n_19167;
wire n_19168;
wire n_19169;
wire n_1917;
wire n_19170;
wire n_19171;
wire n_19172;
wire n_19173;
wire n_19174;
wire n_19175;
wire n_19176;
wire n_19177;
wire n_19178;
wire n_19179;
wire n_1918;
wire n_19180;
wire n_19181;
wire n_19182;
wire n_19183;
wire n_19184;
wire n_19185;
wire n_19186;
wire n_19187;
wire n_19188;
wire n_19189;
wire n_1919;
wire n_19190;
wire n_19191;
wire n_19192;
wire n_19193;
wire n_19194;
wire n_19195;
wire n_19196;
wire n_19197;
wire n_19198;
wire n_19199;
wire n_192;
wire n_1920;
wire n_19200;
wire n_19201;
wire n_19202;
wire n_19203;
wire n_19204;
wire n_19205;
wire n_19206;
wire n_19207;
wire n_19208;
wire n_19209;
wire n_1921;
wire n_19210;
wire n_19211;
wire n_19212;
wire n_19213;
wire n_19214;
wire n_19215;
wire n_19216;
wire n_19217;
wire n_19218;
wire n_19219;
wire n_1922;
wire n_19220;
wire n_19221;
wire n_19222;
wire n_19223;
wire n_19224;
wire n_19225;
wire n_19226;
wire n_19227;
wire n_19228;
wire n_19229;
wire n_1923;
wire n_19230;
wire n_19231;
wire n_19232;
wire n_19233;
wire n_19234;
wire n_19235;
wire n_19236;
wire n_19237;
wire n_19238;
wire n_19239;
wire n_1924;
wire n_19240;
wire n_19241;
wire n_19242;
wire n_19243;
wire n_19244;
wire n_19245;
wire n_19246;
wire n_19247;
wire n_19248;
wire n_19249;
wire n_1925;
wire n_19250;
wire n_19251;
wire n_19252;
wire n_19253;
wire n_19254;
wire n_19255;
wire n_19256;
wire n_19257;
wire n_19258;
wire n_19259;
wire n_1926;
wire n_19260;
wire n_19261;
wire n_19262;
wire n_19263;
wire n_19264;
wire n_19265;
wire n_19266;
wire n_19267;
wire n_19268;
wire n_19269;
wire n_1927;
wire n_19270;
wire n_19271;
wire n_19272;
wire n_19273;
wire n_19274;
wire n_19275;
wire n_19276;
wire n_19277;
wire n_19278;
wire n_19279;
wire n_1928;
wire n_19280;
wire n_19281;
wire n_19282;
wire n_19283;
wire n_19284;
wire n_19285;
wire n_19286;
wire n_19287;
wire n_19288;
wire n_19289;
wire n_1929;
wire n_19290;
wire n_19291;
wire n_19292;
wire n_19293;
wire n_19294;
wire n_19295;
wire n_19296;
wire n_19297;
wire n_19298;
wire n_19299;
wire n_193;
wire n_1930;
wire n_19300;
wire n_19301;
wire n_19302;
wire n_19303;
wire n_19304;
wire n_19305;
wire n_19306;
wire n_19307;
wire n_19308;
wire n_19309;
wire n_1931;
wire n_19310;
wire n_19311;
wire n_19312;
wire n_19313;
wire n_19314;
wire n_19315;
wire n_19316;
wire n_19317;
wire n_19318;
wire n_19319;
wire n_1932;
wire n_19320;
wire n_19321;
wire n_19322;
wire n_19323;
wire n_19324;
wire n_19325;
wire n_19326;
wire n_19327;
wire n_19328;
wire n_19329;
wire n_1933;
wire n_19330;
wire n_19331;
wire n_19332;
wire n_19333;
wire n_19334;
wire n_19335;
wire n_19336;
wire n_19337;
wire n_19338;
wire n_19339;
wire n_1934;
wire n_19340;
wire n_19341;
wire n_19342;
wire n_19343;
wire n_19344;
wire n_19345;
wire n_19346;
wire n_19347;
wire n_19348;
wire n_19349;
wire n_1935;
wire n_19350;
wire n_19351;
wire n_19352;
wire n_19353;
wire n_19354;
wire n_19355;
wire n_19356;
wire n_19357;
wire n_19358;
wire n_19359;
wire n_1936;
wire n_19360;
wire n_19361;
wire n_19362;
wire n_19363;
wire n_19364;
wire n_19365;
wire n_19366;
wire n_19367;
wire n_19368;
wire n_19369;
wire n_1937;
wire n_19370;
wire n_19371;
wire n_19372;
wire n_19373;
wire n_19374;
wire n_19375;
wire n_19376;
wire n_19377;
wire n_19378;
wire n_19379;
wire n_1938;
wire n_19380;
wire n_19381;
wire n_19382;
wire n_19383;
wire n_19384;
wire n_19385;
wire n_19386;
wire n_19387;
wire n_19388;
wire n_19389;
wire n_1939;
wire n_19390;
wire n_19391;
wire n_19392;
wire n_19393;
wire n_19394;
wire n_19395;
wire n_19396;
wire n_19397;
wire n_19398;
wire n_19399;
wire n_194;
wire n_1940;
wire n_19400;
wire n_19401;
wire n_19402;
wire n_19403;
wire n_19404;
wire n_19405;
wire n_19406;
wire n_19407;
wire n_19408;
wire n_19409;
wire n_1941;
wire n_19410;
wire n_19411;
wire n_19412;
wire n_19413;
wire n_19414;
wire n_19415;
wire n_19416;
wire n_19417;
wire n_19418;
wire n_19419;
wire n_1942;
wire n_19420;
wire n_19421;
wire n_19422;
wire n_19423;
wire n_19424;
wire n_19425;
wire n_19426;
wire n_19427;
wire n_19428;
wire n_19429;
wire n_1943;
wire n_19430;
wire n_19431;
wire n_19432;
wire n_19433;
wire n_19434;
wire n_19435;
wire n_19436;
wire n_19437;
wire n_19438;
wire n_19439;
wire n_1944;
wire n_19440;
wire n_19441;
wire n_19442;
wire n_19443;
wire n_19444;
wire n_19445;
wire n_19446;
wire n_19447;
wire n_19448;
wire n_19449;
wire n_1945;
wire n_19450;
wire n_19451;
wire n_19452;
wire n_19453;
wire n_19454;
wire n_19455;
wire n_19456;
wire n_19457;
wire n_19458;
wire n_19459;
wire n_1946;
wire n_19460;
wire n_19461;
wire n_19462;
wire n_19463;
wire n_19464;
wire n_19465;
wire n_19466;
wire n_19467;
wire n_19468;
wire n_19469;
wire n_1947;
wire n_19470;
wire n_19471;
wire n_19472;
wire n_19473;
wire n_19474;
wire n_19475;
wire n_19476;
wire n_19477;
wire n_19478;
wire n_19479;
wire n_1948;
wire n_19480;
wire n_19481;
wire n_19482;
wire n_19483;
wire n_19484;
wire n_19485;
wire n_19486;
wire n_19487;
wire n_19488;
wire n_19489;
wire n_1949;
wire n_19490;
wire n_19491;
wire n_19492;
wire n_19493;
wire n_19494;
wire n_19495;
wire n_19496;
wire n_19497;
wire n_19498;
wire n_19499;
wire n_195;
wire n_1950;
wire n_19500;
wire n_19501;
wire n_19502;
wire n_19503;
wire n_19504;
wire n_19505;
wire n_19506;
wire n_19507;
wire n_19508;
wire n_19509;
wire n_1951;
wire n_19510;
wire n_19511;
wire n_19512;
wire n_19513;
wire n_19514;
wire n_19515;
wire n_19516;
wire n_19517;
wire n_19518;
wire n_19519;
wire n_1952;
wire n_19520;
wire n_19521;
wire n_19522;
wire n_19523;
wire n_19524;
wire n_19525;
wire n_19526;
wire n_19527;
wire n_19528;
wire n_19529;
wire n_1953;
wire n_19530;
wire n_19531;
wire n_19532;
wire n_19533;
wire n_19534;
wire n_19535;
wire n_19536;
wire n_19537;
wire n_19538;
wire n_19539;
wire n_1954;
wire n_19540;
wire n_19541;
wire n_19542;
wire n_19543;
wire n_19544;
wire n_19545;
wire n_19546;
wire n_19547;
wire n_19548;
wire n_19549;
wire n_1955;
wire n_19550;
wire n_19551;
wire n_19552;
wire n_19553;
wire n_19554;
wire n_19555;
wire n_19556;
wire n_19557;
wire n_19558;
wire n_19559;
wire n_1956;
wire n_19560;
wire n_19561;
wire n_19562;
wire n_19563;
wire n_19564;
wire n_19565;
wire n_19566;
wire n_19567;
wire n_19568;
wire n_19569;
wire n_1957;
wire n_19570;
wire n_19571;
wire n_19572;
wire n_19573;
wire n_19574;
wire n_19575;
wire n_19576;
wire n_19577;
wire n_19578;
wire n_19579;
wire n_1958;
wire n_19580;
wire n_19581;
wire n_19582;
wire n_19583;
wire n_19584;
wire n_19585;
wire n_19586;
wire n_19587;
wire n_19588;
wire n_19589;
wire n_1959;
wire n_19590;
wire n_19591;
wire n_19592;
wire n_19593;
wire n_19594;
wire n_19595;
wire n_19596;
wire n_19597;
wire n_19598;
wire n_19599;
wire n_196;
wire n_1960;
wire n_19600;
wire n_19601;
wire n_19602;
wire n_19603;
wire n_19604;
wire n_19605;
wire n_19606;
wire n_19607;
wire n_19608;
wire n_19609;
wire n_1961;
wire n_19610;
wire n_19611;
wire n_19612;
wire n_19613;
wire n_19614;
wire n_19615;
wire n_19616;
wire n_19617;
wire n_19618;
wire n_19619;
wire n_1962;
wire n_19620;
wire n_19621;
wire n_19622;
wire n_19623;
wire n_19624;
wire n_19625;
wire n_19626;
wire n_19627;
wire n_19628;
wire n_19629;
wire n_1963;
wire n_19630;
wire n_19631;
wire n_19632;
wire n_19633;
wire n_19634;
wire n_19635;
wire n_19636;
wire n_19637;
wire n_19638;
wire n_19639;
wire n_1964;
wire n_19640;
wire n_19641;
wire n_19642;
wire n_19643;
wire n_19644;
wire n_19645;
wire n_19646;
wire n_19647;
wire n_19648;
wire n_19649;
wire n_1965;
wire n_19650;
wire n_19651;
wire n_19652;
wire n_19653;
wire n_19654;
wire n_19655;
wire n_19656;
wire n_19657;
wire n_19658;
wire n_19659;
wire n_1966;
wire n_19660;
wire n_19661;
wire n_19662;
wire n_19663;
wire n_19664;
wire n_19665;
wire n_19666;
wire n_19667;
wire n_19668;
wire n_19669;
wire n_1967;
wire n_19670;
wire n_19671;
wire n_19672;
wire n_19673;
wire n_19674;
wire n_19675;
wire n_19676;
wire n_19677;
wire n_19678;
wire n_19679;
wire n_1968;
wire n_19680;
wire n_19681;
wire n_19682;
wire n_19683;
wire n_19684;
wire n_19685;
wire n_19686;
wire n_19687;
wire n_19688;
wire n_19689;
wire n_1969;
wire n_19690;
wire n_19691;
wire n_19692;
wire n_19693;
wire n_19694;
wire n_19695;
wire n_19696;
wire n_19697;
wire n_19698;
wire n_19699;
wire n_197;
wire n_1970;
wire n_19700;
wire n_19701;
wire n_19702;
wire n_19703;
wire n_19704;
wire n_19705;
wire n_19706;
wire n_19707;
wire n_19708;
wire n_19709;
wire n_1971;
wire n_19710;
wire n_19711;
wire n_19712;
wire n_19713;
wire n_19714;
wire n_19715;
wire n_19716;
wire n_19717;
wire n_19718;
wire n_19719;
wire n_1972;
wire n_19720;
wire n_19721;
wire n_19722;
wire n_19723;
wire n_19724;
wire n_19725;
wire n_19726;
wire n_19727;
wire n_19728;
wire n_19729;
wire n_1973;
wire n_19730;
wire n_19731;
wire n_19732;
wire n_19733;
wire n_19734;
wire n_19735;
wire n_19736;
wire n_19737;
wire n_19738;
wire n_19739;
wire n_1974;
wire n_19740;
wire n_19741;
wire n_19742;
wire n_19743;
wire n_19744;
wire n_19745;
wire n_19746;
wire n_19747;
wire n_19748;
wire n_19749;
wire n_1975;
wire n_19750;
wire n_19751;
wire n_19752;
wire n_19753;
wire n_19754;
wire n_19755;
wire n_19756;
wire n_19757;
wire n_19758;
wire n_19759;
wire n_1976;
wire n_19760;
wire n_19761;
wire n_19762;
wire n_19763;
wire n_19764;
wire n_19765;
wire n_19766;
wire n_19767;
wire n_19768;
wire n_19769;
wire n_1977;
wire n_19770;
wire n_19771;
wire n_19772;
wire n_19773;
wire n_19774;
wire n_19775;
wire n_19776;
wire n_19777;
wire n_19778;
wire n_19779;
wire n_1978;
wire n_19780;
wire n_19781;
wire n_19782;
wire n_19783;
wire n_19784;
wire n_19785;
wire n_19786;
wire n_19787;
wire n_19788;
wire n_19789;
wire n_1979;
wire n_19790;
wire n_19791;
wire n_19792;
wire n_19793;
wire n_19794;
wire n_19795;
wire n_19796;
wire n_19797;
wire n_19798;
wire n_19799;
wire n_198;
wire n_1980;
wire n_19800;
wire n_19801;
wire n_19802;
wire n_19803;
wire n_19804;
wire n_19805;
wire n_19806;
wire n_19807;
wire n_19808;
wire n_19809;
wire n_1981;
wire n_19810;
wire n_19811;
wire n_19812;
wire n_19813;
wire n_19814;
wire n_19815;
wire n_19816;
wire n_19817;
wire n_19818;
wire n_19819;
wire n_1982;
wire n_19820;
wire n_19821;
wire n_19822;
wire n_19823;
wire n_19824;
wire n_19825;
wire n_19826;
wire n_19827;
wire n_19828;
wire n_19829;
wire n_19830;
wire n_19831;
wire n_19832;
wire n_19833;
wire n_19834;
wire n_19835;
wire n_19836;
wire n_19837;
wire n_19838;
wire n_19839;
wire n_1984;
wire n_19840;
wire n_19841;
wire n_19842;
wire n_19843;
wire n_19844;
wire n_19845;
wire n_19846;
wire n_19847;
wire n_19848;
wire n_19849;
wire n_1985;
wire n_19850;
wire n_19851;
wire n_19852;
wire n_19853;
wire n_19854;
wire n_19855;
wire n_19856;
wire n_19857;
wire n_19858;
wire n_19859;
wire n_1986;
wire n_19860;
wire n_19861;
wire n_19862;
wire n_19863;
wire n_19864;
wire n_19865;
wire n_19866;
wire n_19867;
wire n_19868;
wire n_19869;
wire n_1987;
wire n_19870;
wire n_19871;
wire n_19872;
wire n_19873;
wire n_19874;
wire n_19875;
wire n_19876;
wire n_19877;
wire n_19878;
wire n_19879;
wire n_1988;
wire n_19880;
wire n_19881;
wire n_19882;
wire n_19883;
wire n_19884;
wire n_19885;
wire n_19886;
wire n_19887;
wire n_19888;
wire n_19889;
wire n_1989;
wire n_19890;
wire n_19891;
wire n_19892;
wire n_19893;
wire n_19894;
wire n_19895;
wire n_19896;
wire n_19897;
wire n_19898;
wire n_19899;
wire n_199;
wire n_1990;
wire n_19900;
wire n_19901;
wire n_19902;
wire n_19903;
wire n_19904;
wire n_19905;
wire n_19906;
wire n_19907;
wire n_19908;
wire n_19909;
wire n_1991;
wire n_19910;
wire n_19911;
wire n_19912;
wire n_19913;
wire n_19914;
wire n_19915;
wire n_19916;
wire n_19918;
wire n_19919;
wire n_1992;
wire n_19920;
wire n_19921;
wire n_19922;
wire n_19923;
wire n_19924;
wire n_19925;
wire n_19926;
wire n_19927;
wire n_19928;
wire n_19929;
wire n_1993;
wire n_19930;
wire n_19931;
wire n_19932;
wire n_19933;
wire n_19934;
wire n_19935;
wire n_19936;
wire n_19937;
wire n_19938;
wire n_19939;
wire n_1994;
wire n_19940;
wire n_19941;
wire n_19942;
wire n_19943;
wire n_19944;
wire n_19945;
wire n_19946;
wire n_19947;
wire n_19948;
wire n_19949;
wire n_1995;
wire n_19950;
wire n_19951;
wire n_19952;
wire n_19953;
wire n_19954;
wire n_19955;
wire n_19956;
wire n_19957;
wire n_19958;
wire n_19959;
wire n_1996;
wire n_19960;
wire n_19961;
wire n_19962;
wire n_19963;
wire n_19964;
wire n_19965;
wire n_19966;
wire n_19967;
wire n_19968;
wire n_19969;
wire n_1997;
wire n_19970;
wire n_19971;
wire n_19972;
wire n_19973;
wire n_19974;
wire n_19975;
wire n_19976;
wire n_19977;
wire n_19978;
wire n_19979;
wire n_1998;
wire n_19980;
wire n_19981;
wire n_19982;
wire n_19983;
wire n_19984;
wire n_19985;
wire n_19986;
wire n_19987;
wire n_19988;
wire n_19989;
wire n_1999;
wire n_19990;
wire n_19991;
wire n_19992;
wire n_19993;
wire n_19994;
wire n_19995;
wire n_19996;
wire n_19997;
wire n_19998;
wire n_19999;
wire n_2;
wire n_20;
wire n_200;
wire n_2000;
wire n_20000;
wire n_20001;
wire n_20002;
wire n_20003;
wire n_20004;
wire n_20005;
wire n_20006;
wire n_20007;
wire n_20008;
wire n_20009;
wire n_2001;
wire n_20010;
wire n_20011;
wire n_20012;
wire n_20013;
wire n_20014;
wire n_20015;
wire n_20016;
wire n_20017;
wire n_20018;
wire n_20019;
wire n_2002;
wire n_20020;
wire n_20021;
wire n_20022;
wire n_20023;
wire n_20024;
wire n_20025;
wire n_20026;
wire n_20027;
wire n_20028;
wire n_20029;
wire n_2003;
wire n_20030;
wire n_20031;
wire n_20032;
wire n_20033;
wire n_20034;
wire n_20035;
wire n_20036;
wire n_20037;
wire n_20038;
wire n_20039;
wire n_2004;
wire n_20040;
wire n_20041;
wire n_20042;
wire n_20043;
wire n_20044;
wire n_20045;
wire n_20046;
wire n_20047;
wire n_20048;
wire n_20049;
wire n_2005;
wire n_20050;
wire n_20051;
wire n_20052;
wire n_20053;
wire n_20054;
wire n_20055;
wire n_20056;
wire n_20057;
wire n_20058;
wire n_20059;
wire n_2006;
wire n_20060;
wire n_20061;
wire n_20062;
wire n_20063;
wire n_20064;
wire n_20065;
wire n_20066;
wire n_20067;
wire n_20068;
wire n_20069;
wire n_2007;
wire n_20070;
wire n_20071;
wire n_20072;
wire n_20073;
wire n_20074;
wire n_20075;
wire n_20076;
wire n_20077;
wire n_20078;
wire n_20079;
wire n_2008;
wire n_20080;
wire n_20081;
wire n_20082;
wire n_20083;
wire n_20084;
wire n_20085;
wire n_20086;
wire n_20087;
wire n_20088;
wire n_20089;
wire n_2009;
wire n_20090;
wire n_20091;
wire n_20092;
wire n_20093;
wire n_20094;
wire n_20095;
wire n_20096;
wire n_20097;
wire n_20098;
wire n_20099;
wire n_201;
wire n_2010;
wire n_20100;
wire n_20101;
wire n_20102;
wire n_20103;
wire n_20104;
wire n_20105;
wire n_20106;
wire n_20107;
wire n_20108;
wire n_20109;
wire n_2011;
wire n_20110;
wire n_20111;
wire n_20112;
wire n_20113;
wire n_20114;
wire n_20115;
wire n_20116;
wire n_20117;
wire n_20118;
wire n_20119;
wire n_2012;
wire n_20120;
wire n_20121;
wire n_20122;
wire n_20123;
wire n_20124;
wire n_20125;
wire n_20126;
wire n_20127;
wire n_20128;
wire n_20129;
wire n_2013;
wire n_20130;
wire n_20131;
wire n_20132;
wire n_20133;
wire n_20134;
wire n_20135;
wire n_20136;
wire n_20137;
wire n_20138;
wire n_20139;
wire n_20140;
wire n_20141;
wire n_20142;
wire n_20143;
wire n_20144;
wire n_20145;
wire n_20146;
wire n_20147;
wire n_20148;
wire n_20149;
wire n_2015;
wire n_20150;
wire n_20151;
wire n_20152;
wire n_20153;
wire n_20154;
wire n_20155;
wire n_20156;
wire n_20157;
wire n_20158;
wire n_20159;
wire n_2016;
wire n_20160;
wire n_20161;
wire n_20162;
wire n_20163;
wire n_20164;
wire n_20165;
wire n_20166;
wire n_20167;
wire n_20168;
wire n_20169;
wire n_2017;
wire n_20170;
wire n_20171;
wire n_20172;
wire n_20173;
wire n_20174;
wire n_20175;
wire n_20176;
wire n_20177;
wire n_20178;
wire n_20179;
wire n_2018;
wire n_20180;
wire n_20181;
wire n_20182;
wire n_20183;
wire n_20184;
wire n_20185;
wire n_20186;
wire n_20187;
wire n_20188;
wire n_20189;
wire n_2019;
wire n_20190;
wire n_20191;
wire n_20192;
wire n_20193;
wire n_20194;
wire n_20195;
wire n_20196;
wire n_20197;
wire n_20198;
wire n_20199;
wire n_202;
wire n_2020;
wire n_20200;
wire n_20201;
wire n_20202;
wire n_20203;
wire n_20204;
wire n_20205;
wire n_20206;
wire n_20207;
wire n_20208;
wire n_20209;
wire n_2021;
wire n_20210;
wire n_20211;
wire n_20212;
wire n_20213;
wire n_20214;
wire n_20215;
wire n_20216;
wire n_20217;
wire n_20218;
wire n_20219;
wire n_2022;
wire n_20220;
wire n_20221;
wire n_20222;
wire n_20223;
wire n_20224;
wire n_20225;
wire n_20226;
wire n_20227;
wire n_20228;
wire n_20229;
wire n_2023;
wire n_20230;
wire n_20231;
wire n_20232;
wire n_20233;
wire n_20234;
wire n_20235;
wire n_20236;
wire n_20237;
wire n_20238;
wire n_20239;
wire n_2024;
wire n_20240;
wire n_20241;
wire n_20242;
wire n_20243;
wire n_20244;
wire n_20245;
wire n_20246;
wire n_20247;
wire n_20248;
wire n_20249;
wire n_2025;
wire n_20250;
wire n_20251;
wire n_20252;
wire n_20253;
wire n_20254;
wire n_20255;
wire n_20256;
wire n_20257;
wire n_20258;
wire n_20259;
wire n_2026;
wire n_20260;
wire n_20261;
wire n_20262;
wire n_20263;
wire n_20264;
wire n_20265;
wire n_20266;
wire n_20267;
wire n_20268;
wire n_20269;
wire n_2027;
wire n_20270;
wire n_20271;
wire n_20272;
wire n_20273;
wire n_20274;
wire n_20275;
wire n_20276;
wire n_20277;
wire n_20278;
wire n_20279;
wire n_2028;
wire n_20280;
wire n_20281;
wire n_20282;
wire n_20283;
wire n_20284;
wire n_20285;
wire n_20286;
wire n_20287;
wire n_20288;
wire n_20289;
wire n_2029;
wire n_20290;
wire n_20291;
wire n_20292;
wire n_20293;
wire n_20294;
wire n_20295;
wire n_20296;
wire n_20297;
wire n_20298;
wire n_20299;
wire n_203;
wire n_2030;
wire n_20300;
wire n_20301;
wire n_20302;
wire n_20303;
wire n_20304;
wire n_20305;
wire n_20306;
wire n_20307;
wire n_20308;
wire n_20309;
wire n_2031;
wire n_20310;
wire n_20311;
wire n_20312;
wire n_20313;
wire n_20314;
wire n_20315;
wire n_20316;
wire n_20317;
wire n_20318;
wire n_20319;
wire n_2032;
wire n_20320;
wire n_20321;
wire n_20322;
wire n_20323;
wire n_20324;
wire n_20325;
wire n_20326;
wire n_20327;
wire n_20328;
wire n_20329;
wire n_2033;
wire n_20330;
wire n_20331;
wire n_20332;
wire n_20333;
wire n_20334;
wire n_20335;
wire n_20336;
wire n_20337;
wire n_20338;
wire n_20339;
wire n_2034;
wire n_20340;
wire n_20341;
wire n_20342;
wire n_20343;
wire n_20344;
wire n_20345;
wire n_20346;
wire n_20347;
wire n_20348;
wire n_20349;
wire n_2035;
wire n_20350;
wire n_20351;
wire n_20352;
wire n_20353;
wire n_20354;
wire n_20355;
wire n_20356;
wire n_20357;
wire n_20358;
wire n_20359;
wire n_2036;
wire n_20360;
wire n_20361;
wire n_20362;
wire n_20363;
wire n_20364;
wire n_20365;
wire n_20366;
wire n_20367;
wire n_20368;
wire n_20369;
wire n_2037;
wire n_20370;
wire n_20371;
wire n_20372;
wire n_20373;
wire n_20374;
wire n_20375;
wire n_20376;
wire n_20377;
wire n_20378;
wire n_20379;
wire n_2038;
wire n_20380;
wire n_20381;
wire n_20382;
wire n_20383;
wire n_20384;
wire n_20385;
wire n_20386;
wire n_20387;
wire n_20388;
wire n_20389;
wire n_2039;
wire n_20390;
wire n_20391;
wire n_20392;
wire n_20393;
wire n_20394;
wire n_20395;
wire n_20396;
wire n_20397;
wire n_20398;
wire n_20399;
wire n_204;
wire n_2040;
wire n_20400;
wire n_20401;
wire n_20402;
wire n_20403;
wire n_20404;
wire n_20405;
wire n_20406;
wire n_20407;
wire n_20408;
wire n_20409;
wire n_2041;
wire n_20410;
wire n_20411;
wire n_20412;
wire n_20413;
wire n_20414;
wire n_20415;
wire n_20416;
wire n_20417;
wire n_20418;
wire n_20419;
wire n_2042;
wire n_20420;
wire n_20421;
wire n_20422;
wire n_20423;
wire n_20424;
wire n_20425;
wire n_20426;
wire n_20427;
wire n_20428;
wire n_20429;
wire n_2043;
wire n_20430;
wire n_20431;
wire n_20432;
wire n_20433;
wire n_20434;
wire n_20435;
wire n_20436;
wire n_20437;
wire n_20438;
wire n_20439;
wire n_2044;
wire n_20440;
wire n_20441;
wire n_20442;
wire n_20443;
wire n_20444;
wire n_20445;
wire n_20446;
wire n_20447;
wire n_20448;
wire n_20449;
wire n_2045;
wire n_20450;
wire n_20451;
wire n_20452;
wire n_20453;
wire n_20454;
wire n_20455;
wire n_20456;
wire n_20457;
wire n_20458;
wire n_20459;
wire n_2046;
wire n_20460;
wire n_20461;
wire n_20462;
wire n_20463;
wire n_20464;
wire n_20465;
wire n_20466;
wire n_20467;
wire n_20468;
wire n_20469;
wire n_2047;
wire n_20470;
wire n_20471;
wire n_20472;
wire n_20473;
wire n_20474;
wire n_20475;
wire n_20476;
wire n_20477;
wire n_20478;
wire n_20479;
wire n_2048;
wire n_20480;
wire n_20481;
wire n_20482;
wire n_20483;
wire n_20484;
wire n_20485;
wire n_20486;
wire n_20487;
wire n_20488;
wire n_20489;
wire n_2049;
wire n_20490;
wire n_20491;
wire n_20492;
wire n_20493;
wire n_20494;
wire n_20495;
wire n_20496;
wire n_20497;
wire n_20498;
wire n_20499;
wire n_205;
wire n_2050;
wire n_20500;
wire n_20501;
wire n_20502;
wire n_20503;
wire n_20504;
wire n_20505;
wire n_20506;
wire n_20507;
wire n_20508;
wire n_20509;
wire n_2051;
wire n_20510;
wire n_20511;
wire n_20512;
wire n_20513;
wire n_20514;
wire n_20515;
wire n_20516;
wire n_20517;
wire n_20518;
wire n_20519;
wire n_2052;
wire n_20520;
wire n_20521;
wire n_20522;
wire n_20523;
wire n_20524;
wire n_20525;
wire n_20526;
wire n_20527;
wire n_20528;
wire n_20529;
wire n_2053;
wire n_20530;
wire n_20531;
wire n_20532;
wire n_20533;
wire n_20534;
wire n_20536;
wire n_20538;
wire n_20539;
wire n_2054;
wire n_20540;
wire n_20541;
wire n_20542;
wire n_20543;
wire n_20544;
wire n_20545;
wire n_20546;
wire n_20547;
wire n_20548;
wire n_20549;
wire n_2055;
wire n_20550;
wire n_20551;
wire n_20552;
wire n_20553;
wire n_20554;
wire n_20555;
wire n_20556;
wire n_20557;
wire n_20558;
wire n_20559;
wire n_2056;
wire n_20560;
wire n_20561;
wire n_20562;
wire n_20563;
wire n_20564;
wire n_20565;
wire n_20566;
wire n_20567;
wire n_20568;
wire n_20569;
wire n_2057;
wire n_20570;
wire n_20571;
wire n_20572;
wire n_20573;
wire n_20574;
wire n_20575;
wire n_20576;
wire n_20577;
wire n_20578;
wire n_20579;
wire n_2058;
wire n_20580;
wire n_20581;
wire n_20582;
wire n_20583;
wire n_20584;
wire n_20585;
wire n_20586;
wire n_20587;
wire n_20588;
wire n_20589;
wire n_2059;
wire n_20590;
wire n_20591;
wire n_20592;
wire n_20593;
wire n_20594;
wire n_20595;
wire n_20596;
wire n_20597;
wire n_20598;
wire n_20599;
wire n_206;
wire n_2060;
wire n_20600;
wire n_20601;
wire n_20602;
wire n_20603;
wire n_20604;
wire n_20605;
wire n_20606;
wire n_20607;
wire n_20608;
wire n_20609;
wire n_2061;
wire n_20610;
wire n_20611;
wire n_20612;
wire n_20613;
wire n_20614;
wire n_20615;
wire n_20616;
wire n_20617;
wire n_20618;
wire n_20619;
wire n_2062;
wire n_20620;
wire n_20621;
wire n_20622;
wire n_20623;
wire n_20624;
wire n_20625;
wire n_20626;
wire n_20627;
wire n_20628;
wire n_20629;
wire n_2063;
wire n_20630;
wire n_20631;
wire n_20632;
wire n_20633;
wire n_20634;
wire n_20635;
wire n_20636;
wire n_20637;
wire n_20638;
wire n_20639;
wire n_2064;
wire n_20640;
wire n_20641;
wire n_20642;
wire n_20643;
wire n_20644;
wire n_20645;
wire n_20646;
wire n_20647;
wire n_20648;
wire n_20649;
wire n_2065;
wire n_20650;
wire n_20651;
wire n_20652;
wire n_20653;
wire n_20654;
wire n_20655;
wire n_20656;
wire n_20657;
wire n_20658;
wire n_20659;
wire n_2066;
wire n_20660;
wire n_20661;
wire n_20662;
wire n_20663;
wire n_20664;
wire n_20665;
wire n_20666;
wire n_20667;
wire n_20668;
wire n_20669;
wire n_2067;
wire n_20670;
wire n_20671;
wire n_20672;
wire n_20673;
wire n_20674;
wire n_20675;
wire n_20676;
wire n_20677;
wire n_20678;
wire n_20679;
wire n_2068;
wire n_20680;
wire n_20681;
wire n_20682;
wire n_20683;
wire n_20684;
wire n_20685;
wire n_20686;
wire n_20687;
wire n_20688;
wire n_20689;
wire n_2069;
wire n_20690;
wire n_20691;
wire n_20692;
wire n_20693;
wire n_20694;
wire n_20695;
wire n_20696;
wire n_20697;
wire n_20698;
wire n_20699;
wire n_207;
wire n_2070;
wire n_20700;
wire n_20701;
wire n_20702;
wire n_20703;
wire n_20704;
wire n_20705;
wire n_20706;
wire n_20707;
wire n_20708;
wire n_20709;
wire n_2071;
wire n_20710;
wire n_20711;
wire n_20712;
wire n_20713;
wire n_20714;
wire n_20715;
wire n_20716;
wire n_20717;
wire n_20718;
wire n_20719;
wire n_2072;
wire n_20720;
wire n_20721;
wire n_20722;
wire n_20723;
wire n_20724;
wire n_20725;
wire n_20726;
wire n_20727;
wire n_20728;
wire n_20729;
wire n_2073;
wire n_20730;
wire n_20731;
wire n_20732;
wire n_20733;
wire n_20734;
wire n_20735;
wire n_20736;
wire n_20737;
wire n_20738;
wire n_20739;
wire n_2074;
wire n_20740;
wire n_20741;
wire n_20742;
wire n_20743;
wire n_20744;
wire n_20745;
wire n_20746;
wire n_20747;
wire n_20748;
wire n_20749;
wire n_2075;
wire n_20750;
wire n_20751;
wire n_20752;
wire n_20753;
wire n_20754;
wire n_20755;
wire n_20756;
wire n_20757;
wire n_20758;
wire n_20759;
wire n_2076;
wire n_20760;
wire n_20761;
wire n_20762;
wire n_20763;
wire n_20764;
wire n_20765;
wire n_20766;
wire n_20767;
wire n_20768;
wire n_20769;
wire n_2077;
wire n_20770;
wire n_20771;
wire n_20772;
wire n_20773;
wire n_20774;
wire n_20775;
wire n_20776;
wire n_20777;
wire n_20778;
wire n_20779;
wire n_2078;
wire n_20780;
wire n_20781;
wire n_20782;
wire n_20783;
wire n_20784;
wire n_20785;
wire n_20786;
wire n_20787;
wire n_20788;
wire n_20789;
wire n_2079;
wire n_20790;
wire n_20791;
wire n_20792;
wire n_20793;
wire n_20794;
wire n_20795;
wire n_20796;
wire n_20797;
wire n_20798;
wire n_20799;
wire n_208;
wire n_2080;
wire n_20800;
wire n_20801;
wire n_20802;
wire n_20803;
wire n_20804;
wire n_20805;
wire n_20806;
wire n_20807;
wire n_20808;
wire n_20809;
wire n_2081;
wire n_20810;
wire n_20811;
wire n_20812;
wire n_20813;
wire n_20814;
wire n_20815;
wire n_20816;
wire n_20817;
wire n_20818;
wire n_20819;
wire n_2082;
wire n_20820;
wire n_20821;
wire n_20822;
wire n_20823;
wire n_20824;
wire n_20825;
wire n_20826;
wire n_20827;
wire n_20828;
wire n_20829;
wire n_20830;
wire n_20831;
wire n_20832;
wire n_20833;
wire n_20834;
wire n_20835;
wire n_20836;
wire n_20837;
wire n_20838;
wire n_20839;
wire n_2084;
wire n_20840;
wire n_20841;
wire n_20842;
wire n_20843;
wire n_20844;
wire n_20845;
wire n_20846;
wire n_20847;
wire n_20848;
wire n_20849;
wire n_2085;
wire n_20850;
wire n_20851;
wire n_20852;
wire n_20853;
wire n_20854;
wire n_20855;
wire n_20856;
wire n_20857;
wire n_20858;
wire n_20859;
wire n_2086;
wire n_20860;
wire n_20861;
wire n_20862;
wire n_20863;
wire n_20864;
wire n_20865;
wire n_20866;
wire n_20867;
wire n_20868;
wire n_20869;
wire n_2087;
wire n_20870;
wire n_20871;
wire n_20872;
wire n_20873;
wire n_20874;
wire n_20875;
wire n_20876;
wire n_20877;
wire n_20878;
wire n_20879;
wire n_2088;
wire n_20880;
wire n_20881;
wire n_20882;
wire n_20883;
wire n_20885;
wire n_20886;
wire n_20887;
wire n_20888;
wire n_20889;
wire n_2089;
wire n_20890;
wire n_20891;
wire n_20892;
wire n_20893;
wire n_20894;
wire n_20895;
wire n_20896;
wire n_20897;
wire n_20898;
wire n_20899;
wire n_209;
wire n_2090;
wire n_20900;
wire n_20901;
wire n_20902;
wire n_20903;
wire n_20904;
wire n_20905;
wire n_20906;
wire n_20907;
wire n_20908;
wire n_20909;
wire n_2091;
wire n_20910;
wire n_20911;
wire n_20912;
wire n_20913;
wire n_20914;
wire n_20915;
wire n_20916;
wire n_20917;
wire n_20918;
wire n_20919;
wire n_2092;
wire n_20920;
wire n_20921;
wire n_20922;
wire n_20923;
wire n_20924;
wire n_20925;
wire n_20926;
wire n_20927;
wire n_20928;
wire n_20929;
wire n_2093;
wire n_20930;
wire n_20931;
wire n_20932;
wire n_20933;
wire n_20934;
wire n_20935;
wire n_20936;
wire n_20937;
wire n_20938;
wire n_20939;
wire n_2094;
wire n_20940;
wire n_20941;
wire n_20942;
wire n_20943;
wire n_20944;
wire n_20945;
wire n_20946;
wire n_20947;
wire n_20948;
wire n_20949;
wire n_2095;
wire n_20950;
wire n_20951;
wire n_20952;
wire n_20953;
wire n_20954;
wire n_20955;
wire n_20956;
wire n_20957;
wire n_20958;
wire n_20959;
wire n_2096;
wire n_20960;
wire n_20961;
wire n_20962;
wire n_20963;
wire n_20964;
wire n_20965;
wire n_20966;
wire n_20967;
wire n_20968;
wire n_20969;
wire n_2097;
wire n_20970;
wire n_20971;
wire n_20972;
wire n_20973;
wire n_20974;
wire n_20975;
wire n_20976;
wire n_20977;
wire n_20978;
wire n_20979;
wire n_2098;
wire n_20980;
wire n_20981;
wire n_20982;
wire n_20983;
wire n_20984;
wire n_20985;
wire n_20986;
wire n_20987;
wire n_20988;
wire n_20989;
wire n_2099;
wire n_20990;
wire n_20991;
wire n_20992;
wire n_20993;
wire n_20994;
wire n_20995;
wire n_20996;
wire n_20997;
wire n_20998;
wire n_20999;
wire n_21;
wire n_210;
wire n_2100;
wire n_21000;
wire n_21001;
wire n_21002;
wire n_21003;
wire n_21004;
wire n_21005;
wire n_21006;
wire n_21007;
wire n_21008;
wire n_21009;
wire n_2101;
wire n_21010;
wire n_21011;
wire n_21012;
wire n_21013;
wire n_21014;
wire n_21015;
wire n_21016;
wire n_21017;
wire n_21018;
wire n_21019;
wire n_2102;
wire n_21020;
wire n_21021;
wire n_21022;
wire n_21023;
wire n_21024;
wire n_21025;
wire n_21026;
wire n_21027;
wire n_21028;
wire n_21029;
wire n_2103;
wire n_21030;
wire n_21031;
wire n_21032;
wire n_21033;
wire n_21034;
wire n_21035;
wire n_21036;
wire n_21037;
wire n_21038;
wire n_21039;
wire n_2104;
wire n_21040;
wire n_21041;
wire n_21042;
wire n_21043;
wire n_21044;
wire n_21045;
wire n_21046;
wire n_21047;
wire n_21048;
wire n_21049;
wire n_2105;
wire n_21050;
wire n_21051;
wire n_21052;
wire n_21053;
wire n_21054;
wire n_21055;
wire n_21056;
wire n_21057;
wire n_21058;
wire n_21059;
wire n_2106;
wire n_21060;
wire n_21061;
wire n_21062;
wire n_21063;
wire n_21064;
wire n_21065;
wire n_21066;
wire n_21067;
wire n_21068;
wire n_21069;
wire n_2107;
wire n_21070;
wire n_21071;
wire n_21072;
wire n_21073;
wire n_21074;
wire n_21075;
wire n_21076;
wire n_21077;
wire n_21078;
wire n_21079;
wire n_2108;
wire n_21080;
wire n_21081;
wire n_21082;
wire n_21083;
wire n_21084;
wire n_21085;
wire n_21086;
wire n_21087;
wire n_21088;
wire n_21089;
wire n_2109;
wire n_21090;
wire n_21091;
wire n_21092;
wire n_21093;
wire n_21094;
wire n_21095;
wire n_21096;
wire n_21097;
wire n_21098;
wire n_21099;
wire n_211;
wire n_2110;
wire n_21100;
wire n_21102;
wire n_21103;
wire n_21104;
wire n_21105;
wire n_21106;
wire n_21107;
wire n_21108;
wire n_21109;
wire n_2111;
wire n_21110;
wire n_21111;
wire n_21112;
wire n_21113;
wire n_21114;
wire n_21115;
wire n_21116;
wire n_21117;
wire n_21118;
wire n_21119;
wire n_2112;
wire n_21120;
wire n_21121;
wire n_21122;
wire n_21123;
wire n_21124;
wire n_21125;
wire n_21126;
wire n_21127;
wire n_21128;
wire n_21129;
wire n_2113;
wire n_21130;
wire n_21131;
wire n_21132;
wire n_21133;
wire n_21134;
wire n_21135;
wire n_21136;
wire n_21137;
wire n_21138;
wire n_21139;
wire n_2114;
wire n_21140;
wire n_21141;
wire n_21142;
wire n_21143;
wire n_21144;
wire n_21145;
wire n_21146;
wire n_21147;
wire n_21148;
wire n_21149;
wire n_2115;
wire n_21150;
wire n_21151;
wire n_21152;
wire n_21153;
wire n_21154;
wire n_21155;
wire n_21156;
wire n_21157;
wire n_21158;
wire n_21159;
wire n_2116;
wire n_21160;
wire n_21161;
wire n_21162;
wire n_21163;
wire n_21164;
wire n_21165;
wire n_21166;
wire n_21167;
wire n_21168;
wire n_21169;
wire n_21170;
wire n_21171;
wire n_21172;
wire n_21173;
wire n_21174;
wire n_21175;
wire n_21176;
wire n_21177;
wire n_21178;
wire n_21179;
wire n_2118;
wire n_21180;
wire n_21181;
wire n_21182;
wire n_21183;
wire n_21184;
wire n_21185;
wire n_21186;
wire n_21187;
wire n_21188;
wire n_21189;
wire n_2119;
wire n_21190;
wire n_21191;
wire n_21192;
wire n_21193;
wire n_21194;
wire n_21195;
wire n_21196;
wire n_21197;
wire n_21198;
wire n_21199;
wire n_212;
wire n_2120;
wire n_21200;
wire n_21201;
wire n_21202;
wire n_21203;
wire n_21204;
wire n_21205;
wire n_21206;
wire n_21207;
wire n_21208;
wire n_21209;
wire n_2121;
wire n_21210;
wire n_21211;
wire n_21212;
wire n_21213;
wire n_21214;
wire n_21215;
wire n_21216;
wire n_21217;
wire n_21218;
wire n_21219;
wire n_2122;
wire n_21220;
wire n_21221;
wire n_21222;
wire n_21223;
wire n_21224;
wire n_21225;
wire n_21226;
wire n_21227;
wire n_21228;
wire n_21229;
wire n_2123;
wire n_21230;
wire n_21231;
wire n_21232;
wire n_21233;
wire n_21234;
wire n_21235;
wire n_21236;
wire n_21237;
wire n_21238;
wire n_21239;
wire n_2124;
wire n_21240;
wire n_21241;
wire n_21242;
wire n_21243;
wire n_21244;
wire n_21245;
wire n_21246;
wire n_21247;
wire n_21248;
wire n_21249;
wire n_2125;
wire n_21250;
wire n_21251;
wire n_21252;
wire n_21253;
wire n_21254;
wire n_21255;
wire n_21256;
wire n_21257;
wire n_21258;
wire n_21259;
wire n_2126;
wire n_21260;
wire n_21261;
wire n_21262;
wire n_21263;
wire n_21264;
wire n_21265;
wire n_21266;
wire n_21267;
wire n_21268;
wire n_21269;
wire n_2127;
wire n_21270;
wire n_21271;
wire n_21272;
wire n_21273;
wire n_21274;
wire n_21275;
wire n_21276;
wire n_21277;
wire n_21278;
wire n_21279;
wire n_2128;
wire n_21280;
wire n_21281;
wire n_21282;
wire n_21283;
wire n_21284;
wire n_21285;
wire n_21286;
wire n_21287;
wire n_21288;
wire n_21289;
wire n_2129;
wire n_21290;
wire n_21291;
wire n_21292;
wire n_21293;
wire n_21294;
wire n_21295;
wire n_21296;
wire n_21297;
wire n_21298;
wire n_21299;
wire n_213;
wire n_2130;
wire n_21300;
wire n_21301;
wire n_21302;
wire n_21303;
wire n_21304;
wire n_21305;
wire n_21306;
wire n_21307;
wire n_21308;
wire n_21309;
wire n_2131;
wire n_21310;
wire n_21311;
wire n_21312;
wire n_21313;
wire n_21314;
wire n_21315;
wire n_21316;
wire n_21317;
wire n_21318;
wire n_21319;
wire n_2132;
wire n_21320;
wire n_21321;
wire n_21322;
wire n_21323;
wire n_21324;
wire n_21325;
wire n_21326;
wire n_21327;
wire n_21328;
wire n_21329;
wire n_2133;
wire n_21330;
wire n_21331;
wire n_21332;
wire n_21333;
wire n_21334;
wire n_21335;
wire n_21336;
wire n_21337;
wire n_21338;
wire n_21339;
wire n_2134;
wire n_21340;
wire n_21341;
wire n_21342;
wire n_21343;
wire n_21344;
wire n_21345;
wire n_21346;
wire n_21347;
wire n_21348;
wire n_21349;
wire n_2135;
wire n_21350;
wire n_21351;
wire n_21352;
wire n_21353;
wire n_21354;
wire n_21355;
wire n_21356;
wire n_21357;
wire n_21358;
wire n_21359;
wire n_2136;
wire n_21360;
wire n_21361;
wire n_21362;
wire n_21363;
wire n_21364;
wire n_21365;
wire n_21366;
wire n_21367;
wire n_21368;
wire n_21369;
wire n_2137;
wire n_21370;
wire n_21371;
wire n_21372;
wire n_21373;
wire n_21374;
wire n_21375;
wire n_21376;
wire n_21377;
wire n_21378;
wire n_21379;
wire n_2138;
wire n_21380;
wire n_21381;
wire n_21382;
wire n_21383;
wire n_21384;
wire n_21385;
wire n_21386;
wire n_21387;
wire n_21388;
wire n_21389;
wire n_2139;
wire n_21390;
wire n_21391;
wire n_21392;
wire n_21393;
wire n_21394;
wire n_21395;
wire n_21396;
wire n_21397;
wire n_21398;
wire n_21399;
wire n_214;
wire n_2140;
wire n_21400;
wire n_21401;
wire n_21402;
wire n_21403;
wire n_21404;
wire n_21405;
wire n_21406;
wire n_21407;
wire n_21408;
wire n_21409;
wire n_2141;
wire n_21410;
wire n_21411;
wire n_21412;
wire n_21413;
wire n_21414;
wire n_21415;
wire n_21416;
wire n_21417;
wire n_21418;
wire n_21419;
wire n_2142;
wire n_21420;
wire n_21421;
wire n_21422;
wire n_21423;
wire n_21424;
wire n_21425;
wire n_21426;
wire n_21427;
wire n_21428;
wire n_21429;
wire n_2143;
wire n_21430;
wire n_21431;
wire n_21432;
wire n_21433;
wire n_21434;
wire n_21435;
wire n_21436;
wire n_21437;
wire n_21438;
wire n_21439;
wire n_2144;
wire n_21440;
wire n_21441;
wire n_21442;
wire n_21443;
wire n_21444;
wire n_21445;
wire n_21446;
wire n_21447;
wire n_21448;
wire n_21449;
wire n_2145;
wire n_21450;
wire n_21451;
wire n_21452;
wire n_21453;
wire n_21454;
wire n_21455;
wire n_21456;
wire n_21457;
wire n_21458;
wire n_21459;
wire n_2146;
wire n_21460;
wire n_21461;
wire n_21462;
wire n_21463;
wire n_21464;
wire n_21465;
wire n_21466;
wire n_21467;
wire n_21468;
wire n_21469;
wire n_2147;
wire n_21470;
wire n_21471;
wire n_21472;
wire n_21473;
wire n_21474;
wire n_21475;
wire n_21476;
wire n_21477;
wire n_21478;
wire n_21479;
wire n_2148;
wire n_21480;
wire n_21481;
wire n_21482;
wire n_21483;
wire n_21484;
wire n_21485;
wire n_21486;
wire n_21487;
wire n_21488;
wire n_21489;
wire n_2149;
wire n_21490;
wire n_21491;
wire n_21492;
wire n_21493;
wire n_21494;
wire n_21495;
wire n_21496;
wire n_21497;
wire n_21498;
wire n_21499;
wire n_215;
wire n_2150;
wire n_21500;
wire n_21501;
wire n_21502;
wire n_21503;
wire n_21504;
wire n_21505;
wire n_21506;
wire n_21507;
wire n_21508;
wire n_21509;
wire n_2151;
wire n_21510;
wire n_21511;
wire n_21512;
wire n_21513;
wire n_21514;
wire n_21515;
wire n_21516;
wire n_21517;
wire n_21518;
wire n_21519;
wire n_2152;
wire n_21520;
wire n_21521;
wire n_21522;
wire n_21523;
wire n_21524;
wire n_21525;
wire n_21526;
wire n_21527;
wire n_21528;
wire n_21529;
wire n_2153;
wire n_21530;
wire n_21531;
wire n_21532;
wire n_21533;
wire n_21534;
wire n_21535;
wire n_21536;
wire n_21537;
wire n_21538;
wire n_21539;
wire n_2154;
wire n_21540;
wire n_21541;
wire n_21542;
wire n_21543;
wire n_21544;
wire n_21545;
wire n_21546;
wire n_21547;
wire n_21548;
wire n_21549;
wire n_2155;
wire n_21550;
wire n_21551;
wire n_21552;
wire n_21553;
wire n_21554;
wire n_21555;
wire n_21556;
wire n_21557;
wire n_21558;
wire n_21559;
wire n_2156;
wire n_21560;
wire n_21561;
wire n_21562;
wire n_21563;
wire n_21564;
wire n_21565;
wire n_21566;
wire n_21567;
wire n_21568;
wire n_21569;
wire n_2157;
wire n_21570;
wire n_21571;
wire n_21572;
wire n_21573;
wire n_21574;
wire n_21575;
wire n_21576;
wire n_21577;
wire n_21578;
wire n_21579;
wire n_2158;
wire n_21580;
wire n_21581;
wire n_21582;
wire n_21583;
wire n_21584;
wire n_21585;
wire n_21586;
wire n_21587;
wire n_21588;
wire n_21589;
wire n_2159;
wire n_21590;
wire n_21591;
wire n_21592;
wire n_21593;
wire n_21594;
wire n_21595;
wire n_21596;
wire n_21597;
wire n_21598;
wire n_21599;
wire n_216;
wire n_2160;
wire n_21600;
wire n_21601;
wire n_21602;
wire n_21603;
wire n_21604;
wire n_21605;
wire n_21606;
wire n_21607;
wire n_21609;
wire n_2161;
wire n_21610;
wire n_21611;
wire n_21612;
wire n_21613;
wire n_21614;
wire n_21615;
wire n_21616;
wire n_21617;
wire n_21618;
wire n_21619;
wire n_2162;
wire n_21620;
wire n_21621;
wire n_21622;
wire n_21623;
wire n_21624;
wire n_21625;
wire n_21626;
wire n_21627;
wire n_21628;
wire n_21629;
wire n_2163;
wire n_21630;
wire n_21631;
wire n_21632;
wire n_21633;
wire n_21634;
wire n_21635;
wire n_21636;
wire n_21637;
wire n_21639;
wire n_2164;
wire n_21640;
wire n_21641;
wire n_21643;
wire n_21644;
wire n_21645;
wire n_21646;
wire n_21647;
wire n_21648;
wire n_21649;
wire n_2165;
wire n_21650;
wire n_21651;
wire n_21652;
wire n_21653;
wire n_21654;
wire n_21655;
wire n_21656;
wire n_21657;
wire n_21658;
wire n_21659;
wire n_2166;
wire n_21660;
wire n_21661;
wire n_21662;
wire n_21663;
wire n_21664;
wire n_21665;
wire n_21666;
wire n_21667;
wire n_21668;
wire n_21669;
wire n_2167;
wire n_21670;
wire n_21671;
wire n_21672;
wire n_21673;
wire n_21674;
wire n_21675;
wire n_21676;
wire n_21677;
wire n_21678;
wire n_21679;
wire n_2168;
wire n_21680;
wire n_21681;
wire n_21682;
wire n_21683;
wire n_21684;
wire n_21685;
wire n_21686;
wire n_21687;
wire n_21688;
wire n_21689;
wire n_2169;
wire n_21690;
wire n_21691;
wire n_21692;
wire n_21693;
wire n_21694;
wire n_21695;
wire n_21696;
wire n_21697;
wire n_21698;
wire n_21699;
wire n_217;
wire n_2170;
wire n_21700;
wire n_21701;
wire n_21702;
wire n_21703;
wire n_21704;
wire n_21705;
wire n_21706;
wire n_21707;
wire n_21708;
wire n_21709;
wire n_2171;
wire n_21710;
wire n_21711;
wire n_21712;
wire n_21713;
wire n_21714;
wire n_21715;
wire n_21716;
wire n_21717;
wire n_21718;
wire n_21719;
wire n_2172;
wire n_21720;
wire n_21721;
wire n_21722;
wire n_21723;
wire n_21724;
wire n_21725;
wire n_21726;
wire n_21727;
wire n_21728;
wire n_21729;
wire n_2173;
wire n_21730;
wire n_21731;
wire n_21732;
wire n_21733;
wire n_21734;
wire n_21735;
wire n_21736;
wire n_21737;
wire n_21738;
wire n_21739;
wire n_2174;
wire n_21740;
wire n_21741;
wire n_21742;
wire n_21743;
wire n_21744;
wire n_21745;
wire n_21746;
wire n_21747;
wire n_21748;
wire n_21749;
wire n_2175;
wire n_21750;
wire n_21751;
wire n_21752;
wire n_21753;
wire n_21754;
wire n_21755;
wire n_21756;
wire n_21757;
wire n_21758;
wire n_21759;
wire n_2176;
wire n_21760;
wire n_21761;
wire n_21762;
wire n_21763;
wire n_21764;
wire n_21765;
wire n_21766;
wire n_21767;
wire n_21768;
wire n_21769;
wire n_2177;
wire n_21770;
wire n_21771;
wire n_21772;
wire n_21773;
wire n_21774;
wire n_21775;
wire n_21776;
wire n_21777;
wire n_21778;
wire n_21779;
wire n_2178;
wire n_21780;
wire n_21781;
wire n_21782;
wire n_21783;
wire n_21784;
wire n_21785;
wire n_21786;
wire n_21787;
wire n_21788;
wire n_21789;
wire n_2179;
wire n_21790;
wire n_21791;
wire n_21792;
wire n_21793;
wire n_21794;
wire n_21795;
wire n_21796;
wire n_21797;
wire n_21798;
wire n_21799;
wire n_218;
wire n_2180;
wire n_21800;
wire n_21801;
wire n_21802;
wire n_21803;
wire n_21804;
wire n_21805;
wire n_21806;
wire n_21807;
wire n_21808;
wire n_21809;
wire n_2181;
wire n_21810;
wire n_21811;
wire n_21812;
wire n_21813;
wire n_21814;
wire n_21815;
wire n_21816;
wire n_21817;
wire n_21818;
wire n_21819;
wire n_2182;
wire n_21820;
wire n_21821;
wire n_21822;
wire n_21823;
wire n_21824;
wire n_21825;
wire n_21826;
wire n_21827;
wire n_21828;
wire n_21829;
wire n_2183;
wire n_21830;
wire n_21831;
wire n_21832;
wire n_21833;
wire n_21834;
wire n_21835;
wire n_21836;
wire n_21837;
wire n_21838;
wire n_21839;
wire n_2184;
wire n_21840;
wire n_21841;
wire n_21842;
wire n_21843;
wire n_21844;
wire n_21845;
wire n_21846;
wire n_21847;
wire n_21848;
wire n_21849;
wire n_2185;
wire n_21850;
wire n_21851;
wire n_21852;
wire n_21853;
wire n_21854;
wire n_21855;
wire n_21856;
wire n_21857;
wire n_21858;
wire n_21859;
wire n_2186;
wire n_21860;
wire n_21861;
wire n_21862;
wire n_21863;
wire n_21864;
wire n_21865;
wire n_21866;
wire n_21867;
wire n_21868;
wire n_21869;
wire n_2187;
wire n_21870;
wire n_21871;
wire n_21872;
wire n_21873;
wire n_21874;
wire n_21875;
wire n_21876;
wire n_21877;
wire n_21878;
wire n_21879;
wire n_2188;
wire n_21880;
wire n_21881;
wire n_21882;
wire n_21883;
wire n_21884;
wire n_21885;
wire n_21886;
wire n_21887;
wire n_21888;
wire n_21889;
wire n_2189;
wire n_21890;
wire n_21891;
wire n_21892;
wire n_21893;
wire n_21894;
wire n_21895;
wire n_21896;
wire n_21897;
wire n_21898;
wire n_21899;
wire n_219;
wire n_2190;
wire n_21900;
wire n_21901;
wire n_21902;
wire n_21903;
wire n_21904;
wire n_21905;
wire n_21906;
wire n_21907;
wire n_21908;
wire n_21909;
wire n_2191;
wire n_21910;
wire n_21911;
wire n_21912;
wire n_21913;
wire n_21914;
wire n_21915;
wire n_21916;
wire n_21917;
wire n_21918;
wire n_21919;
wire n_2192;
wire n_21920;
wire n_21921;
wire n_21922;
wire n_21923;
wire n_21924;
wire n_21925;
wire n_21926;
wire n_21927;
wire n_21928;
wire n_21929;
wire n_2193;
wire n_21930;
wire n_21931;
wire n_21932;
wire n_21933;
wire n_21934;
wire n_21935;
wire n_21936;
wire n_21937;
wire n_21938;
wire n_21939;
wire n_2194;
wire n_21940;
wire n_21941;
wire n_21942;
wire n_21943;
wire n_21944;
wire n_21945;
wire n_21946;
wire n_21947;
wire n_21948;
wire n_21949;
wire n_2195;
wire n_21950;
wire n_21951;
wire n_21952;
wire n_21953;
wire n_21954;
wire n_21955;
wire n_21956;
wire n_21957;
wire n_21958;
wire n_21959;
wire n_2196;
wire n_21960;
wire n_21961;
wire n_21962;
wire n_21963;
wire n_21964;
wire n_21965;
wire n_21966;
wire n_21967;
wire n_21968;
wire n_21969;
wire n_2197;
wire n_21970;
wire n_21971;
wire n_21972;
wire n_21973;
wire n_21974;
wire n_21975;
wire n_21976;
wire n_21977;
wire n_21978;
wire n_21979;
wire n_2198;
wire n_21980;
wire n_21981;
wire n_21982;
wire n_21983;
wire n_21984;
wire n_21985;
wire n_21986;
wire n_21987;
wire n_21988;
wire n_21989;
wire n_2199;
wire n_21990;
wire n_21991;
wire n_21992;
wire n_21993;
wire n_21994;
wire n_21995;
wire n_21996;
wire n_21997;
wire n_21998;
wire n_21999;
wire n_22;
wire n_220;
wire n_22000;
wire n_22001;
wire n_22002;
wire n_22003;
wire n_22004;
wire n_22005;
wire n_22006;
wire n_22007;
wire n_22008;
wire n_22009;
wire n_22010;
wire n_22011;
wire n_22012;
wire n_22013;
wire n_22014;
wire n_22015;
wire n_22016;
wire n_22017;
wire n_22018;
wire n_22019;
wire n_2202;
wire n_22020;
wire n_22021;
wire n_22022;
wire n_22023;
wire n_22024;
wire n_22025;
wire n_22026;
wire n_22027;
wire n_22028;
wire n_22029;
wire n_2203;
wire n_22030;
wire n_22031;
wire n_22032;
wire n_22033;
wire n_22034;
wire n_22035;
wire n_22036;
wire n_22037;
wire n_22038;
wire n_22039;
wire n_2204;
wire n_22040;
wire n_22041;
wire n_22042;
wire n_22043;
wire n_22044;
wire n_22045;
wire n_22046;
wire n_22047;
wire n_22048;
wire n_2205;
wire n_22050;
wire n_22051;
wire n_22052;
wire n_22053;
wire n_22054;
wire n_22055;
wire n_22056;
wire n_22057;
wire n_22058;
wire n_22059;
wire n_2206;
wire n_22060;
wire n_22061;
wire n_22062;
wire n_22063;
wire n_22064;
wire n_22065;
wire n_22066;
wire n_22067;
wire n_22068;
wire n_22069;
wire n_2207;
wire n_22070;
wire n_22072;
wire n_22073;
wire n_22074;
wire n_22075;
wire n_22076;
wire n_22077;
wire n_22078;
wire n_22079;
wire n_2208;
wire n_22080;
wire n_22081;
wire n_22082;
wire n_22083;
wire n_22084;
wire n_22085;
wire n_22086;
wire n_22087;
wire n_22088;
wire n_22089;
wire n_2209;
wire n_22090;
wire n_22091;
wire n_22092;
wire n_22093;
wire n_22094;
wire n_22095;
wire n_22096;
wire n_22097;
wire n_22098;
wire n_22099;
wire n_221;
wire n_2210;
wire n_22100;
wire n_22101;
wire n_22102;
wire n_22103;
wire n_22104;
wire n_22105;
wire n_22106;
wire n_22107;
wire n_22108;
wire n_22109;
wire n_2211;
wire n_22110;
wire n_22112;
wire n_22113;
wire n_22114;
wire n_22115;
wire n_22116;
wire n_22117;
wire n_22118;
wire n_22119;
wire n_2212;
wire n_22120;
wire n_22121;
wire n_22122;
wire n_22123;
wire n_22124;
wire n_22125;
wire n_22126;
wire n_22127;
wire n_22128;
wire n_22129;
wire n_2213;
wire n_22130;
wire n_22131;
wire n_22132;
wire n_22133;
wire n_22134;
wire n_22135;
wire n_22136;
wire n_22137;
wire n_22138;
wire n_22139;
wire n_2214;
wire n_22140;
wire n_22141;
wire n_22142;
wire n_22143;
wire n_22144;
wire n_22145;
wire n_22146;
wire n_22147;
wire n_22148;
wire n_22149;
wire n_2215;
wire n_22150;
wire n_22151;
wire n_22152;
wire n_22153;
wire n_22154;
wire n_22155;
wire n_22156;
wire n_22157;
wire n_22158;
wire n_22159;
wire n_2216;
wire n_22160;
wire n_22161;
wire n_22162;
wire n_22163;
wire n_22164;
wire n_22165;
wire n_22166;
wire n_22167;
wire n_22168;
wire n_22169;
wire n_2217;
wire n_22170;
wire n_22171;
wire n_22172;
wire n_22173;
wire n_22174;
wire n_22175;
wire n_22176;
wire n_22177;
wire n_22178;
wire n_22179;
wire n_2218;
wire n_22180;
wire n_22181;
wire n_22182;
wire n_22183;
wire n_22184;
wire n_22185;
wire n_22186;
wire n_22187;
wire n_22188;
wire n_22189;
wire n_2219;
wire n_22190;
wire n_22191;
wire n_22192;
wire n_22193;
wire n_22194;
wire n_22195;
wire n_22196;
wire n_22197;
wire n_22198;
wire n_22199;
wire n_222;
wire n_2220;
wire n_22200;
wire n_22201;
wire n_22202;
wire n_22203;
wire n_22204;
wire n_22205;
wire n_22206;
wire n_22207;
wire n_22208;
wire n_22209;
wire n_2221;
wire n_22210;
wire n_22211;
wire n_22212;
wire n_22213;
wire n_22214;
wire n_22215;
wire n_22216;
wire n_22217;
wire n_22218;
wire n_22219;
wire n_2222;
wire n_22220;
wire n_22221;
wire n_22222;
wire n_22223;
wire n_22224;
wire n_22225;
wire n_22226;
wire n_22227;
wire n_22228;
wire n_22229;
wire n_2223;
wire n_22230;
wire n_22231;
wire n_22232;
wire n_22233;
wire n_22234;
wire n_22235;
wire n_22236;
wire n_22237;
wire n_22238;
wire n_22239;
wire n_2224;
wire n_22240;
wire n_22241;
wire n_22242;
wire n_22243;
wire n_22244;
wire n_22245;
wire n_22246;
wire n_22247;
wire n_22248;
wire n_22249;
wire n_2225;
wire n_22250;
wire n_22251;
wire n_22252;
wire n_22253;
wire n_22254;
wire n_22255;
wire n_22256;
wire n_22257;
wire n_22258;
wire n_22259;
wire n_2226;
wire n_22260;
wire n_22261;
wire n_22262;
wire n_22263;
wire n_22264;
wire n_22265;
wire n_22266;
wire n_22267;
wire n_22268;
wire n_22269;
wire n_2227;
wire n_22270;
wire n_22271;
wire n_22272;
wire n_22273;
wire n_22274;
wire n_22275;
wire n_22276;
wire n_22278;
wire n_22279;
wire n_2228;
wire n_22280;
wire n_22281;
wire n_22282;
wire n_22283;
wire n_22284;
wire n_22285;
wire n_22286;
wire n_22287;
wire n_22288;
wire n_22289;
wire n_22290;
wire n_22291;
wire n_22292;
wire n_22293;
wire n_22294;
wire n_22295;
wire n_22296;
wire n_22297;
wire n_22298;
wire n_22299;
wire n_223;
wire n_2230;
wire n_22300;
wire n_22301;
wire n_22302;
wire n_22303;
wire n_22304;
wire n_22305;
wire n_22306;
wire n_22307;
wire n_22308;
wire n_22309;
wire n_2231;
wire n_22311;
wire n_22312;
wire n_22313;
wire n_22314;
wire n_22315;
wire n_22316;
wire n_22317;
wire n_22318;
wire n_22319;
wire n_2232;
wire n_22320;
wire n_22321;
wire n_22322;
wire n_22323;
wire n_22324;
wire n_22325;
wire n_22326;
wire n_22327;
wire n_22328;
wire n_22329;
wire n_2233;
wire n_22330;
wire n_22331;
wire n_22332;
wire n_22333;
wire n_22334;
wire n_22335;
wire n_22336;
wire n_22337;
wire n_22338;
wire n_22339;
wire n_2234;
wire n_22340;
wire n_22341;
wire n_22342;
wire n_22343;
wire n_22344;
wire n_22345;
wire n_22346;
wire n_22347;
wire n_22348;
wire n_22349;
wire n_2235;
wire n_22350;
wire n_22351;
wire n_22352;
wire n_22353;
wire n_22354;
wire n_22355;
wire n_22356;
wire n_22357;
wire n_22358;
wire n_22359;
wire n_2236;
wire n_22360;
wire n_22361;
wire n_22362;
wire n_22363;
wire n_22364;
wire n_22365;
wire n_22366;
wire n_22367;
wire n_22368;
wire n_22369;
wire n_2237;
wire n_22371;
wire n_22373;
wire n_22374;
wire n_22375;
wire n_22376;
wire n_22377;
wire n_22378;
wire n_22379;
wire n_2238;
wire n_22380;
wire n_22381;
wire n_22382;
wire n_22383;
wire n_22384;
wire n_22385;
wire n_22386;
wire n_22387;
wire n_22388;
wire n_22389;
wire n_2239;
wire n_22390;
wire n_22391;
wire n_22392;
wire n_22393;
wire n_22394;
wire n_22395;
wire n_22396;
wire n_22397;
wire n_22398;
wire n_22399;
wire n_224;
wire n_2240;
wire n_22400;
wire n_22401;
wire n_22402;
wire n_22403;
wire n_22404;
wire n_22405;
wire n_22406;
wire n_22407;
wire n_22408;
wire n_22409;
wire n_2241;
wire n_22410;
wire n_22411;
wire n_22412;
wire n_22413;
wire n_22414;
wire n_22415;
wire n_22416;
wire n_22417;
wire n_22418;
wire n_22419;
wire n_2242;
wire n_22420;
wire n_22421;
wire n_22422;
wire n_22423;
wire n_22424;
wire n_22425;
wire n_22426;
wire n_22427;
wire n_22428;
wire n_22429;
wire n_2243;
wire n_22430;
wire n_22431;
wire n_22432;
wire n_22433;
wire n_22434;
wire n_22435;
wire n_22436;
wire n_22437;
wire n_22438;
wire n_22439;
wire n_2244;
wire n_22440;
wire n_22441;
wire n_22442;
wire n_22443;
wire n_22444;
wire n_22445;
wire n_22446;
wire n_22447;
wire n_22448;
wire n_22449;
wire n_2245;
wire n_22450;
wire n_22451;
wire n_22452;
wire n_22453;
wire n_22454;
wire n_22455;
wire n_22456;
wire n_22457;
wire n_22458;
wire n_22459;
wire n_2246;
wire n_22460;
wire n_22461;
wire n_22462;
wire n_22463;
wire n_22464;
wire n_22465;
wire n_22466;
wire n_22467;
wire n_22468;
wire n_22469;
wire n_2247;
wire n_22470;
wire n_22471;
wire n_22472;
wire n_22473;
wire n_22474;
wire n_22475;
wire n_22476;
wire n_22477;
wire n_22478;
wire n_22479;
wire n_2248;
wire n_22480;
wire n_22481;
wire n_22482;
wire n_22483;
wire n_22484;
wire n_22485;
wire n_22486;
wire n_22487;
wire n_22488;
wire n_22489;
wire n_2249;
wire n_22490;
wire n_22491;
wire n_22492;
wire n_22493;
wire n_22494;
wire n_22495;
wire n_22496;
wire n_22497;
wire n_22498;
wire n_22499;
wire n_225;
wire n_2250;
wire n_22500;
wire n_22501;
wire n_22502;
wire n_22503;
wire n_22504;
wire n_22505;
wire n_22506;
wire n_22507;
wire n_22508;
wire n_22509;
wire n_2251;
wire n_22510;
wire n_22511;
wire n_22512;
wire n_22513;
wire n_22514;
wire n_22515;
wire n_22516;
wire n_22517;
wire n_22518;
wire n_22519;
wire n_2252;
wire n_22520;
wire n_22521;
wire n_22522;
wire n_22523;
wire n_22524;
wire n_22525;
wire n_22526;
wire n_22527;
wire n_22528;
wire n_22529;
wire n_2253;
wire n_22530;
wire n_22531;
wire n_22532;
wire n_22533;
wire n_22534;
wire n_22535;
wire n_22536;
wire n_22537;
wire n_22538;
wire n_22539;
wire n_2254;
wire n_22540;
wire n_22541;
wire n_22542;
wire n_22543;
wire n_22544;
wire n_22545;
wire n_22546;
wire n_22547;
wire n_22548;
wire n_22549;
wire n_2255;
wire n_22550;
wire n_22551;
wire n_22552;
wire n_22553;
wire n_22554;
wire n_22555;
wire n_22556;
wire n_22557;
wire n_22558;
wire n_22559;
wire n_2256;
wire n_22560;
wire n_22561;
wire n_22562;
wire n_22563;
wire n_22564;
wire n_22565;
wire n_22566;
wire n_22567;
wire n_22568;
wire n_22569;
wire n_2257;
wire n_22570;
wire n_22571;
wire n_22572;
wire n_22573;
wire n_22574;
wire n_22575;
wire n_22576;
wire n_22577;
wire n_22578;
wire n_22579;
wire n_2258;
wire n_22580;
wire n_22581;
wire n_22582;
wire n_22583;
wire n_22584;
wire n_22585;
wire n_22586;
wire n_22587;
wire n_22589;
wire n_2259;
wire n_22590;
wire n_22591;
wire n_22592;
wire n_22593;
wire n_22594;
wire n_22595;
wire n_22596;
wire n_22597;
wire n_22598;
wire n_22599;
wire n_226;
wire n_2260;
wire n_22600;
wire n_22601;
wire n_22602;
wire n_22603;
wire n_22604;
wire n_22605;
wire n_22606;
wire n_22607;
wire n_22609;
wire n_2261;
wire n_22610;
wire n_22611;
wire n_22612;
wire n_22613;
wire n_22614;
wire n_22615;
wire n_22616;
wire n_22617;
wire n_22618;
wire n_22619;
wire n_2262;
wire n_22620;
wire n_22621;
wire n_22622;
wire n_22623;
wire n_22624;
wire n_22625;
wire n_22626;
wire n_22627;
wire n_22628;
wire n_22629;
wire n_2263;
wire n_22630;
wire n_22631;
wire n_22632;
wire n_22633;
wire n_22634;
wire n_22635;
wire n_22636;
wire n_22637;
wire n_22638;
wire n_22639;
wire n_2264;
wire n_22640;
wire n_22641;
wire n_22642;
wire n_22643;
wire n_22644;
wire n_22645;
wire n_22646;
wire n_22647;
wire n_22648;
wire n_22649;
wire n_2265;
wire n_22650;
wire n_22651;
wire n_22652;
wire n_22653;
wire n_22654;
wire n_22655;
wire n_22656;
wire n_22657;
wire n_22658;
wire n_22659;
wire n_2266;
wire n_22660;
wire n_22661;
wire n_22662;
wire n_22663;
wire n_22664;
wire n_22665;
wire n_22666;
wire n_22667;
wire n_22668;
wire n_22669;
wire n_2267;
wire n_22670;
wire n_22671;
wire n_22672;
wire n_22673;
wire n_22674;
wire n_22675;
wire n_22676;
wire n_22677;
wire n_22678;
wire n_22679;
wire n_2268;
wire n_22680;
wire n_22681;
wire n_22682;
wire n_22683;
wire n_22684;
wire n_22685;
wire n_22686;
wire n_22687;
wire n_22688;
wire n_22689;
wire n_2269;
wire n_22690;
wire n_22691;
wire n_22692;
wire n_22693;
wire n_22694;
wire n_22695;
wire n_22696;
wire n_22697;
wire n_22698;
wire n_22699;
wire n_227;
wire n_2270;
wire n_22700;
wire n_22701;
wire n_22702;
wire n_22703;
wire n_22704;
wire n_22705;
wire n_22706;
wire n_22707;
wire n_22708;
wire n_22709;
wire n_2271;
wire n_22710;
wire n_22711;
wire n_22712;
wire n_22713;
wire n_22714;
wire n_22715;
wire n_22716;
wire n_22717;
wire n_22718;
wire n_22719;
wire n_2272;
wire n_22720;
wire n_22721;
wire n_22722;
wire n_22723;
wire n_22724;
wire n_22725;
wire n_22726;
wire n_22727;
wire n_22728;
wire n_22729;
wire n_2273;
wire n_22730;
wire n_22731;
wire n_22732;
wire n_22733;
wire n_22734;
wire n_22735;
wire n_22736;
wire n_22737;
wire n_22738;
wire n_22739;
wire n_2274;
wire n_22740;
wire n_22741;
wire n_22742;
wire n_22743;
wire n_22744;
wire n_22745;
wire n_22746;
wire n_22747;
wire n_22748;
wire n_22749;
wire n_2275;
wire n_22750;
wire n_22751;
wire n_22752;
wire n_22753;
wire n_22754;
wire n_22755;
wire n_22756;
wire n_22757;
wire n_22758;
wire n_22759;
wire n_2276;
wire n_22760;
wire n_22761;
wire n_22762;
wire n_22763;
wire n_22764;
wire n_22765;
wire n_22766;
wire n_22767;
wire n_22768;
wire n_22769;
wire n_2277;
wire n_22770;
wire n_22771;
wire n_22772;
wire n_22773;
wire n_22774;
wire n_22775;
wire n_22776;
wire n_22777;
wire n_22778;
wire n_22779;
wire n_2278;
wire n_22780;
wire n_22781;
wire n_22782;
wire n_22783;
wire n_22784;
wire n_22785;
wire n_22786;
wire n_22787;
wire n_22788;
wire n_22789;
wire n_2279;
wire n_22790;
wire n_22791;
wire n_22792;
wire n_22793;
wire n_22794;
wire n_22795;
wire n_22796;
wire n_22797;
wire n_22798;
wire n_22799;
wire n_228;
wire n_2280;
wire n_22800;
wire n_22801;
wire n_22802;
wire n_22803;
wire n_22804;
wire n_22805;
wire n_22806;
wire n_22807;
wire n_22808;
wire n_22809;
wire n_2281;
wire n_22810;
wire n_22811;
wire n_22812;
wire n_22813;
wire n_22814;
wire n_22815;
wire n_22816;
wire n_22817;
wire n_22818;
wire n_22819;
wire n_2282;
wire n_22820;
wire n_22821;
wire n_22822;
wire n_22823;
wire n_22824;
wire n_22825;
wire n_22826;
wire n_22827;
wire n_22828;
wire n_22829;
wire n_2283;
wire n_22830;
wire n_22831;
wire n_22832;
wire n_22833;
wire n_22834;
wire n_22835;
wire n_22836;
wire n_22837;
wire n_22838;
wire n_22839;
wire n_2284;
wire n_22840;
wire n_22841;
wire n_22842;
wire n_22843;
wire n_22844;
wire n_22845;
wire n_22846;
wire n_22847;
wire n_22848;
wire n_22849;
wire n_2285;
wire n_22850;
wire n_22851;
wire n_22852;
wire n_22853;
wire n_22854;
wire n_22855;
wire n_22856;
wire n_22857;
wire n_22858;
wire n_22859;
wire n_2286;
wire n_22860;
wire n_22861;
wire n_22862;
wire n_22863;
wire n_22864;
wire n_22865;
wire n_22866;
wire n_22867;
wire n_22868;
wire n_22869;
wire n_2287;
wire n_22870;
wire n_22871;
wire n_22872;
wire n_22873;
wire n_22874;
wire n_22875;
wire n_22876;
wire n_22877;
wire n_22878;
wire n_22879;
wire n_2288;
wire n_22880;
wire n_22881;
wire n_22882;
wire n_22883;
wire n_22884;
wire n_22885;
wire n_22886;
wire n_22887;
wire n_22888;
wire n_22889;
wire n_2289;
wire n_22890;
wire n_22891;
wire n_22892;
wire n_22893;
wire n_22894;
wire n_22895;
wire n_22896;
wire n_22897;
wire n_22898;
wire n_22899;
wire n_229;
wire n_2290;
wire n_22900;
wire n_22901;
wire n_22902;
wire n_22903;
wire n_22904;
wire n_22905;
wire n_22906;
wire n_22907;
wire n_22908;
wire n_22909;
wire n_2291;
wire n_22910;
wire n_22911;
wire n_22912;
wire n_22913;
wire n_22914;
wire n_22915;
wire n_22916;
wire n_22917;
wire n_22918;
wire n_22919;
wire n_2292;
wire n_22920;
wire n_22921;
wire n_22922;
wire n_22923;
wire n_22924;
wire n_22925;
wire n_22926;
wire n_22927;
wire n_22928;
wire n_22929;
wire n_2293;
wire n_22930;
wire n_22931;
wire n_22932;
wire n_22933;
wire n_22934;
wire n_22935;
wire n_22936;
wire n_22937;
wire n_22938;
wire n_22939;
wire n_2294;
wire n_22940;
wire n_22941;
wire n_22942;
wire n_22943;
wire n_22944;
wire n_22945;
wire n_22946;
wire n_22947;
wire n_22949;
wire n_2295;
wire n_22950;
wire n_22951;
wire n_22952;
wire n_22953;
wire n_22954;
wire n_22955;
wire n_22957;
wire n_22958;
wire n_22959;
wire n_2296;
wire n_22960;
wire n_22961;
wire n_22962;
wire n_22963;
wire n_22964;
wire n_22965;
wire n_22966;
wire n_22967;
wire n_22968;
wire n_22969;
wire n_2297;
wire n_22970;
wire n_22971;
wire n_22972;
wire n_22973;
wire n_22974;
wire n_22975;
wire n_22976;
wire n_22977;
wire n_22978;
wire n_22979;
wire n_2298;
wire n_22980;
wire n_22981;
wire n_22982;
wire n_22983;
wire n_22984;
wire n_22985;
wire n_22986;
wire n_22987;
wire n_22988;
wire n_22989;
wire n_2299;
wire n_22990;
wire n_22991;
wire n_22992;
wire n_22993;
wire n_22994;
wire n_22995;
wire n_22996;
wire n_22997;
wire n_22998;
wire n_22999;
wire n_23;
wire n_230;
wire n_2300;
wire n_23000;
wire n_23001;
wire n_23002;
wire n_23003;
wire n_23004;
wire n_23005;
wire n_23006;
wire n_23007;
wire n_23008;
wire n_23009;
wire n_2301;
wire n_23010;
wire n_23011;
wire n_23012;
wire n_23013;
wire n_23014;
wire n_23015;
wire n_23016;
wire n_23017;
wire n_23018;
wire n_23019;
wire n_2302;
wire n_23020;
wire n_23021;
wire n_23022;
wire n_23023;
wire n_23024;
wire n_23025;
wire n_23026;
wire n_23027;
wire n_23028;
wire n_23029;
wire n_2303;
wire n_23030;
wire n_23031;
wire n_23032;
wire n_23033;
wire n_23034;
wire n_23035;
wire n_23036;
wire n_23037;
wire n_23038;
wire n_23039;
wire n_2304;
wire n_23040;
wire n_23041;
wire n_23042;
wire n_23043;
wire n_23044;
wire n_23045;
wire n_23047;
wire n_23048;
wire n_23049;
wire n_23050;
wire n_23051;
wire n_23052;
wire n_23053;
wire n_23054;
wire n_23055;
wire n_23056;
wire n_23057;
wire n_23058;
wire n_23059;
wire n_2306;
wire n_23060;
wire n_23061;
wire n_23062;
wire n_23063;
wire n_23064;
wire n_23065;
wire n_23066;
wire n_23067;
wire n_23068;
wire n_23069;
wire n_2307;
wire n_23070;
wire n_23071;
wire n_23072;
wire n_23073;
wire n_23074;
wire n_23075;
wire n_23077;
wire n_23078;
wire n_23079;
wire n_23080;
wire n_23081;
wire n_23082;
wire n_23083;
wire n_23084;
wire n_23085;
wire n_23086;
wire n_23087;
wire n_23088;
wire n_23089;
wire n_2309;
wire n_23090;
wire n_23091;
wire n_23092;
wire n_23093;
wire n_23094;
wire n_23095;
wire n_23096;
wire n_23097;
wire n_23098;
wire n_23099;
wire n_231;
wire n_2310;
wire n_23100;
wire n_23101;
wire n_23102;
wire n_23103;
wire n_23104;
wire n_23105;
wire n_23106;
wire n_23107;
wire n_23108;
wire n_23109;
wire n_2311;
wire n_23110;
wire n_23111;
wire n_23112;
wire n_23113;
wire n_23114;
wire n_23115;
wire n_23116;
wire n_23117;
wire n_23118;
wire n_23119;
wire n_2312;
wire n_23120;
wire n_23121;
wire n_23122;
wire n_23123;
wire n_23124;
wire n_23125;
wire n_23126;
wire n_23127;
wire n_23128;
wire n_23129;
wire n_2313;
wire n_23130;
wire n_23131;
wire n_23132;
wire n_23133;
wire n_23134;
wire n_23135;
wire n_23136;
wire n_23137;
wire n_23138;
wire n_23139;
wire n_2314;
wire n_23140;
wire n_23141;
wire n_23142;
wire n_23143;
wire n_23144;
wire n_23145;
wire n_23146;
wire n_23147;
wire n_23148;
wire n_23149;
wire n_2315;
wire n_23150;
wire n_23151;
wire n_23152;
wire n_23153;
wire n_23154;
wire n_23155;
wire n_23156;
wire n_23157;
wire n_23158;
wire n_23159;
wire n_2316;
wire n_23160;
wire n_23161;
wire n_23162;
wire n_23163;
wire n_23164;
wire n_23165;
wire n_23166;
wire n_23167;
wire n_23168;
wire n_23169;
wire n_2317;
wire n_23170;
wire n_23171;
wire n_23172;
wire n_23173;
wire n_23174;
wire n_23175;
wire n_23176;
wire n_23177;
wire n_23178;
wire n_23179;
wire n_2318;
wire n_23180;
wire n_23181;
wire n_23182;
wire n_23183;
wire n_23184;
wire n_23185;
wire n_23186;
wire n_23187;
wire n_23188;
wire n_23189;
wire n_2319;
wire n_23190;
wire n_23191;
wire n_23192;
wire n_23193;
wire n_23194;
wire n_23195;
wire n_23196;
wire n_23197;
wire n_23198;
wire n_23199;
wire n_232;
wire n_2320;
wire n_23200;
wire n_23201;
wire n_23202;
wire n_23203;
wire n_23204;
wire n_23205;
wire n_23206;
wire n_23207;
wire n_23208;
wire n_23209;
wire n_2321;
wire n_23210;
wire n_23211;
wire n_23212;
wire n_23213;
wire n_23214;
wire n_23215;
wire n_23216;
wire n_23217;
wire n_23218;
wire n_23219;
wire n_2322;
wire n_23220;
wire n_23221;
wire n_23222;
wire n_23223;
wire n_23224;
wire n_23225;
wire n_23226;
wire n_23227;
wire n_23228;
wire n_23229;
wire n_2323;
wire n_23230;
wire n_23231;
wire n_23232;
wire n_23233;
wire n_23234;
wire n_23235;
wire n_23236;
wire n_23237;
wire n_23238;
wire n_23239;
wire n_2324;
wire n_23240;
wire n_23241;
wire n_23242;
wire n_23243;
wire n_23244;
wire n_23245;
wire n_23246;
wire n_23247;
wire n_23248;
wire n_23249;
wire n_2325;
wire n_23250;
wire n_23251;
wire n_23252;
wire n_23253;
wire n_23254;
wire n_23255;
wire n_23256;
wire n_23257;
wire n_23258;
wire n_23259;
wire n_2326;
wire n_23260;
wire n_23261;
wire n_23262;
wire n_23263;
wire n_23264;
wire n_23265;
wire n_23266;
wire n_23267;
wire n_23268;
wire n_23269;
wire n_2327;
wire n_23270;
wire n_23271;
wire n_23272;
wire n_23273;
wire n_23274;
wire n_23275;
wire n_23276;
wire n_23277;
wire n_23278;
wire n_23279;
wire n_2328;
wire n_23280;
wire n_23281;
wire n_23282;
wire n_23283;
wire n_23284;
wire n_23285;
wire n_23286;
wire n_23287;
wire n_23288;
wire n_23289;
wire n_2329;
wire n_23290;
wire n_23291;
wire n_23292;
wire n_23293;
wire n_23294;
wire n_23295;
wire n_23296;
wire n_23297;
wire n_23298;
wire n_23299;
wire n_233;
wire n_2330;
wire n_23300;
wire n_23301;
wire n_23302;
wire n_23305;
wire n_23306;
wire n_23307;
wire n_23308;
wire n_23309;
wire n_2331;
wire n_23310;
wire n_23311;
wire n_23312;
wire n_23313;
wire n_23314;
wire n_23315;
wire n_23316;
wire n_23317;
wire n_23318;
wire n_23319;
wire n_2332;
wire n_23320;
wire n_23321;
wire n_23322;
wire n_23323;
wire n_23324;
wire n_23325;
wire n_23326;
wire n_23327;
wire n_23328;
wire n_23329;
wire n_2333;
wire n_23330;
wire n_23331;
wire n_23332;
wire n_23333;
wire n_23334;
wire n_23335;
wire n_23336;
wire n_23337;
wire n_23338;
wire n_23339;
wire n_2334;
wire n_23340;
wire n_23341;
wire n_23342;
wire n_23343;
wire n_23344;
wire n_23345;
wire n_23346;
wire n_23347;
wire n_23348;
wire n_23349;
wire n_2335;
wire n_23350;
wire n_23351;
wire n_23352;
wire n_23353;
wire n_23354;
wire n_23355;
wire n_23356;
wire n_23357;
wire n_23358;
wire n_23359;
wire n_2336;
wire n_23360;
wire n_23361;
wire n_23362;
wire n_23363;
wire n_23364;
wire n_23365;
wire n_23366;
wire n_23367;
wire n_23369;
wire n_2337;
wire n_23370;
wire n_23371;
wire n_23372;
wire n_23373;
wire n_23374;
wire n_23375;
wire n_23376;
wire n_23377;
wire n_23378;
wire n_23379;
wire n_2338;
wire n_23380;
wire n_23381;
wire n_23382;
wire n_23383;
wire n_23384;
wire n_23385;
wire n_23386;
wire n_23387;
wire n_23388;
wire n_23389;
wire n_2339;
wire n_23390;
wire n_23391;
wire n_23392;
wire n_23393;
wire n_23394;
wire n_23395;
wire n_23396;
wire n_23397;
wire n_23398;
wire n_23399;
wire n_234;
wire n_2340;
wire n_23400;
wire n_23401;
wire n_23402;
wire n_23403;
wire n_23404;
wire n_23405;
wire n_23406;
wire n_23408;
wire n_23409;
wire n_2341;
wire n_23410;
wire n_23411;
wire n_23412;
wire n_23413;
wire n_23414;
wire n_23415;
wire n_23416;
wire n_23417;
wire n_23418;
wire n_23419;
wire n_2342;
wire n_23420;
wire n_23421;
wire n_23422;
wire n_23423;
wire n_23424;
wire n_23425;
wire n_23426;
wire n_23427;
wire n_23428;
wire n_23429;
wire n_2343;
wire n_23430;
wire n_23431;
wire n_23432;
wire n_23433;
wire n_23434;
wire n_23435;
wire n_23436;
wire n_23437;
wire n_23438;
wire n_23439;
wire n_2344;
wire n_23440;
wire n_23441;
wire n_23442;
wire n_23443;
wire n_23444;
wire n_23445;
wire n_23446;
wire n_23447;
wire n_23448;
wire n_23449;
wire n_2345;
wire n_23450;
wire n_23451;
wire n_23452;
wire n_23453;
wire n_23454;
wire n_23455;
wire n_23456;
wire n_23457;
wire n_23458;
wire n_23459;
wire n_2346;
wire n_23460;
wire n_23461;
wire n_23462;
wire n_23463;
wire n_23464;
wire n_23465;
wire n_23466;
wire n_23467;
wire n_23468;
wire n_23469;
wire n_2347;
wire n_23470;
wire n_23471;
wire n_23472;
wire n_23473;
wire n_23474;
wire n_23475;
wire n_23476;
wire n_23477;
wire n_23478;
wire n_23479;
wire n_2348;
wire n_23480;
wire n_23481;
wire n_23482;
wire n_23483;
wire n_23484;
wire n_23485;
wire n_23486;
wire n_23487;
wire n_23488;
wire n_23489;
wire n_2349;
wire n_23490;
wire n_23491;
wire n_23492;
wire n_23493;
wire n_23494;
wire n_23495;
wire n_23496;
wire n_23497;
wire n_23498;
wire n_23499;
wire n_235;
wire n_2350;
wire n_23500;
wire n_23501;
wire n_23502;
wire n_23503;
wire n_23504;
wire n_23505;
wire n_23506;
wire n_23507;
wire n_23508;
wire n_23509;
wire n_2351;
wire n_23510;
wire n_23511;
wire n_23512;
wire n_23513;
wire n_23514;
wire n_23515;
wire n_23516;
wire n_23517;
wire n_23518;
wire n_23519;
wire n_2352;
wire n_23520;
wire n_23521;
wire n_23522;
wire n_23523;
wire n_23524;
wire n_23525;
wire n_23526;
wire n_23527;
wire n_23528;
wire n_23529;
wire n_2353;
wire n_23530;
wire n_23531;
wire n_23532;
wire n_23533;
wire n_23534;
wire n_23535;
wire n_23536;
wire n_23537;
wire n_23538;
wire n_23539;
wire n_2354;
wire n_23540;
wire n_23541;
wire n_23542;
wire n_23543;
wire n_23544;
wire n_23545;
wire n_23546;
wire n_23547;
wire n_23548;
wire n_23549;
wire n_2355;
wire n_23551;
wire n_23552;
wire n_23553;
wire n_23554;
wire n_23555;
wire n_23556;
wire n_23557;
wire n_23558;
wire n_23559;
wire n_2356;
wire n_23560;
wire n_23561;
wire n_23562;
wire n_23563;
wire n_23564;
wire n_23565;
wire n_23566;
wire n_23567;
wire n_23568;
wire n_23569;
wire n_2357;
wire n_23570;
wire n_23571;
wire n_23572;
wire n_23573;
wire n_23574;
wire n_23575;
wire n_23576;
wire n_23577;
wire n_23578;
wire n_23579;
wire n_23580;
wire n_23581;
wire n_23582;
wire n_23583;
wire n_23584;
wire n_23585;
wire n_23586;
wire n_23587;
wire n_23588;
wire n_23589;
wire n_2359;
wire n_23590;
wire n_23591;
wire n_23592;
wire n_23593;
wire n_23594;
wire n_23595;
wire n_23596;
wire n_23597;
wire n_23598;
wire n_23599;
wire n_236;
wire n_2360;
wire n_23600;
wire n_23601;
wire n_23602;
wire n_23603;
wire n_23604;
wire n_23605;
wire n_23606;
wire n_23607;
wire n_23609;
wire n_2361;
wire n_23610;
wire n_23611;
wire n_23612;
wire n_23614;
wire n_23615;
wire n_23616;
wire n_23617;
wire n_23618;
wire n_23619;
wire n_2362;
wire n_23620;
wire n_23621;
wire n_23622;
wire n_23623;
wire n_23624;
wire n_23625;
wire n_23626;
wire n_23627;
wire n_23628;
wire n_23629;
wire n_2363;
wire n_23630;
wire n_23631;
wire n_23632;
wire n_23633;
wire n_23634;
wire n_23635;
wire n_23636;
wire n_23637;
wire n_23638;
wire n_23639;
wire n_2364;
wire n_23640;
wire n_23641;
wire n_23642;
wire n_23643;
wire n_23644;
wire n_23645;
wire n_23646;
wire n_23647;
wire n_23648;
wire n_23649;
wire n_2365;
wire n_23650;
wire n_23651;
wire n_23652;
wire n_23653;
wire n_23655;
wire n_23656;
wire n_23657;
wire n_23658;
wire n_23659;
wire n_2366;
wire n_23660;
wire n_23661;
wire n_23662;
wire n_23663;
wire n_23664;
wire n_23665;
wire n_23666;
wire n_23667;
wire n_23668;
wire n_23669;
wire n_2367;
wire n_23670;
wire n_23671;
wire n_23672;
wire n_23673;
wire n_23674;
wire n_23675;
wire n_23676;
wire n_23677;
wire n_23678;
wire n_23679;
wire n_2368;
wire n_23680;
wire n_23681;
wire n_23682;
wire n_23683;
wire n_23684;
wire n_23685;
wire n_23686;
wire n_23687;
wire n_23688;
wire n_23689;
wire n_2369;
wire n_23690;
wire n_23691;
wire n_23692;
wire n_23693;
wire n_23694;
wire n_23695;
wire n_23696;
wire n_23697;
wire n_23698;
wire n_23699;
wire n_237;
wire n_2370;
wire n_23700;
wire n_23701;
wire n_23702;
wire n_23703;
wire n_23704;
wire n_23705;
wire n_23706;
wire n_23707;
wire n_23708;
wire n_23709;
wire n_2371;
wire n_23710;
wire n_23711;
wire n_23713;
wire n_23714;
wire n_23715;
wire n_23716;
wire n_23717;
wire n_23718;
wire n_23719;
wire n_2372;
wire n_23720;
wire n_23721;
wire n_23722;
wire n_23723;
wire n_23724;
wire n_23725;
wire n_23726;
wire n_23727;
wire n_23728;
wire n_23729;
wire n_2373;
wire n_23730;
wire n_23731;
wire n_23732;
wire n_23733;
wire n_23734;
wire n_23735;
wire n_23736;
wire n_23737;
wire n_23738;
wire n_23739;
wire n_2374;
wire n_23740;
wire n_23741;
wire n_23742;
wire n_23743;
wire n_23744;
wire n_23745;
wire n_23746;
wire n_23747;
wire n_23748;
wire n_23749;
wire n_2375;
wire n_23750;
wire n_23751;
wire n_23752;
wire n_23753;
wire n_23754;
wire n_23755;
wire n_23756;
wire n_23757;
wire n_23758;
wire n_23759;
wire n_2376;
wire n_23760;
wire n_23761;
wire n_23762;
wire n_23763;
wire n_23764;
wire n_23765;
wire n_23766;
wire n_23767;
wire n_23768;
wire n_23769;
wire n_2377;
wire n_23770;
wire n_23771;
wire n_23772;
wire n_23773;
wire n_23774;
wire n_23775;
wire n_23776;
wire n_23777;
wire n_23778;
wire n_23779;
wire n_2378;
wire n_23780;
wire n_23781;
wire n_23782;
wire n_23783;
wire n_23784;
wire n_23785;
wire n_23786;
wire n_23787;
wire n_23788;
wire n_23789;
wire n_2379;
wire n_23790;
wire n_23791;
wire n_23792;
wire n_23793;
wire n_23794;
wire n_23795;
wire n_23796;
wire n_23797;
wire n_23798;
wire n_23799;
wire n_238;
wire n_2380;
wire n_23800;
wire n_23801;
wire n_23802;
wire n_23803;
wire n_23804;
wire n_23806;
wire n_23807;
wire n_23808;
wire n_23809;
wire n_2381;
wire n_23810;
wire n_23811;
wire n_23812;
wire n_23813;
wire n_23814;
wire n_23815;
wire n_23816;
wire n_23817;
wire n_23818;
wire n_23819;
wire n_2382;
wire n_23820;
wire n_23821;
wire n_23822;
wire n_23823;
wire n_23824;
wire n_23825;
wire n_23826;
wire n_23827;
wire n_23828;
wire n_23829;
wire n_2383;
wire n_23830;
wire n_23831;
wire n_23832;
wire n_23833;
wire n_23834;
wire n_23835;
wire n_23836;
wire n_23837;
wire n_23838;
wire n_23839;
wire n_2384;
wire n_23840;
wire n_23841;
wire n_23842;
wire n_23843;
wire n_23844;
wire n_23845;
wire n_23846;
wire n_23847;
wire n_23848;
wire n_23849;
wire n_2385;
wire n_23850;
wire n_23851;
wire n_23852;
wire n_23853;
wire n_23854;
wire n_23855;
wire n_23856;
wire n_23857;
wire n_23858;
wire n_23859;
wire n_23860;
wire n_23861;
wire n_23862;
wire n_23863;
wire n_23864;
wire n_23865;
wire n_23866;
wire n_23867;
wire n_23868;
wire n_23869;
wire n_2387;
wire n_23870;
wire n_23871;
wire n_23872;
wire n_23873;
wire n_23874;
wire n_23875;
wire n_23876;
wire n_23877;
wire n_23878;
wire n_23879;
wire n_2388;
wire n_23880;
wire n_23881;
wire n_23882;
wire n_23883;
wire n_23884;
wire n_23885;
wire n_23886;
wire n_23887;
wire n_23888;
wire n_23889;
wire n_2389;
wire n_23890;
wire n_23891;
wire n_23892;
wire n_23893;
wire n_23894;
wire n_23895;
wire n_23896;
wire n_23897;
wire n_23898;
wire n_23899;
wire n_239;
wire n_2390;
wire n_23900;
wire n_23901;
wire n_23902;
wire n_23903;
wire n_23904;
wire n_23905;
wire n_23906;
wire n_23907;
wire n_23908;
wire n_23909;
wire n_2391;
wire n_23910;
wire n_23911;
wire n_23912;
wire n_23913;
wire n_23914;
wire n_23915;
wire n_23916;
wire n_23917;
wire n_23918;
wire n_23919;
wire n_2392;
wire n_23920;
wire n_23921;
wire n_23922;
wire n_23923;
wire n_23924;
wire n_23925;
wire n_23926;
wire n_23927;
wire n_23928;
wire n_23929;
wire n_2393;
wire n_23930;
wire n_23931;
wire n_23932;
wire n_23933;
wire n_23934;
wire n_23936;
wire n_23937;
wire n_23938;
wire n_23939;
wire n_2394;
wire n_23940;
wire n_23941;
wire n_23942;
wire n_23943;
wire n_23944;
wire n_23945;
wire n_23946;
wire n_23947;
wire n_23948;
wire n_23949;
wire n_2395;
wire n_23950;
wire n_23951;
wire n_23952;
wire n_23953;
wire n_23954;
wire n_23955;
wire n_23956;
wire n_23957;
wire n_23958;
wire n_23959;
wire n_2396;
wire n_23960;
wire n_23961;
wire n_23962;
wire n_23963;
wire n_23964;
wire n_23965;
wire n_23966;
wire n_23967;
wire n_23968;
wire n_23969;
wire n_2397;
wire n_23970;
wire n_23971;
wire n_23972;
wire n_23973;
wire n_23974;
wire n_23975;
wire n_23976;
wire n_23977;
wire n_23978;
wire n_23979;
wire n_2398;
wire n_23980;
wire n_23981;
wire n_23982;
wire n_23983;
wire n_23984;
wire n_23985;
wire n_23986;
wire n_23987;
wire n_23988;
wire n_23989;
wire n_2399;
wire n_23990;
wire n_23991;
wire n_23992;
wire n_23993;
wire n_23994;
wire n_23995;
wire n_23996;
wire n_23997;
wire n_23998;
wire n_23999;
wire n_24;
wire n_240;
wire n_2400;
wire n_24000;
wire n_24001;
wire n_24002;
wire n_24003;
wire n_24004;
wire n_24005;
wire n_24006;
wire n_24007;
wire n_24008;
wire n_24009;
wire n_2401;
wire n_24010;
wire n_24011;
wire n_24012;
wire n_24013;
wire n_24014;
wire n_24015;
wire n_24016;
wire n_24017;
wire n_24018;
wire n_24019;
wire n_2402;
wire n_24020;
wire n_24021;
wire n_24022;
wire n_24023;
wire n_24024;
wire n_24025;
wire n_24026;
wire n_24027;
wire n_24028;
wire n_24029;
wire n_2403;
wire n_24030;
wire n_24031;
wire n_24032;
wire n_24033;
wire n_24034;
wire n_24035;
wire n_24036;
wire n_24037;
wire n_24038;
wire n_24039;
wire n_2404;
wire n_24040;
wire n_24041;
wire n_24042;
wire n_24043;
wire n_24044;
wire n_24045;
wire n_24046;
wire n_24047;
wire n_24048;
wire n_24049;
wire n_2405;
wire n_24050;
wire n_24051;
wire n_24052;
wire n_24053;
wire n_24054;
wire n_24055;
wire n_24056;
wire n_24057;
wire n_24058;
wire n_24059;
wire n_2406;
wire n_24060;
wire n_24061;
wire n_24062;
wire n_24063;
wire n_24064;
wire n_24065;
wire n_24066;
wire n_24067;
wire n_24068;
wire n_24069;
wire n_2407;
wire n_24070;
wire n_24071;
wire n_24072;
wire n_24073;
wire n_24074;
wire n_24075;
wire n_24076;
wire n_24077;
wire n_24078;
wire n_24079;
wire n_2408;
wire n_24080;
wire n_24081;
wire n_24082;
wire n_24083;
wire n_24084;
wire n_24085;
wire n_24086;
wire n_24087;
wire n_24088;
wire n_24089;
wire n_2409;
wire n_24090;
wire n_24091;
wire n_24092;
wire n_24093;
wire n_24094;
wire n_24095;
wire n_24096;
wire n_24097;
wire n_24098;
wire n_24099;
wire n_241;
wire n_2410;
wire n_24100;
wire n_24101;
wire n_24102;
wire n_24103;
wire n_24104;
wire n_24105;
wire n_24106;
wire n_24107;
wire n_24108;
wire n_24109;
wire n_2411;
wire n_24110;
wire n_24111;
wire n_24112;
wire n_24113;
wire n_24114;
wire n_24115;
wire n_24116;
wire n_24117;
wire n_24118;
wire n_24119;
wire n_2412;
wire n_24120;
wire n_24121;
wire n_24122;
wire n_24123;
wire n_24124;
wire n_24125;
wire n_24126;
wire n_24127;
wire n_24128;
wire n_24129;
wire n_2413;
wire n_24130;
wire n_24131;
wire n_24132;
wire n_24133;
wire n_24134;
wire n_24135;
wire n_24136;
wire n_24137;
wire n_24138;
wire n_24139;
wire n_2414;
wire n_24140;
wire n_24141;
wire n_24142;
wire n_24143;
wire n_24144;
wire n_24145;
wire n_24146;
wire n_24147;
wire n_24148;
wire n_24149;
wire n_2415;
wire n_24150;
wire n_24151;
wire n_24152;
wire n_24153;
wire n_24154;
wire n_24155;
wire n_24156;
wire n_24157;
wire n_24158;
wire n_24159;
wire n_2416;
wire n_24160;
wire n_24161;
wire n_24162;
wire n_24163;
wire n_24164;
wire n_24166;
wire n_24167;
wire n_24168;
wire n_24169;
wire n_2417;
wire n_24170;
wire n_24171;
wire n_24172;
wire n_24173;
wire n_24174;
wire n_24175;
wire n_24176;
wire n_24177;
wire n_24178;
wire n_24179;
wire n_24180;
wire n_24181;
wire n_24182;
wire n_24183;
wire n_24184;
wire n_24185;
wire n_24186;
wire n_24187;
wire n_24188;
wire n_24189;
wire n_2419;
wire n_24190;
wire n_24191;
wire n_24192;
wire n_24193;
wire n_24194;
wire n_24195;
wire n_24196;
wire n_24197;
wire n_24198;
wire n_24199;
wire n_242;
wire n_2420;
wire n_24200;
wire n_24201;
wire n_24202;
wire n_24203;
wire n_24204;
wire n_24205;
wire n_24206;
wire n_24207;
wire n_24208;
wire n_24209;
wire n_2421;
wire n_24210;
wire n_24211;
wire n_24212;
wire n_24213;
wire n_24214;
wire n_24215;
wire n_24216;
wire n_24217;
wire n_24218;
wire n_24219;
wire n_2422;
wire n_24220;
wire n_24221;
wire n_24222;
wire n_24223;
wire n_24224;
wire n_24225;
wire n_24226;
wire n_24227;
wire n_24228;
wire n_24229;
wire n_2423;
wire n_24230;
wire n_24231;
wire n_24232;
wire n_24233;
wire n_24234;
wire n_24235;
wire n_24236;
wire n_24237;
wire n_24238;
wire n_24239;
wire n_2424;
wire n_24240;
wire n_24241;
wire n_24242;
wire n_24243;
wire n_24244;
wire n_24245;
wire n_24246;
wire n_24247;
wire n_24248;
wire n_24249;
wire n_2425;
wire n_24250;
wire n_24251;
wire n_24252;
wire n_24253;
wire n_24254;
wire n_24255;
wire n_24256;
wire n_24257;
wire n_24258;
wire n_24259;
wire n_2426;
wire n_24260;
wire n_24261;
wire n_24262;
wire n_24263;
wire n_24264;
wire n_24265;
wire n_24266;
wire n_24267;
wire n_24268;
wire n_24269;
wire n_24270;
wire n_24271;
wire n_24272;
wire n_24273;
wire n_24274;
wire n_24275;
wire n_24276;
wire n_24277;
wire n_24278;
wire n_24279;
wire n_2428;
wire n_24280;
wire n_24281;
wire n_24282;
wire n_24283;
wire n_24284;
wire n_24285;
wire n_24286;
wire n_24287;
wire n_24288;
wire n_24289;
wire n_2429;
wire n_24290;
wire n_24291;
wire n_24292;
wire n_24293;
wire n_24294;
wire n_24295;
wire n_24296;
wire n_24297;
wire n_24298;
wire n_24299;
wire n_243;
wire n_2430;
wire n_24300;
wire n_24301;
wire n_24302;
wire n_24303;
wire n_24304;
wire n_24305;
wire n_24306;
wire n_24307;
wire n_24308;
wire n_24309;
wire n_2431;
wire n_24310;
wire n_24311;
wire n_24312;
wire n_24313;
wire n_24314;
wire n_24315;
wire n_24316;
wire n_24317;
wire n_24318;
wire n_24319;
wire n_2432;
wire n_24320;
wire n_24321;
wire n_24322;
wire n_24323;
wire n_24324;
wire n_24325;
wire n_24326;
wire n_24327;
wire n_24328;
wire n_24329;
wire n_2433;
wire n_24330;
wire n_24331;
wire n_24332;
wire n_24333;
wire n_24334;
wire n_24335;
wire n_24336;
wire n_24337;
wire n_24338;
wire n_24339;
wire n_2434;
wire n_24340;
wire n_24341;
wire n_24342;
wire n_24343;
wire n_24344;
wire n_24345;
wire n_24346;
wire n_24347;
wire n_24348;
wire n_24349;
wire n_2435;
wire n_24350;
wire n_24351;
wire n_24352;
wire n_24353;
wire n_24354;
wire n_24355;
wire n_24356;
wire n_24357;
wire n_24358;
wire n_24359;
wire n_2436;
wire n_24360;
wire n_24361;
wire n_24362;
wire n_24363;
wire n_24364;
wire n_24365;
wire n_24366;
wire n_24367;
wire n_24368;
wire n_24369;
wire n_2437;
wire n_24370;
wire n_24371;
wire n_24372;
wire n_24373;
wire n_24374;
wire n_24375;
wire n_24376;
wire n_24377;
wire n_24378;
wire n_24379;
wire n_2438;
wire n_24380;
wire n_24381;
wire n_24382;
wire n_24383;
wire n_24384;
wire n_24385;
wire n_24386;
wire n_24387;
wire n_24388;
wire n_24389;
wire n_2439;
wire n_24390;
wire n_24391;
wire n_24392;
wire n_24393;
wire n_24394;
wire n_24395;
wire n_24396;
wire n_24397;
wire n_24398;
wire n_24399;
wire n_244;
wire n_2440;
wire n_24400;
wire n_24401;
wire n_24402;
wire n_24403;
wire n_24404;
wire n_24405;
wire n_24406;
wire n_24408;
wire n_24409;
wire n_2441;
wire n_24410;
wire n_24411;
wire n_24412;
wire n_24413;
wire n_24414;
wire n_24415;
wire n_24416;
wire n_24417;
wire n_24418;
wire n_24419;
wire n_2442;
wire n_24420;
wire n_24421;
wire n_24422;
wire n_24423;
wire n_24424;
wire n_24425;
wire n_24426;
wire n_24427;
wire n_24428;
wire n_24429;
wire n_2443;
wire n_24430;
wire n_24431;
wire n_24432;
wire n_24433;
wire n_24434;
wire n_24435;
wire n_24436;
wire n_24437;
wire n_24438;
wire n_24439;
wire n_2444;
wire n_24440;
wire n_24441;
wire n_24442;
wire n_24443;
wire n_24444;
wire n_24445;
wire n_24446;
wire n_24447;
wire n_24448;
wire n_24449;
wire n_2445;
wire n_24450;
wire n_24451;
wire n_24452;
wire n_24453;
wire n_24454;
wire n_24455;
wire n_24456;
wire n_24457;
wire n_24458;
wire n_24459;
wire n_2446;
wire n_24460;
wire n_24461;
wire n_24462;
wire n_24463;
wire n_24464;
wire n_24465;
wire n_24466;
wire n_24467;
wire n_24468;
wire n_24469;
wire n_2447;
wire n_24470;
wire n_24471;
wire n_24472;
wire n_24473;
wire n_24474;
wire n_24475;
wire n_24476;
wire n_24477;
wire n_24478;
wire n_24479;
wire n_2448;
wire n_24480;
wire n_24481;
wire n_24482;
wire n_24483;
wire n_24484;
wire n_24485;
wire n_24486;
wire n_24487;
wire n_24488;
wire n_24489;
wire n_2449;
wire n_24490;
wire n_24491;
wire n_24492;
wire n_24493;
wire n_24494;
wire n_24495;
wire n_24496;
wire n_24497;
wire n_24498;
wire n_24499;
wire n_245;
wire n_2450;
wire n_24500;
wire n_24501;
wire n_24502;
wire n_24503;
wire n_24504;
wire n_24505;
wire n_24506;
wire n_24507;
wire n_24508;
wire n_24509;
wire n_2451;
wire n_24510;
wire n_24511;
wire n_24512;
wire n_24513;
wire n_24514;
wire n_24515;
wire n_24516;
wire n_24517;
wire n_24518;
wire n_2452;
wire n_24520;
wire n_24521;
wire n_24522;
wire n_24523;
wire n_24524;
wire n_24525;
wire n_24526;
wire n_24527;
wire n_24528;
wire n_24529;
wire n_2453;
wire n_24530;
wire n_24531;
wire n_24532;
wire n_24533;
wire n_24534;
wire n_24535;
wire n_24536;
wire n_24537;
wire n_24538;
wire n_24539;
wire n_2454;
wire n_24540;
wire n_24541;
wire n_24542;
wire n_24543;
wire n_24544;
wire n_24545;
wire n_24546;
wire n_24547;
wire n_24548;
wire n_24549;
wire n_2455;
wire n_24550;
wire n_24551;
wire n_24552;
wire n_24553;
wire n_24554;
wire n_24555;
wire n_24556;
wire n_24557;
wire n_24558;
wire n_24559;
wire n_2456;
wire n_24560;
wire n_24561;
wire n_24562;
wire n_24563;
wire n_24564;
wire n_24565;
wire n_24566;
wire n_24567;
wire n_24568;
wire n_24569;
wire n_2457;
wire n_24570;
wire n_24571;
wire n_24572;
wire n_24573;
wire n_24574;
wire n_24575;
wire n_24576;
wire n_24577;
wire n_24578;
wire n_24579;
wire n_2458;
wire n_24580;
wire n_24581;
wire n_24582;
wire n_24583;
wire n_24584;
wire n_24585;
wire n_24586;
wire n_24587;
wire n_24588;
wire n_24589;
wire n_2459;
wire n_24590;
wire n_24591;
wire n_24592;
wire n_24593;
wire n_24594;
wire n_24595;
wire n_24596;
wire n_24598;
wire n_246;
wire n_2460;
wire n_24600;
wire n_24601;
wire n_24603;
wire n_24604;
wire n_24605;
wire n_24606;
wire n_24608;
wire n_24609;
wire n_2461;
wire n_24610;
wire n_24611;
wire n_24612;
wire n_24613;
wire n_24614;
wire n_24616;
wire n_24617;
wire n_24618;
wire n_24619;
wire n_2462;
wire n_24620;
wire n_24621;
wire n_24623;
wire n_24624;
wire n_24625;
wire n_24626;
wire n_24627;
wire n_24628;
wire n_24629;
wire n_2463;
wire n_24630;
wire n_24631;
wire n_24632;
wire n_24633;
wire n_24634;
wire n_24635;
wire n_24636;
wire n_24637;
wire n_24638;
wire n_24639;
wire n_2464;
wire n_24640;
wire n_24641;
wire n_24642;
wire n_24643;
wire n_24644;
wire n_24645;
wire n_24646;
wire n_24647;
wire n_24648;
wire n_24649;
wire n_2465;
wire n_24650;
wire n_24651;
wire n_24652;
wire n_24653;
wire n_24654;
wire n_24655;
wire n_24656;
wire n_24657;
wire n_24658;
wire n_24659;
wire n_2466;
wire n_24660;
wire n_24661;
wire n_24662;
wire n_24663;
wire n_24665;
wire n_24666;
wire n_24667;
wire n_24668;
wire n_24669;
wire n_2467;
wire n_24670;
wire n_24671;
wire n_24672;
wire n_24673;
wire n_24674;
wire n_24675;
wire n_24676;
wire n_24677;
wire n_24678;
wire n_24679;
wire n_2468;
wire n_24680;
wire n_24681;
wire n_24682;
wire n_24683;
wire n_24684;
wire n_24685;
wire n_24686;
wire n_24687;
wire n_24688;
wire n_24689;
wire n_2469;
wire n_24690;
wire n_24691;
wire n_24692;
wire n_24693;
wire n_24694;
wire n_24695;
wire n_24697;
wire n_24698;
wire n_24699;
wire n_247;
wire n_2470;
wire n_24700;
wire n_24701;
wire n_24702;
wire n_24703;
wire n_24704;
wire n_24705;
wire n_24706;
wire n_24707;
wire n_24708;
wire n_24709;
wire n_2471;
wire n_24711;
wire n_24712;
wire n_24713;
wire n_24714;
wire n_24715;
wire n_24716;
wire n_24717;
wire n_24718;
wire n_24719;
wire n_2472;
wire n_24720;
wire n_24721;
wire n_24722;
wire n_24723;
wire n_24724;
wire n_24725;
wire n_24726;
wire n_24727;
wire n_24728;
wire n_24729;
wire n_2473;
wire n_24730;
wire n_24731;
wire n_24732;
wire n_24733;
wire n_24734;
wire n_24735;
wire n_24736;
wire n_24737;
wire n_24738;
wire n_24739;
wire n_2474;
wire n_24740;
wire n_24742;
wire n_24743;
wire n_24744;
wire n_24745;
wire n_24746;
wire n_24747;
wire n_24748;
wire n_24749;
wire n_2475;
wire n_24750;
wire n_24751;
wire n_24752;
wire n_24753;
wire n_24754;
wire n_24755;
wire n_24756;
wire n_24757;
wire n_24758;
wire n_24759;
wire n_2476;
wire n_24760;
wire n_24761;
wire n_24762;
wire n_24763;
wire n_24764;
wire n_24765;
wire n_24766;
wire n_24767;
wire n_24768;
wire n_24769;
wire n_2477;
wire n_24770;
wire n_24771;
wire n_24772;
wire n_24773;
wire n_24774;
wire n_24775;
wire n_24776;
wire n_24777;
wire n_24778;
wire n_24779;
wire n_2478;
wire n_24780;
wire n_24781;
wire n_24782;
wire n_24783;
wire n_24784;
wire n_24785;
wire n_24786;
wire n_24787;
wire n_24788;
wire n_24789;
wire n_2479;
wire n_24790;
wire n_24791;
wire n_24792;
wire n_24793;
wire n_24794;
wire n_24795;
wire n_24796;
wire n_24797;
wire n_24798;
wire n_24799;
wire n_248;
wire n_2480;
wire n_24800;
wire n_24801;
wire n_24802;
wire n_24803;
wire n_24804;
wire n_24805;
wire n_24806;
wire n_24807;
wire n_24808;
wire n_24809;
wire n_2481;
wire n_24810;
wire n_24811;
wire n_24812;
wire n_24813;
wire n_24814;
wire n_24815;
wire n_24816;
wire n_24817;
wire n_24819;
wire n_2482;
wire n_24820;
wire n_24821;
wire n_24822;
wire n_24823;
wire n_24824;
wire n_24825;
wire n_24826;
wire n_24827;
wire n_24828;
wire n_24829;
wire n_2483;
wire n_24830;
wire n_24831;
wire n_24832;
wire n_24833;
wire n_24834;
wire n_24835;
wire n_24837;
wire n_24838;
wire n_24839;
wire n_2484;
wire n_24840;
wire n_24841;
wire n_24842;
wire n_24843;
wire n_24844;
wire n_24845;
wire n_24846;
wire n_24847;
wire n_24848;
wire n_24849;
wire n_2485;
wire n_24850;
wire n_24851;
wire n_24852;
wire n_24853;
wire n_24854;
wire n_24855;
wire n_24856;
wire n_24857;
wire n_24858;
wire n_24859;
wire n_2486;
wire n_24860;
wire n_24861;
wire n_24862;
wire n_24863;
wire n_24864;
wire n_24865;
wire n_24866;
wire n_24867;
wire n_24868;
wire n_24869;
wire n_2487;
wire n_24870;
wire n_24871;
wire n_24872;
wire n_24873;
wire n_24874;
wire n_24875;
wire n_24876;
wire n_24877;
wire n_24878;
wire n_24879;
wire n_2488;
wire n_24880;
wire n_24881;
wire n_24882;
wire n_24883;
wire n_24884;
wire n_24885;
wire n_24886;
wire n_24887;
wire n_24888;
wire n_24889;
wire n_2489;
wire n_24890;
wire n_24891;
wire n_24892;
wire n_24893;
wire n_24894;
wire n_24895;
wire n_24896;
wire n_24897;
wire n_24898;
wire n_24899;
wire n_249;
wire n_2490;
wire n_24900;
wire n_24901;
wire n_24902;
wire n_24903;
wire n_24904;
wire n_24905;
wire n_24906;
wire n_24907;
wire n_24908;
wire n_24909;
wire n_2491;
wire n_24910;
wire n_24911;
wire n_24912;
wire n_24913;
wire n_24914;
wire n_24915;
wire n_24916;
wire n_24917;
wire n_24918;
wire n_24919;
wire n_2492;
wire n_24920;
wire n_24921;
wire n_24923;
wire n_24924;
wire n_24925;
wire n_24926;
wire n_24927;
wire n_24928;
wire n_24929;
wire n_2493;
wire n_24930;
wire n_24931;
wire n_24932;
wire n_24933;
wire n_24934;
wire n_24935;
wire n_24936;
wire n_24937;
wire n_24938;
wire n_24939;
wire n_2494;
wire n_24940;
wire n_24941;
wire n_24942;
wire n_24943;
wire n_24944;
wire n_24945;
wire n_24946;
wire n_24947;
wire n_24948;
wire n_24949;
wire n_2495;
wire n_24950;
wire n_24951;
wire n_24952;
wire n_24953;
wire n_24954;
wire n_24955;
wire n_24956;
wire n_24957;
wire n_24958;
wire n_24959;
wire n_2496;
wire n_24960;
wire n_24961;
wire n_24962;
wire n_24963;
wire n_24964;
wire n_24965;
wire n_24966;
wire n_24967;
wire n_24968;
wire n_24969;
wire n_2497;
wire n_24970;
wire n_24971;
wire n_24972;
wire n_24973;
wire n_24974;
wire n_24975;
wire n_24976;
wire n_24977;
wire n_24978;
wire n_24979;
wire n_2498;
wire n_24980;
wire n_24981;
wire n_24982;
wire n_24983;
wire n_24985;
wire n_24986;
wire n_24987;
wire n_24988;
wire n_24989;
wire n_2499;
wire n_24990;
wire n_24991;
wire n_24992;
wire n_24993;
wire n_24994;
wire n_24995;
wire n_24996;
wire n_24997;
wire n_24998;
wire n_24999;
wire n_25;
wire n_250;
wire n_2500;
wire n_25000;
wire n_25001;
wire n_25002;
wire n_25003;
wire n_25004;
wire n_25005;
wire n_25006;
wire n_25007;
wire n_25008;
wire n_25009;
wire n_2501;
wire n_25010;
wire n_25011;
wire n_25012;
wire n_25013;
wire n_25014;
wire n_25015;
wire n_25016;
wire n_25017;
wire n_25018;
wire n_25019;
wire n_2502;
wire n_25020;
wire n_25021;
wire n_25022;
wire n_25023;
wire n_25024;
wire n_25025;
wire n_25026;
wire n_25027;
wire n_25028;
wire n_25029;
wire n_2503;
wire n_25030;
wire n_25031;
wire n_25032;
wire n_25033;
wire n_25034;
wire n_25035;
wire n_25036;
wire n_25038;
wire n_25039;
wire n_2504;
wire n_25040;
wire n_25041;
wire n_25042;
wire n_25043;
wire n_25044;
wire n_25045;
wire n_25046;
wire n_25047;
wire n_25048;
wire n_25049;
wire n_2505;
wire n_25050;
wire n_25051;
wire n_25052;
wire n_25053;
wire n_25054;
wire n_25055;
wire n_25056;
wire n_25057;
wire n_25058;
wire n_25059;
wire n_2506;
wire n_25060;
wire n_25061;
wire n_25062;
wire n_25063;
wire n_25064;
wire n_25065;
wire n_25066;
wire n_25067;
wire n_25068;
wire n_25069;
wire n_2507;
wire n_25070;
wire n_25071;
wire n_25072;
wire n_25073;
wire n_25074;
wire n_25075;
wire n_25076;
wire n_25077;
wire n_25078;
wire n_25079;
wire n_2508;
wire n_25080;
wire n_25081;
wire n_25082;
wire n_25083;
wire n_25084;
wire n_25085;
wire n_25086;
wire n_25087;
wire n_25088;
wire n_25089;
wire n_2509;
wire n_25090;
wire n_25091;
wire n_25092;
wire n_25093;
wire n_25095;
wire n_25096;
wire n_25097;
wire n_25098;
wire n_25099;
wire n_251;
wire n_25100;
wire n_25101;
wire n_25102;
wire n_25103;
wire n_25104;
wire n_25105;
wire n_25106;
wire n_25107;
wire n_25108;
wire n_25109;
wire n_2511;
wire n_25110;
wire n_25111;
wire n_25112;
wire n_25113;
wire n_25114;
wire n_25115;
wire n_25116;
wire n_25117;
wire n_25118;
wire n_25119;
wire n_2512;
wire n_25120;
wire n_25121;
wire n_25122;
wire n_25123;
wire n_25124;
wire n_25125;
wire n_25126;
wire n_25127;
wire n_25128;
wire n_25129;
wire n_2513;
wire n_25130;
wire n_25131;
wire n_25132;
wire n_25133;
wire n_25134;
wire n_25135;
wire n_25136;
wire n_25137;
wire n_25138;
wire n_25139;
wire n_2514;
wire n_25140;
wire n_25141;
wire n_25142;
wire n_25143;
wire n_25144;
wire n_25145;
wire n_25146;
wire n_25147;
wire n_25148;
wire n_25149;
wire n_2515;
wire n_25150;
wire n_25151;
wire n_25152;
wire n_25153;
wire n_25154;
wire n_25155;
wire n_25156;
wire n_25157;
wire n_25158;
wire n_25159;
wire n_2516;
wire n_25160;
wire n_25161;
wire n_25162;
wire n_25163;
wire n_25164;
wire n_25165;
wire n_25166;
wire n_25167;
wire n_25168;
wire n_25169;
wire n_2517;
wire n_25170;
wire n_25171;
wire n_25172;
wire n_25173;
wire n_25174;
wire n_25175;
wire n_25176;
wire n_25177;
wire n_25178;
wire n_25179;
wire n_2518;
wire n_25180;
wire n_25181;
wire n_25182;
wire n_25183;
wire n_25184;
wire n_25185;
wire n_25186;
wire n_25187;
wire n_25188;
wire n_25189;
wire n_2519;
wire n_25190;
wire n_25191;
wire n_25192;
wire n_25193;
wire n_25194;
wire n_25195;
wire n_25196;
wire n_25197;
wire n_25198;
wire n_25199;
wire n_252;
wire n_2520;
wire n_25200;
wire n_25201;
wire n_25202;
wire n_25203;
wire n_25204;
wire n_25205;
wire n_25206;
wire n_25207;
wire n_25208;
wire n_25209;
wire n_2521;
wire n_25210;
wire n_25211;
wire n_25212;
wire n_25213;
wire n_25214;
wire n_25215;
wire n_25216;
wire n_25217;
wire n_25218;
wire n_25219;
wire n_2522;
wire n_25220;
wire n_25221;
wire n_25222;
wire n_25223;
wire n_25224;
wire n_25225;
wire n_25226;
wire n_25227;
wire n_25228;
wire n_25229;
wire n_2523;
wire n_25230;
wire n_25231;
wire n_25233;
wire n_25234;
wire n_25235;
wire n_25236;
wire n_25237;
wire n_25238;
wire n_25239;
wire n_2524;
wire n_25240;
wire n_25241;
wire n_25242;
wire n_25243;
wire n_25244;
wire n_25245;
wire n_25246;
wire n_25247;
wire n_25248;
wire n_25249;
wire n_2525;
wire n_25250;
wire n_25251;
wire n_25253;
wire n_25254;
wire n_25255;
wire n_25256;
wire n_25257;
wire n_25258;
wire n_25259;
wire n_2526;
wire n_25260;
wire n_25261;
wire n_25262;
wire n_25263;
wire n_25264;
wire n_25265;
wire n_25266;
wire n_25267;
wire n_25268;
wire n_25269;
wire n_2527;
wire n_25270;
wire n_25271;
wire n_25272;
wire n_25273;
wire n_25274;
wire n_25275;
wire n_25276;
wire n_25277;
wire n_25278;
wire n_25279;
wire n_2528;
wire n_25280;
wire n_25282;
wire n_25283;
wire n_25284;
wire n_25286;
wire n_25287;
wire n_25288;
wire n_25289;
wire n_2529;
wire n_25290;
wire n_25291;
wire n_25292;
wire n_25293;
wire n_25294;
wire n_25295;
wire n_25296;
wire n_25297;
wire n_25298;
wire n_25299;
wire n_253;
wire n_2530;
wire n_25300;
wire n_25301;
wire n_25302;
wire n_25303;
wire n_25304;
wire n_25305;
wire n_25306;
wire n_25307;
wire n_25308;
wire n_25309;
wire n_2531;
wire n_25310;
wire n_25311;
wire n_25312;
wire n_25313;
wire n_25314;
wire n_25315;
wire n_25316;
wire n_25317;
wire n_25318;
wire n_25319;
wire n_2532;
wire n_25320;
wire n_25321;
wire n_25322;
wire n_25323;
wire n_25324;
wire n_25325;
wire n_25326;
wire n_25327;
wire n_25328;
wire n_25329;
wire n_2533;
wire n_25330;
wire n_25331;
wire n_25332;
wire n_25333;
wire n_25334;
wire n_25335;
wire n_25336;
wire n_25337;
wire n_25338;
wire n_25339;
wire n_2534;
wire n_25340;
wire n_25341;
wire n_25342;
wire n_25343;
wire n_25344;
wire n_25345;
wire n_25346;
wire n_25347;
wire n_25348;
wire n_25349;
wire n_2535;
wire n_25351;
wire n_25353;
wire n_25355;
wire n_25356;
wire n_25357;
wire n_25358;
wire n_25359;
wire n_2536;
wire n_25360;
wire n_25361;
wire n_25362;
wire n_25363;
wire n_25364;
wire n_25365;
wire n_25366;
wire n_25367;
wire n_25368;
wire n_25369;
wire n_2537;
wire n_25370;
wire n_25371;
wire n_25372;
wire n_25374;
wire n_25375;
wire n_25376;
wire n_25377;
wire n_25378;
wire n_25379;
wire n_2538;
wire n_25380;
wire n_25381;
wire n_25382;
wire n_25383;
wire n_25384;
wire n_25385;
wire n_25386;
wire n_25387;
wire n_25388;
wire n_25389;
wire n_2539;
wire n_25390;
wire n_25391;
wire n_25392;
wire n_25393;
wire n_25394;
wire n_25395;
wire n_25396;
wire n_25397;
wire n_25398;
wire n_254;
wire n_2540;
wire n_25400;
wire n_25402;
wire n_25403;
wire n_25404;
wire n_25405;
wire n_25406;
wire n_25407;
wire n_25408;
wire n_25409;
wire n_2541;
wire n_25410;
wire n_25411;
wire n_25412;
wire n_25413;
wire n_25414;
wire n_25415;
wire n_25416;
wire n_25417;
wire n_25418;
wire n_25419;
wire n_2542;
wire n_25420;
wire n_25421;
wire n_25422;
wire n_25423;
wire n_25424;
wire n_25425;
wire n_25427;
wire n_25428;
wire n_25429;
wire n_2543;
wire n_25430;
wire n_25431;
wire n_25432;
wire n_25433;
wire n_25434;
wire n_25435;
wire n_25436;
wire n_25437;
wire n_25438;
wire n_25439;
wire n_2544;
wire n_25440;
wire n_25441;
wire n_25442;
wire n_25443;
wire n_25444;
wire n_25445;
wire n_25446;
wire n_25447;
wire n_25448;
wire n_25449;
wire n_2545;
wire n_25450;
wire n_25451;
wire n_25452;
wire n_25453;
wire n_25454;
wire n_25455;
wire n_25456;
wire n_25457;
wire n_25458;
wire n_25459;
wire n_2546;
wire n_25460;
wire n_25461;
wire n_25462;
wire n_25463;
wire n_25464;
wire n_25465;
wire n_25466;
wire n_25467;
wire n_25468;
wire n_25469;
wire n_2547;
wire n_25470;
wire n_25471;
wire n_25472;
wire n_25473;
wire n_25474;
wire n_25475;
wire n_25476;
wire n_25477;
wire n_25478;
wire n_25479;
wire n_2548;
wire n_25480;
wire n_25481;
wire n_25482;
wire n_25483;
wire n_25484;
wire n_25485;
wire n_25486;
wire n_25487;
wire n_25488;
wire n_25489;
wire n_2549;
wire n_25490;
wire n_25491;
wire n_25492;
wire n_25493;
wire n_25494;
wire n_25495;
wire n_25496;
wire n_25497;
wire n_25498;
wire n_25499;
wire n_255;
wire n_2550;
wire n_25500;
wire n_25501;
wire n_25502;
wire n_25503;
wire n_25504;
wire n_25505;
wire n_25506;
wire n_25507;
wire n_25508;
wire n_25509;
wire n_2551;
wire n_25510;
wire n_25511;
wire n_25512;
wire n_25513;
wire n_25514;
wire n_25516;
wire n_25517;
wire n_25518;
wire n_25519;
wire n_2552;
wire n_25520;
wire n_25521;
wire n_25522;
wire n_25523;
wire n_25524;
wire n_25525;
wire n_25526;
wire n_25527;
wire n_25528;
wire n_25529;
wire n_2553;
wire n_25530;
wire n_25531;
wire n_25532;
wire n_25533;
wire n_25534;
wire n_25535;
wire n_25536;
wire n_25537;
wire n_25538;
wire n_25539;
wire n_2554;
wire n_25540;
wire n_25541;
wire n_25542;
wire n_25543;
wire n_25544;
wire n_25545;
wire n_25547;
wire n_25548;
wire n_25549;
wire n_2555;
wire n_25550;
wire n_25551;
wire n_25552;
wire n_25553;
wire n_25554;
wire n_25555;
wire n_25556;
wire n_25557;
wire n_25558;
wire n_25559;
wire n_2556;
wire n_25560;
wire n_25561;
wire n_25562;
wire n_25563;
wire n_25564;
wire n_25565;
wire n_25566;
wire n_25567;
wire n_25568;
wire n_25569;
wire n_2557;
wire n_25570;
wire n_25571;
wire n_25572;
wire n_25573;
wire n_25574;
wire n_25575;
wire n_25576;
wire n_25577;
wire n_25578;
wire n_25579;
wire n_2558;
wire n_25580;
wire n_25581;
wire n_25582;
wire n_25583;
wire n_25584;
wire n_25585;
wire n_25586;
wire n_25587;
wire n_25588;
wire n_25589;
wire n_2559;
wire n_25590;
wire n_25591;
wire n_25592;
wire n_25593;
wire n_25594;
wire n_25595;
wire n_25596;
wire n_25597;
wire n_25598;
wire n_25599;
wire n_256;
wire n_2560;
wire n_25600;
wire n_25601;
wire n_25602;
wire n_25603;
wire n_25604;
wire n_25605;
wire n_25606;
wire n_25607;
wire n_25608;
wire n_25609;
wire n_2561;
wire n_25610;
wire n_25611;
wire n_25612;
wire n_25613;
wire n_25614;
wire n_25615;
wire n_25616;
wire n_25617;
wire n_25618;
wire n_25619;
wire n_2562;
wire n_25620;
wire n_25621;
wire n_25622;
wire n_25623;
wire n_25624;
wire n_25625;
wire n_25626;
wire n_25627;
wire n_25628;
wire n_25629;
wire n_2563;
wire n_25630;
wire n_25631;
wire n_25632;
wire n_25633;
wire n_25634;
wire n_25635;
wire n_25636;
wire n_25637;
wire n_25638;
wire n_25639;
wire n_2564;
wire n_25640;
wire n_25641;
wire n_25642;
wire n_25643;
wire n_25644;
wire n_25645;
wire n_25646;
wire n_25647;
wire n_25648;
wire n_25649;
wire n_2565;
wire n_25650;
wire n_25651;
wire n_25652;
wire n_25653;
wire n_25654;
wire n_25655;
wire n_25656;
wire n_25658;
wire n_25659;
wire n_2566;
wire n_25660;
wire n_25661;
wire n_25663;
wire n_25664;
wire n_25666;
wire n_25667;
wire n_25668;
wire n_25669;
wire n_2567;
wire n_25670;
wire n_25671;
wire n_25672;
wire n_25673;
wire n_25675;
wire n_25676;
wire n_25678;
wire n_25679;
wire n_2568;
wire n_25680;
wire n_25681;
wire n_25682;
wire n_25684;
wire n_25685;
wire n_25686;
wire n_25687;
wire n_25688;
wire n_25689;
wire n_2569;
wire n_25690;
wire n_25691;
wire n_25692;
wire n_25693;
wire n_25694;
wire n_25695;
wire n_25696;
wire n_25697;
wire n_25698;
wire n_25699;
wire n_257;
wire n_2570;
wire n_25700;
wire n_25701;
wire n_25702;
wire n_25703;
wire n_25704;
wire n_25705;
wire n_25706;
wire n_25707;
wire n_25708;
wire n_25709;
wire n_2571;
wire n_25710;
wire n_25711;
wire n_25712;
wire n_25713;
wire n_25714;
wire n_25715;
wire n_25716;
wire n_25717;
wire n_25718;
wire n_25719;
wire n_2572;
wire n_25720;
wire n_25721;
wire n_25722;
wire n_25723;
wire n_25724;
wire n_25725;
wire n_25726;
wire n_25727;
wire n_25728;
wire n_25729;
wire n_2573;
wire n_25730;
wire n_25731;
wire n_25732;
wire n_25733;
wire n_25734;
wire n_25735;
wire n_25736;
wire n_25737;
wire n_25738;
wire n_25739;
wire n_2574;
wire n_25740;
wire n_25741;
wire n_25743;
wire n_25744;
wire n_25745;
wire n_25746;
wire n_25747;
wire n_25748;
wire n_25749;
wire n_2575;
wire n_25750;
wire n_25751;
wire n_25752;
wire n_25753;
wire n_25754;
wire n_25755;
wire n_25756;
wire n_25757;
wire n_25758;
wire n_25759;
wire n_2576;
wire n_25760;
wire n_25761;
wire n_25762;
wire n_25763;
wire n_25764;
wire n_25765;
wire n_25766;
wire n_25767;
wire n_25768;
wire n_25769;
wire n_2577;
wire n_25770;
wire n_25771;
wire n_25772;
wire n_25773;
wire n_25774;
wire n_25775;
wire n_25776;
wire n_25777;
wire n_25778;
wire n_25779;
wire n_2578;
wire n_25780;
wire n_25781;
wire n_25782;
wire n_25783;
wire n_25784;
wire n_25785;
wire n_25786;
wire n_25787;
wire n_25788;
wire n_25789;
wire n_2579;
wire n_25790;
wire n_25791;
wire n_25792;
wire n_25793;
wire n_25794;
wire n_25795;
wire n_25796;
wire n_25797;
wire n_25798;
wire n_25799;
wire n_258;
wire n_2580;
wire n_25800;
wire n_25801;
wire n_25802;
wire n_25803;
wire n_25804;
wire n_25805;
wire n_25806;
wire n_25807;
wire n_25808;
wire n_25809;
wire n_2581;
wire n_25810;
wire n_25811;
wire n_25812;
wire n_25813;
wire n_25814;
wire n_25815;
wire n_25816;
wire n_25817;
wire n_25818;
wire n_25819;
wire n_2582;
wire n_25820;
wire n_25821;
wire n_25822;
wire n_25823;
wire n_25824;
wire n_25825;
wire n_25826;
wire n_25827;
wire n_25828;
wire n_25829;
wire n_2583;
wire n_25830;
wire n_25831;
wire n_25832;
wire n_25833;
wire n_25834;
wire n_25835;
wire n_25836;
wire n_25837;
wire n_25838;
wire n_25839;
wire n_2584;
wire n_25840;
wire n_25841;
wire n_25842;
wire n_25843;
wire n_25844;
wire n_25845;
wire n_25846;
wire n_25847;
wire n_25848;
wire n_25849;
wire n_2585;
wire n_25850;
wire n_25851;
wire n_25852;
wire n_25853;
wire n_25854;
wire n_25855;
wire n_25856;
wire n_25857;
wire n_25858;
wire n_25859;
wire n_2586;
wire n_25860;
wire n_25861;
wire n_25862;
wire n_25863;
wire n_25864;
wire n_25865;
wire n_25866;
wire n_25867;
wire n_25868;
wire n_25869;
wire n_2587;
wire n_25870;
wire n_25871;
wire n_25872;
wire n_25873;
wire n_25874;
wire n_25875;
wire n_25876;
wire n_25878;
wire n_25879;
wire n_2588;
wire n_25880;
wire n_25881;
wire n_25883;
wire n_25884;
wire n_25886;
wire n_25887;
wire n_25888;
wire n_25889;
wire n_2589;
wire n_25890;
wire n_25891;
wire n_25892;
wire n_25893;
wire n_25894;
wire n_25896;
wire n_25897;
wire n_25898;
wire n_25899;
wire n_259;
wire n_2590;
wire n_25900;
wire n_25902;
wire n_25904;
wire n_25905;
wire n_25906;
wire n_25907;
wire n_25908;
wire n_25909;
wire n_2591;
wire n_25910;
wire n_25911;
wire n_25912;
wire n_25913;
wire n_25914;
wire n_25915;
wire n_25916;
wire n_25917;
wire n_25918;
wire n_25919;
wire n_2592;
wire n_25920;
wire n_25921;
wire n_25922;
wire n_25923;
wire n_25924;
wire n_25925;
wire n_25926;
wire n_25927;
wire n_25928;
wire n_25929;
wire n_2593;
wire n_25930;
wire n_25931;
wire n_25932;
wire n_25933;
wire n_25934;
wire n_25935;
wire n_25936;
wire n_25937;
wire n_25938;
wire n_25939;
wire n_2594;
wire n_25940;
wire n_25941;
wire n_25942;
wire n_25943;
wire n_25944;
wire n_25945;
wire n_25946;
wire n_25947;
wire n_25948;
wire n_25949;
wire n_2595;
wire n_25950;
wire n_25951;
wire n_25952;
wire n_25953;
wire n_25954;
wire n_25955;
wire n_25956;
wire n_25957;
wire n_25958;
wire n_25959;
wire n_2596;
wire n_25960;
wire n_25961;
wire n_25962;
wire n_25963;
wire n_25964;
wire n_25965;
wire n_25966;
wire n_25967;
wire n_25968;
wire n_25969;
wire n_2597;
wire n_25970;
wire n_25971;
wire n_25972;
wire n_25973;
wire n_25974;
wire n_25975;
wire n_25976;
wire n_25977;
wire n_25978;
wire n_25979;
wire n_2598;
wire n_25980;
wire n_25981;
wire n_25982;
wire n_25983;
wire n_25984;
wire n_25985;
wire n_25986;
wire n_25987;
wire n_25988;
wire n_25989;
wire n_2599;
wire n_25990;
wire n_25991;
wire n_25992;
wire n_25993;
wire n_25994;
wire n_25995;
wire n_25996;
wire n_25997;
wire n_25998;
wire n_25999;
wire n_26;
wire n_260;
wire n_2600;
wire n_26000;
wire n_26001;
wire n_26002;
wire n_26003;
wire n_26004;
wire n_26005;
wire n_26006;
wire n_26007;
wire n_26008;
wire n_26009;
wire n_2601;
wire n_26010;
wire n_26011;
wire n_26012;
wire n_26013;
wire n_26014;
wire n_26016;
wire n_26017;
wire n_26018;
wire n_26019;
wire n_2602;
wire n_26020;
wire n_26021;
wire n_26022;
wire n_26023;
wire n_26024;
wire n_26025;
wire n_26026;
wire n_26027;
wire n_26028;
wire n_26029;
wire n_2603;
wire n_26030;
wire n_26031;
wire n_26032;
wire n_26033;
wire n_26034;
wire n_26035;
wire n_26036;
wire n_26037;
wire n_26038;
wire n_26039;
wire n_2604;
wire n_26040;
wire n_26041;
wire n_26042;
wire n_26043;
wire n_26044;
wire n_26045;
wire n_26046;
wire n_26047;
wire n_26048;
wire n_26049;
wire n_2605;
wire n_26050;
wire n_26051;
wire n_26052;
wire n_26053;
wire n_26054;
wire n_26055;
wire n_26056;
wire n_26057;
wire n_26058;
wire n_26059;
wire n_2606;
wire n_26060;
wire n_26061;
wire n_26062;
wire n_26063;
wire n_26064;
wire n_26065;
wire n_26066;
wire n_26067;
wire n_26068;
wire n_26069;
wire n_2607;
wire n_26070;
wire n_26071;
wire n_26072;
wire n_26073;
wire n_26074;
wire n_26075;
wire n_26076;
wire n_26077;
wire n_26078;
wire n_26079;
wire n_2608;
wire n_26080;
wire n_26081;
wire n_26082;
wire n_26083;
wire n_26084;
wire n_26085;
wire n_26086;
wire n_26087;
wire n_26088;
wire n_26089;
wire n_2609;
wire n_26090;
wire n_26091;
wire n_26092;
wire n_26093;
wire n_26094;
wire n_26095;
wire n_26096;
wire n_26097;
wire n_26098;
wire n_26099;
wire n_261;
wire n_2610;
wire n_26100;
wire n_26101;
wire n_26102;
wire n_26103;
wire n_26104;
wire n_26105;
wire n_26106;
wire n_26107;
wire n_26108;
wire n_26109;
wire n_2611;
wire n_26110;
wire n_26111;
wire n_26112;
wire n_26113;
wire n_26114;
wire n_26115;
wire n_26116;
wire n_26117;
wire n_26118;
wire n_26119;
wire n_2612;
wire n_26121;
wire n_26122;
wire n_26123;
wire n_26124;
wire n_26125;
wire n_26126;
wire n_26127;
wire n_26128;
wire n_26129;
wire n_2613;
wire n_26130;
wire n_26131;
wire n_26132;
wire n_26133;
wire n_26134;
wire n_26135;
wire n_26136;
wire n_26137;
wire n_26138;
wire n_26139;
wire n_2614;
wire n_26140;
wire n_26141;
wire n_26142;
wire n_26143;
wire n_26144;
wire n_26145;
wire n_26146;
wire n_26147;
wire n_26148;
wire n_26149;
wire n_2615;
wire n_26150;
wire n_26151;
wire n_26152;
wire n_26153;
wire n_26154;
wire n_26155;
wire n_26156;
wire n_26157;
wire n_26158;
wire n_26159;
wire n_2616;
wire n_26160;
wire n_26161;
wire n_26162;
wire n_26163;
wire n_26164;
wire n_26165;
wire n_26166;
wire n_26167;
wire n_26168;
wire n_26169;
wire n_2617;
wire n_26170;
wire n_26171;
wire n_26172;
wire n_26173;
wire n_26174;
wire n_26175;
wire n_26176;
wire n_26177;
wire n_26178;
wire n_26179;
wire n_2618;
wire n_26180;
wire n_26181;
wire n_26182;
wire n_26183;
wire n_26184;
wire n_26185;
wire n_26186;
wire n_26187;
wire n_26188;
wire n_26189;
wire n_2619;
wire n_26190;
wire n_26191;
wire n_26192;
wire n_26193;
wire n_26194;
wire n_26195;
wire n_26196;
wire n_26197;
wire n_26198;
wire n_26199;
wire n_262;
wire n_2620;
wire n_26200;
wire n_26201;
wire n_26202;
wire n_26203;
wire n_26204;
wire n_26205;
wire n_26206;
wire n_26207;
wire n_26208;
wire n_26209;
wire n_2621;
wire n_26210;
wire n_26211;
wire n_26212;
wire n_26213;
wire n_26214;
wire n_26215;
wire n_26216;
wire n_26217;
wire n_26218;
wire n_26219;
wire n_2622;
wire n_26220;
wire n_26221;
wire n_26222;
wire n_26223;
wire n_26224;
wire n_26225;
wire n_26226;
wire n_26227;
wire n_26228;
wire n_26229;
wire n_2623;
wire n_26231;
wire n_26233;
wire n_26234;
wire n_26235;
wire n_26237;
wire n_26238;
wire n_26239;
wire n_2624;
wire n_26240;
wire n_26241;
wire n_26242;
wire n_26243;
wire n_26244;
wire n_26245;
wire n_26246;
wire n_26247;
wire n_26248;
wire n_26249;
wire n_2625;
wire n_26250;
wire n_26251;
wire n_26252;
wire n_26253;
wire n_26254;
wire n_26255;
wire n_26256;
wire n_26257;
wire n_26258;
wire n_26259;
wire n_2626;
wire n_26260;
wire n_26261;
wire n_26262;
wire n_26263;
wire n_26264;
wire n_26265;
wire n_26266;
wire n_26267;
wire n_26268;
wire n_26269;
wire n_2627;
wire n_26270;
wire n_26271;
wire n_26272;
wire n_26273;
wire n_26274;
wire n_26275;
wire n_26276;
wire n_26277;
wire n_26278;
wire n_26279;
wire n_2628;
wire n_26280;
wire n_26281;
wire n_26282;
wire n_26283;
wire n_26284;
wire n_26285;
wire n_26286;
wire n_26287;
wire n_26288;
wire n_26289;
wire n_2629;
wire n_26290;
wire n_26291;
wire n_26292;
wire n_26293;
wire n_26294;
wire n_26295;
wire n_26296;
wire n_26297;
wire n_26298;
wire n_26299;
wire n_263;
wire n_2630;
wire n_26300;
wire n_26301;
wire n_26302;
wire n_26303;
wire n_26304;
wire n_26306;
wire n_26307;
wire n_26308;
wire n_26309;
wire n_2631;
wire n_26310;
wire n_26311;
wire n_26312;
wire n_26313;
wire n_26314;
wire n_26315;
wire n_26316;
wire n_26317;
wire n_26318;
wire n_26319;
wire n_2632;
wire n_26320;
wire n_26321;
wire n_26322;
wire n_26323;
wire n_26324;
wire n_26325;
wire n_26326;
wire n_26327;
wire n_26328;
wire n_26329;
wire n_2633;
wire n_26330;
wire n_26331;
wire n_26332;
wire n_26333;
wire n_26334;
wire n_26335;
wire n_26336;
wire n_26337;
wire n_26338;
wire n_26339;
wire n_2634;
wire n_26340;
wire n_26341;
wire n_26342;
wire n_26343;
wire n_26344;
wire n_26345;
wire n_26346;
wire n_26347;
wire n_26348;
wire n_26349;
wire n_2635;
wire n_26350;
wire n_26351;
wire n_26352;
wire n_26353;
wire n_26354;
wire n_26355;
wire n_26356;
wire n_26357;
wire n_26358;
wire n_26359;
wire n_2636;
wire n_26360;
wire n_26361;
wire n_26362;
wire n_26363;
wire n_26364;
wire n_26365;
wire n_26366;
wire n_26367;
wire n_26368;
wire n_26369;
wire n_2637;
wire n_26370;
wire n_26371;
wire n_26372;
wire n_26373;
wire n_26374;
wire n_26375;
wire n_26376;
wire n_26377;
wire n_26378;
wire n_26379;
wire n_2638;
wire n_26380;
wire n_26381;
wire n_26382;
wire n_26383;
wire n_26384;
wire n_26385;
wire n_26386;
wire n_26387;
wire n_26388;
wire n_26389;
wire n_2639;
wire n_26390;
wire n_26391;
wire n_26392;
wire n_26393;
wire n_26394;
wire n_26395;
wire n_26396;
wire n_26397;
wire n_26398;
wire n_26399;
wire n_264;
wire n_2640;
wire n_26400;
wire n_26401;
wire n_26402;
wire n_26403;
wire n_26404;
wire n_26405;
wire n_26406;
wire n_26407;
wire n_26408;
wire n_26409;
wire n_2641;
wire n_26410;
wire n_26411;
wire n_26412;
wire n_26413;
wire n_26414;
wire n_26415;
wire n_26416;
wire n_26417;
wire n_26418;
wire n_26419;
wire n_2642;
wire n_26420;
wire n_26421;
wire n_26422;
wire n_26423;
wire n_26424;
wire n_26425;
wire n_26426;
wire n_26427;
wire n_26428;
wire n_26429;
wire n_2643;
wire n_26430;
wire n_26431;
wire n_26432;
wire n_26433;
wire n_26434;
wire n_26435;
wire n_26436;
wire n_26437;
wire n_26438;
wire n_26439;
wire n_2644;
wire n_26440;
wire n_26441;
wire n_26442;
wire n_26443;
wire n_26444;
wire n_26445;
wire n_26446;
wire n_26447;
wire n_26448;
wire n_26449;
wire n_2645;
wire n_26450;
wire n_26451;
wire n_26452;
wire n_26453;
wire n_26454;
wire n_26455;
wire n_26456;
wire n_26457;
wire n_26458;
wire n_26459;
wire n_2646;
wire n_26460;
wire n_26461;
wire n_26462;
wire n_26463;
wire n_26464;
wire n_26465;
wire n_26466;
wire n_26467;
wire n_26468;
wire n_26469;
wire n_2647;
wire n_26470;
wire n_26471;
wire n_26472;
wire n_26473;
wire n_26474;
wire n_26475;
wire n_26476;
wire n_26477;
wire n_26478;
wire n_26479;
wire n_26480;
wire n_26481;
wire n_26482;
wire n_26483;
wire n_26484;
wire n_26485;
wire n_26486;
wire n_26487;
wire n_26488;
wire n_26489;
wire n_2649;
wire n_26490;
wire n_26491;
wire n_26492;
wire n_26493;
wire n_26494;
wire n_26495;
wire n_26496;
wire n_26497;
wire n_26498;
wire n_26499;
wire n_265;
wire n_2650;
wire n_26500;
wire n_26501;
wire n_26502;
wire n_26503;
wire n_26504;
wire n_26505;
wire n_26506;
wire n_26507;
wire n_26508;
wire n_26509;
wire n_2651;
wire n_26510;
wire n_26511;
wire n_26512;
wire n_26513;
wire n_26514;
wire n_26515;
wire n_26516;
wire n_26517;
wire n_26518;
wire n_26519;
wire n_2652;
wire n_26520;
wire n_26522;
wire n_26523;
wire n_26524;
wire n_26526;
wire n_26528;
wire n_26529;
wire n_2653;
wire n_26530;
wire n_26532;
wire n_26533;
wire n_26534;
wire n_26535;
wire n_26536;
wire n_26537;
wire n_26538;
wire n_26539;
wire n_2654;
wire n_26540;
wire n_26541;
wire n_26542;
wire n_26543;
wire n_26544;
wire n_26545;
wire n_26546;
wire n_26547;
wire n_26548;
wire n_26549;
wire n_2655;
wire n_26550;
wire n_26551;
wire n_26552;
wire n_26553;
wire n_26554;
wire n_26555;
wire n_26556;
wire n_26557;
wire n_26558;
wire n_26559;
wire n_2656;
wire n_26560;
wire n_26561;
wire n_26562;
wire n_26563;
wire n_26564;
wire n_26566;
wire n_26567;
wire n_26568;
wire n_26569;
wire n_2657;
wire n_26570;
wire n_26571;
wire n_26572;
wire n_26573;
wire n_26574;
wire n_26575;
wire n_26576;
wire n_26577;
wire n_26578;
wire n_26579;
wire n_2658;
wire n_26580;
wire n_26581;
wire n_26582;
wire n_26583;
wire n_26584;
wire n_26585;
wire n_26586;
wire n_26587;
wire n_26588;
wire n_26589;
wire n_2659;
wire n_26590;
wire n_26591;
wire n_26592;
wire n_26593;
wire n_26594;
wire n_26595;
wire n_26596;
wire n_26597;
wire n_26598;
wire n_26599;
wire n_266;
wire n_2660;
wire n_26600;
wire n_26601;
wire n_26602;
wire n_26603;
wire n_26604;
wire n_26605;
wire n_26606;
wire n_26607;
wire n_26608;
wire n_26609;
wire n_2661;
wire n_26610;
wire n_26611;
wire n_26612;
wire n_26613;
wire n_26614;
wire n_26615;
wire n_26616;
wire n_26617;
wire n_26618;
wire n_26619;
wire n_2662;
wire n_26620;
wire n_26621;
wire n_26622;
wire n_26623;
wire n_26624;
wire n_26625;
wire n_26626;
wire n_26627;
wire n_26628;
wire n_26629;
wire n_2663;
wire n_26630;
wire n_26631;
wire n_26632;
wire n_26633;
wire n_26634;
wire n_26635;
wire n_26636;
wire n_26637;
wire n_26638;
wire n_26639;
wire n_2664;
wire n_26640;
wire n_26641;
wire n_26642;
wire n_26643;
wire n_26644;
wire n_26645;
wire n_26646;
wire n_26647;
wire n_26648;
wire n_26649;
wire n_2665;
wire n_26650;
wire n_26651;
wire n_26652;
wire n_26653;
wire n_26654;
wire n_26655;
wire n_26656;
wire n_26657;
wire n_26658;
wire n_26659;
wire n_2666;
wire n_26660;
wire n_26661;
wire n_26662;
wire n_26663;
wire n_26664;
wire n_26665;
wire n_26666;
wire n_26667;
wire n_26668;
wire n_26669;
wire n_26670;
wire n_26671;
wire n_26672;
wire n_26673;
wire n_26674;
wire n_26675;
wire n_26676;
wire n_26677;
wire n_26678;
wire n_26679;
wire n_2668;
wire n_26680;
wire n_26681;
wire n_26682;
wire n_26683;
wire n_26684;
wire n_26685;
wire n_26686;
wire n_26687;
wire n_26688;
wire n_26689;
wire n_2669;
wire n_26690;
wire n_26691;
wire n_26692;
wire n_26693;
wire n_26694;
wire n_26695;
wire n_26696;
wire n_26697;
wire n_26698;
wire n_26699;
wire n_267;
wire n_26700;
wire n_26701;
wire n_26702;
wire n_26703;
wire n_26704;
wire n_26705;
wire n_26706;
wire n_26707;
wire n_26708;
wire n_26709;
wire n_2671;
wire n_26710;
wire n_26711;
wire n_26712;
wire n_26713;
wire n_26714;
wire n_26715;
wire n_26716;
wire n_26717;
wire n_26718;
wire n_26719;
wire n_2672;
wire n_26720;
wire n_26721;
wire n_26722;
wire n_26723;
wire n_26724;
wire n_26725;
wire n_26726;
wire n_26727;
wire n_26728;
wire n_26729;
wire n_2673;
wire n_26730;
wire n_26731;
wire n_26732;
wire n_26733;
wire n_26734;
wire n_26735;
wire n_26736;
wire n_26737;
wire n_26738;
wire n_26739;
wire n_2674;
wire n_26740;
wire n_26741;
wire n_26742;
wire n_26743;
wire n_26744;
wire n_26745;
wire n_26746;
wire n_26747;
wire n_26748;
wire n_26749;
wire n_2675;
wire n_26750;
wire n_26751;
wire n_26752;
wire n_26753;
wire n_26754;
wire n_26755;
wire n_26756;
wire n_26757;
wire n_26758;
wire n_26759;
wire n_2676;
wire n_26760;
wire n_26761;
wire n_26762;
wire n_26764;
wire n_26765;
wire n_26766;
wire n_26767;
wire n_26768;
wire n_2677;
wire n_26771;
wire n_26772;
wire n_26774;
wire n_26775;
wire n_26776;
wire n_26777;
wire n_26778;
wire n_26779;
wire n_2678;
wire n_26780;
wire n_26781;
wire n_26783;
wire n_26784;
wire n_26785;
wire n_26786;
wire n_26787;
wire n_26788;
wire n_26789;
wire n_2679;
wire n_26790;
wire n_26791;
wire n_26792;
wire n_26793;
wire n_26794;
wire n_26795;
wire n_26796;
wire n_26797;
wire n_26798;
wire n_26799;
wire n_268;
wire n_2680;
wire n_26800;
wire n_26801;
wire n_26803;
wire n_26804;
wire n_26806;
wire n_26807;
wire n_26808;
wire n_26809;
wire n_2681;
wire n_26810;
wire n_26811;
wire n_26812;
wire n_26814;
wire n_26815;
wire n_26816;
wire n_26817;
wire n_26818;
wire n_26819;
wire n_2682;
wire n_26820;
wire n_26821;
wire n_26822;
wire n_26823;
wire n_26824;
wire n_26825;
wire n_26826;
wire n_26827;
wire n_26828;
wire n_26829;
wire n_26830;
wire n_26831;
wire n_26832;
wire n_26833;
wire n_26834;
wire n_26835;
wire n_26836;
wire n_26837;
wire n_26838;
wire n_26839;
wire n_26840;
wire n_26841;
wire n_26842;
wire n_26843;
wire n_26844;
wire n_26845;
wire n_26846;
wire n_26847;
wire n_26848;
wire n_26849;
wire n_2685;
wire n_26850;
wire n_26851;
wire n_26852;
wire n_26853;
wire n_26854;
wire n_26855;
wire n_26856;
wire n_26857;
wire n_26858;
wire n_26859;
wire n_2686;
wire n_26860;
wire n_26861;
wire n_26862;
wire n_26863;
wire n_26864;
wire n_26865;
wire n_26866;
wire n_26867;
wire n_26868;
wire n_26869;
wire n_2687;
wire n_26870;
wire n_26871;
wire n_26872;
wire n_26873;
wire n_26874;
wire n_26875;
wire n_26876;
wire n_26877;
wire n_26878;
wire n_26879;
wire n_26880;
wire n_26881;
wire n_26882;
wire n_26883;
wire n_26884;
wire n_26885;
wire n_26886;
wire n_26887;
wire n_26888;
wire n_26889;
wire n_2689;
wire n_26890;
wire n_26891;
wire n_26892;
wire n_26893;
wire n_26894;
wire n_26895;
wire n_26896;
wire n_26897;
wire n_26898;
wire n_26899;
wire n_269;
wire n_2690;
wire n_26900;
wire n_26901;
wire n_26902;
wire n_26903;
wire n_26904;
wire n_26905;
wire n_26906;
wire n_26907;
wire n_26908;
wire n_26909;
wire n_2691;
wire n_26910;
wire n_26911;
wire n_26912;
wire n_26913;
wire n_26914;
wire n_26915;
wire n_26916;
wire n_26917;
wire n_26918;
wire n_26919;
wire n_2692;
wire n_26920;
wire n_26921;
wire n_26922;
wire n_26923;
wire n_26924;
wire n_26925;
wire n_26926;
wire n_26927;
wire n_26928;
wire n_26929;
wire n_2693;
wire n_26930;
wire n_26931;
wire n_26932;
wire n_26933;
wire n_26934;
wire n_26935;
wire n_26936;
wire n_26937;
wire n_26938;
wire n_26939;
wire n_2694;
wire n_26940;
wire n_26941;
wire n_26942;
wire n_26943;
wire n_26945;
wire n_26946;
wire n_26947;
wire n_26948;
wire n_26949;
wire n_2695;
wire n_26950;
wire n_26951;
wire n_26952;
wire n_26953;
wire n_26954;
wire n_26955;
wire n_26956;
wire n_26957;
wire n_26958;
wire n_26959;
wire n_2696;
wire n_26960;
wire n_26961;
wire n_26962;
wire n_26963;
wire n_26964;
wire n_26965;
wire n_26966;
wire n_26967;
wire n_26968;
wire n_26969;
wire n_2697;
wire n_26970;
wire n_26971;
wire n_26972;
wire n_26973;
wire n_26974;
wire n_26975;
wire n_26976;
wire n_26977;
wire n_26978;
wire n_26979;
wire n_2698;
wire n_26980;
wire n_26981;
wire n_26982;
wire n_26983;
wire n_26984;
wire n_26985;
wire n_26986;
wire n_26987;
wire n_26988;
wire n_26989;
wire n_2699;
wire n_26990;
wire n_26991;
wire n_26992;
wire n_26993;
wire n_26994;
wire n_26995;
wire n_26996;
wire n_26997;
wire n_26998;
wire n_26999;
wire n_27;
wire n_270;
wire n_2700;
wire n_27000;
wire n_27001;
wire n_27002;
wire n_27003;
wire n_27004;
wire n_27005;
wire n_27006;
wire n_27007;
wire n_27008;
wire n_27009;
wire n_27011;
wire n_27012;
wire n_27013;
wire n_27014;
wire n_27015;
wire n_27016;
wire n_27017;
wire n_27018;
wire n_27019;
wire n_2702;
wire n_27020;
wire n_27021;
wire n_27022;
wire n_27023;
wire n_27024;
wire n_27025;
wire n_27026;
wire n_27028;
wire n_27029;
wire n_2703;
wire n_27030;
wire n_27031;
wire n_27032;
wire n_27033;
wire n_27034;
wire n_27035;
wire n_27036;
wire n_27037;
wire n_27038;
wire n_27039;
wire n_2704;
wire n_27040;
wire n_27041;
wire n_27042;
wire n_27043;
wire n_27044;
wire n_27045;
wire n_27046;
wire n_27047;
wire n_27048;
wire n_2705;
wire n_27050;
wire n_27051;
wire n_27052;
wire n_27053;
wire n_27054;
wire n_27055;
wire n_27056;
wire n_27057;
wire n_27058;
wire n_27059;
wire n_2706;
wire n_27060;
wire n_27061;
wire n_27062;
wire n_27063;
wire n_27064;
wire n_27065;
wire n_27066;
wire n_27067;
wire n_27068;
wire n_27069;
wire n_2707;
wire n_27070;
wire n_27071;
wire n_27072;
wire n_27074;
wire n_27075;
wire n_27076;
wire n_27077;
wire n_27078;
wire n_27079;
wire n_2708;
wire n_27080;
wire n_27081;
wire n_27082;
wire n_27083;
wire n_27084;
wire n_27085;
wire n_27086;
wire n_27087;
wire n_27088;
wire n_27089;
wire n_2709;
wire n_27090;
wire n_27091;
wire n_27092;
wire n_27093;
wire n_27094;
wire n_27095;
wire n_27096;
wire n_27097;
wire n_27098;
wire n_27099;
wire n_271;
wire n_2710;
wire n_27100;
wire n_27101;
wire n_27102;
wire n_27103;
wire n_27104;
wire n_27105;
wire n_27106;
wire n_27107;
wire n_27108;
wire n_27109;
wire n_2711;
wire n_27110;
wire n_27111;
wire n_27112;
wire n_27113;
wire n_27114;
wire n_27115;
wire n_27116;
wire n_27117;
wire n_27118;
wire n_27119;
wire n_2712;
wire n_27120;
wire n_27121;
wire n_27122;
wire n_27123;
wire n_27124;
wire n_27125;
wire n_27126;
wire n_27127;
wire n_27128;
wire n_27129;
wire n_2713;
wire n_27130;
wire n_27131;
wire n_27132;
wire n_27133;
wire n_27134;
wire n_27135;
wire n_27136;
wire n_27137;
wire n_27138;
wire n_27139;
wire n_2714;
wire n_27140;
wire n_27141;
wire n_27142;
wire n_27143;
wire n_27144;
wire n_27145;
wire n_27146;
wire n_27147;
wire n_27148;
wire n_27149;
wire n_2715;
wire n_27150;
wire n_27151;
wire n_27152;
wire n_27153;
wire n_27154;
wire n_27155;
wire n_27156;
wire n_27157;
wire n_27158;
wire n_27159;
wire n_2716;
wire n_27160;
wire n_27161;
wire n_27162;
wire n_27163;
wire n_27164;
wire n_27165;
wire n_27166;
wire n_27167;
wire n_27169;
wire n_2717;
wire n_27170;
wire n_27171;
wire n_27172;
wire n_27173;
wire n_27174;
wire n_27175;
wire n_27176;
wire n_27177;
wire n_27178;
wire n_27179;
wire n_2718;
wire n_27180;
wire n_27181;
wire n_27182;
wire n_27183;
wire n_27184;
wire n_27185;
wire n_27186;
wire n_27187;
wire n_27188;
wire n_27189;
wire n_2719;
wire n_27190;
wire n_27191;
wire n_27192;
wire n_27193;
wire n_27194;
wire n_27195;
wire n_27196;
wire n_27197;
wire n_27198;
wire n_27199;
wire n_272;
wire n_2720;
wire n_27200;
wire n_27201;
wire n_27202;
wire n_27203;
wire n_27204;
wire n_27205;
wire n_27206;
wire n_27208;
wire n_27209;
wire n_2721;
wire n_27210;
wire n_27211;
wire n_27212;
wire n_27213;
wire n_27214;
wire n_27215;
wire n_27216;
wire n_27217;
wire n_27218;
wire n_27219;
wire n_2722;
wire n_27220;
wire n_27221;
wire n_27222;
wire n_27223;
wire n_27224;
wire n_27225;
wire n_27226;
wire n_27227;
wire n_27228;
wire n_27229;
wire n_2723;
wire n_27230;
wire n_27231;
wire n_27233;
wire n_27234;
wire n_27235;
wire n_27236;
wire n_27237;
wire n_27238;
wire n_27239;
wire n_2724;
wire n_27240;
wire n_27241;
wire n_27242;
wire n_27243;
wire n_27244;
wire n_27245;
wire n_27246;
wire n_27247;
wire n_27248;
wire n_27249;
wire n_2725;
wire n_27250;
wire n_27252;
wire n_27253;
wire n_27254;
wire n_27255;
wire n_27256;
wire n_27257;
wire n_27258;
wire n_27259;
wire n_2726;
wire n_27260;
wire n_27261;
wire n_27262;
wire n_27263;
wire n_27264;
wire n_27265;
wire n_27267;
wire n_27268;
wire n_27269;
wire n_2727;
wire n_27270;
wire n_27271;
wire n_27272;
wire n_27273;
wire n_27274;
wire n_27275;
wire n_27276;
wire n_27277;
wire n_27278;
wire n_27279;
wire n_2728;
wire n_27280;
wire n_27281;
wire n_27282;
wire n_27283;
wire n_27284;
wire n_27285;
wire n_27286;
wire n_27287;
wire n_27288;
wire n_27289;
wire n_2729;
wire n_27290;
wire n_27291;
wire n_27292;
wire n_27293;
wire n_27294;
wire n_27295;
wire n_27296;
wire n_27297;
wire n_27298;
wire n_27299;
wire n_273;
wire n_2730;
wire n_27300;
wire n_27301;
wire n_27302;
wire n_27303;
wire n_27304;
wire n_27305;
wire n_27306;
wire n_27307;
wire n_27308;
wire n_27309;
wire n_2731;
wire n_27310;
wire n_27311;
wire n_27312;
wire n_27313;
wire n_27314;
wire n_27315;
wire n_27316;
wire n_27317;
wire n_27318;
wire n_27319;
wire n_2732;
wire n_27320;
wire n_27321;
wire n_27322;
wire n_27323;
wire n_27324;
wire n_27325;
wire n_27326;
wire n_27327;
wire n_27328;
wire n_27329;
wire n_2733;
wire n_27330;
wire n_27331;
wire n_27332;
wire n_27333;
wire n_27334;
wire n_27335;
wire n_27336;
wire n_27337;
wire n_27338;
wire n_27339;
wire n_2734;
wire n_27340;
wire n_27341;
wire n_27343;
wire n_27344;
wire n_27346;
wire n_27348;
wire n_27349;
wire n_2735;
wire n_27350;
wire n_27351;
wire n_27352;
wire n_27353;
wire n_27354;
wire n_27355;
wire n_27356;
wire n_27357;
wire n_27358;
wire n_27359;
wire n_2736;
wire n_27360;
wire n_27361;
wire n_27362;
wire n_27363;
wire n_27364;
wire n_27366;
wire n_27367;
wire n_27368;
wire n_27369;
wire n_2737;
wire n_27370;
wire n_27372;
wire n_27373;
wire n_27374;
wire n_27375;
wire n_27376;
wire n_27377;
wire n_27379;
wire n_2738;
wire n_27380;
wire n_27381;
wire n_27382;
wire n_27383;
wire n_27384;
wire n_27385;
wire n_27386;
wire n_27387;
wire n_27388;
wire n_27389;
wire n_2739;
wire n_27390;
wire n_27391;
wire n_27392;
wire n_27393;
wire n_27394;
wire n_27395;
wire n_27396;
wire n_27397;
wire n_27398;
wire n_27399;
wire n_274;
wire n_2740;
wire n_27400;
wire n_27401;
wire n_27402;
wire n_27403;
wire n_27404;
wire n_27405;
wire n_27406;
wire n_27407;
wire n_27408;
wire n_27409;
wire n_2741;
wire n_27410;
wire n_27411;
wire n_27412;
wire n_27413;
wire n_27414;
wire n_27415;
wire n_27416;
wire n_27417;
wire n_27418;
wire n_27419;
wire n_2742;
wire n_27420;
wire n_27421;
wire n_27422;
wire n_27423;
wire n_27424;
wire n_27425;
wire n_27426;
wire n_27427;
wire n_27428;
wire n_27429;
wire n_2743;
wire n_27430;
wire n_27431;
wire n_27432;
wire n_27433;
wire n_27434;
wire n_27435;
wire n_27436;
wire n_27437;
wire n_27438;
wire n_27439;
wire n_2744;
wire n_27440;
wire n_27441;
wire n_27442;
wire n_27443;
wire n_27444;
wire n_27445;
wire n_27446;
wire n_27447;
wire n_27448;
wire n_27449;
wire n_2745;
wire n_27450;
wire n_27451;
wire n_27452;
wire n_27453;
wire n_27454;
wire n_27455;
wire n_27456;
wire n_27457;
wire n_27458;
wire n_27459;
wire n_2746;
wire n_27460;
wire n_27461;
wire n_27462;
wire n_27463;
wire n_27464;
wire n_27465;
wire n_27466;
wire n_27467;
wire n_27468;
wire n_27469;
wire n_2747;
wire n_27470;
wire n_27471;
wire n_27472;
wire n_27473;
wire n_27474;
wire n_27475;
wire n_27476;
wire n_27477;
wire n_27478;
wire n_27479;
wire n_2748;
wire n_27480;
wire n_27481;
wire n_27482;
wire n_27483;
wire n_27484;
wire n_27485;
wire n_27486;
wire n_27487;
wire n_27488;
wire n_27489;
wire n_2749;
wire n_27490;
wire n_27491;
wire n_27492;
wire n_27493;
wire n_27494;
wire n_27495;
wire n_27496;
wire n_27497;
wire n_27498;
wire n_27499;
wire n_275;
wire n_2750;
wire n_27500;
wire n_27501;
wire n_27502;
wire n_27503;
wire n_27504;
wire n_27505;
wire n_27506;
wire n_27507;
wire n_27508;
wire n_27509;
wire n_2751;
wire n_27510;
wire n_27511;
wire n_27512;
wire n_27513;
wire n_27514;
wire n_27515;
wire n_27516;
wire n_27517;
wire n_27518;
wire n_27519;
wire n_2752;
wire n_27520;
wire n_27521;
wire n_27522;
wire n_27523;
wire n_27524;
wire n_27525;
wire n_27526;
wire n_27527;
wire n_27528;
wire n_27529;
wire n_2753;
wire n_27530;
wire n_27531;
wire n_27532;
wire n_27533;
wire n_27534;
wire n_27535;
wire n_27536;
wire n_27537;
wire n_27538;
wire n_27539;
wire n_2754;
wire n_27540;
wire n_27541;
wire n_27542;
wire n_27543;
wire n_27544;
wire n_27546;
wire n_27547;
wire n_27548;
wire n_27549;
wire n_2755;
wire n_27550;
wire n_27551;
wire n_27552;
wire n_27553;
wire n_27554;
wire n_27556;
wire n_27557;
wire n_27559;
wire n_2756;
wire n_27560;
wire n_27561;
wire n_27562;
wire n_27563;
wire n_27564;
wire n_27566;
wire n_27567;
wire n_27568;
wire n_27569;
wire n_2757;
wire n_27570;
wire n_27571;
wire n_27572;
wire n_27573;
wire n_27574;
wire n_27575;
wire n_27576;
wire n_27577;
wire n_27578;
wire n_27579;
wire n_27580;
wire n_27581;
wire n_27582;
wire n_27583;
wire n_27584;
wire n_27585;
wire n_27586;
wire n_27587;
wire n_27588;
wire n_27589;
wire n_2759;
wire n_27590;
wire n_27591;
wire n_27592;
wire n_27593;
wire n_27594;
wire n_27595;
wire n_27596;
wire n_27597;
wire n_27598;
wire n_27599;
wire n_276;
wire n_2760;
wire n_27600;
wire n_27601;
wire n_27602;
wire n_27603;
wire n_27604;
wire n_27605;
wire n_27606;
wire n_27607;
wire n_27609;
wire n_2761;
wire n_27610;
wire n_27611;
wire n_27612;
wire n_27614;
wire n_27615;
wire n_27616;
wire n_27617;
wire n_27618;
wire n_27619;
wire n_2762;
wire n_27620;
wire n_27621;
wire n_27622;
wire n_27623;
wire n_27624;
wire n_27625;
wire n_27626;
wire n_27627;
wire n_27628;
wire n_27629;
wire n_2763;
wire n_27630;
wire n_27631;
wire n_27632;
wire n_27633;
wire n_27634;
wire n_27635;
wire n_27636;
wire n_27637;
wire n_27638;
wire n_27639;
wire n_27640;
wire n_27641;
wire n_27642;
wire n_27643;
wire n_27644;
wire n_27645;
wire n_27646;
wire n_27647;
wire n_27648;
wire n_27649;
wire n_2765;
wire n_27650;
wire n_27651;
wire n_27652;
wire n_27653;
wire n_27654;
wire n_27655;
wire n_27656;
wire n_27657;
wire n_27658;
wire n_27659;
wire n_2766;
wire n_27660;
wire n_27661;
wire n_27662;
wire n_27663;
wire n_27664;
wire n_27665;
wire n_27666;
wire n_27667;
wire n_27668;
wire n_27669;
wire n_2767;
wire n_27670;
wire n_27671;
wire n_27672;
wire n_27673;
wire n_27674;
wire n_27675;
wire n_27676;
wire n_27677;
wire n_27678;
wire n_27679;
wire n_2768;
wire n_27680;
wire n_27681;
wire n_27682;
wire n_27684;
wire n_27685;
wire n_27686;
wire n_27687;
wire n_2769;
wire n_27690;
wire n_27691;
wire n_27692;
wire n_27693;
wire n_27694;
wire n_27695;
wire n_27696;
wire n_27698;
wire n_27699;
wire n_277;
wire n_2770;
wire n_27700;
wire n_27701;
wire n_27702;
wire n_27704;
wire n_27705;
wire n_27706;
wire n_27708;
wire n_27709;
wire n_2771;
wire n_27710;
wire n_27711;
wire n_27713;
wire n_27715;
wire n_27716;
wire n_27717;
wire n_27719;
wire n_2772;
wire n_27720;
wire n_27721;
wire n_27722;
wire n_27723;
wire n_27724;
wire n_27725;
wire n_27726;
wire n_27727;
wire n_27728;
wire n_27729;
wire n_2773;
wire n_27730;
wire n_27731;
wire n_27732;
wire n_27733;
wire n_27734;
wire n_27735;
wire n_27736;
wire n_27737;
wire n_27738;
wire n_27739;
wire n_2774;
wire n_27740;
wire n_27741;
wire n_27742;
wire n_27743;
wire n_27744;
wire n_27745;
wire n_27746;
wire n_27747;
wire n_27748;
wire n_27749;
wire n_2775;
wire n_27750;
wire n_27751;
wire n_27752;
wire n_27753;
wire n_27754;
wire n_27755;
wire n_27756;
wire n_27757;
wire n_27758;
wire n_27759;
wire n_2776;
wire n_27760;
wire n_27761;
wire n_27762;
wire n_27763;
wire n_27764;
wire n_27765;
wire n_27766;
wire n_27767;
wire n_27768;
wire n_27769;
wire n_2777;
wire n_27770;
wire n_27771;
wire n_27772;
wire n_27773;
wire n_27774;
wire n_27775;
wire n_27776;
wire n_27777;
wire n_27778;
wire n_27779;
wire n_2778;
wire n_27780;
wire n_27781;
wire n_27782;
wire n_27783;
wire n_27784;
wire n_27785;
wire n_27786;
wire n_27787;
wire n_27788;
wire n_27789;
wire n_2779;
wire n_27790;
wire n_27791;
wire n_27792;
wire n_27793;
wire n_27794;
wire n_27795;
wire n_27796;
wire n_27797;
wire n_27798;
wire n_27799;
wire n_278;
wire n_2780;
wire n_27800;
wire n_27801;
wire n_27802;
wire n_27803;
wire n_27804;
wire n_27805;
wire n_27806;
wire n_27807;
wire n_27808;
wire n_27809;
wire n_2781;
wire n_27810;
wire n_27811;
wire n_27812;
wire n_27813;
wire n_27814;
wire n_27815;
wire n_27816;
wire n_27817;
wire n_27818;
wire n_27819;
wire n_2782;
wire n_27820;
wire n_27821;
wire n_27822;
wire n_27823;
wire n_27824;
wire n_27825;
wire n_27826;
wire n_27827;
wire n_27828;
wire n_27829;
wire n_2783;
wire n_27830;
wire n_27831;
wire n_27832;
wire n_27833;
wire n_27834;
wire n_27835;
wire n_27836;
wire n_27837;
wire n_27838;
wire n_27839;
wire n_2784;
wire n_27840;
wire n_27841;
wire n_27842;
wire n_27843;
wire n_27844;
wire n_27845;
wire n_27846;
wire n_27847;
wire n_27848;
wire n_27849;
wire n_2785;
wire n_27850;
wire n_27851;
wire n_27852;
wire n_27853;
wire n_27854;
wire n_27855;
wire n_27856;
wire n_27857;
wire n_27858;
wire n_27859;
wire n_2786;
wire n_27860;
wire n_27861;
wire n_27862;
wire n_27863;
wire n_27864;
wire n_27865;
wire n_27866;
wire n_27867;
wire n_27868;
wire n_27869;
wire n_2787;
wire n_27870;
wire n_27871;
wire n_27872;
wire n_27873;
wire n_27874;
wire n_27875;
wire n_27876;
wire n_27877;
wire n_27878;
wire n_27879;
wire n_2788;
wire n_27880;
wire n_27881;
wire n_27882;
wire n_27883;
wire n_27884;
wire n_27885;
wire n_27886;
wire n_27887;
wire n_27888;
wire n_27889;
wire n_2789;
wire n_27890;
wire n_27891;
wire n_27892;
wire n_27893;
wire n_27894;
wire n_27895;
wire n_27897;
wire n_27898;
wire n_27899;
wire n_279;
wire n_2790;
wire n_27900;
wire n_27901;
wire n_27903;
wire n_27904;
wire n_27905;
wire n_27907;
wire n_27908;
wire n_27909;
wire n_2791;
wire n_27910;
wire n_27911;
wire n_27912;
wire n_27913;
wire n_27914;
wire n_27915;
wire n_27916;
wire n_27917;
wire n_27918;
wire n_27919;
wire n_2792;
wire n_27920;
wire n_27921;
wire n_27922;
wire n_27923;
wire n_27924;
wire n_27925;
wire n_27927;
wire n_27928;
wire n_2793;
wire n_27930;
wire n_27931;
wire n_27932;
wire n_27933;
wire n_27934;
wire n_27935;
wire n_27936;
wire n_27937;
wire n_27938;
wire n_27939;
wire n_2794;
wire n_27940;
wire n_27941;
wire n_27942;
wire n_27943;
wire n_27944;
wire n_27945;
wire n_27946;
wire n_27947;
wire n_27948;
wire n_27949;
wire n_2795;
wire n_27950;
wire n_27951;
wire n_27952;
wire n_27953;
wire n_27954;
wire n_27955;
wire n_27956;
wire n_27957;
wire n_27958;
wire n_27959;
wire n_2796;
wire n_27960;
wire n_27961;
wire n_27962;
wire n_27963;
wire n_27964;
wire n_27965;
wire n_27966;
wire n_27967;
wire n_27968;
wire n_27969;
wire n_2797;
wire n_27970;
wire n_27971;
wire n_27972;
wire n_27973;
wire n_27974;
wire n_27975;
wire n_27976;
wire n_27977;
wire n_27978;
wire n_27979;
wire n_2798;
wire n_27980;
wire n_27981;
wire n_27982;
wire n_27983;
wire n_27984;
wire n_27985;
wire n_27986;
wire n_27987;
wire n_27989;
wire n_2799;
wire n_27990;
wire n_27991;
wire n_27992;
wire n_27993;
wire n_27994;
wire n_27995;
wire n_27996;
wire n_27998;
wire n_27999;
wire n_28;
wire n_280;
wire n_2800;
wire n_28000;
wire n_28001;
wire n_28002;
wire n_28003;
wire n_28004;
wire n_28005;
wire n_28006;
wire n_28007;
wire n_28008;
wire n_28009;
wire n_2801;
wire n_28010;
wire n_28011;
wire n_28012;
wire n_28013;
wire n_28015;
wire n_28016;
wire n_28017;
wire n_28018;
wire n_28019;
wire n_2802;
wire n_28020;
wire n_28021;
wire n_28022;
wire n_28023;
wire n_28024;
wire n_28025;
wire n_28026;
wire n_28027;
wire n_28028;
wire n_28029;
wire n_2803;
wire n_28030;
wire n_28031;
wire n_28032;
wire n_28033;
wire n_28034;
wire n_28035;
wire n_28036;
wire n_28037;
wire n_28039;
wire n_2804;
wire n_28040;
wire n_28041;
wire n_28042;
wire n_28043;
wire n_28044;
wire n_28045;
wire n_28046;
wire n_28047;
wire n_28048;
wire n_28049;
wire n_2805;
wire n_28050;
wire n_28051;
wire n_28052;
wire n_28053;
wire n_28054;
wire n_28055;
wire n_28056;
wire n_28057;
wire n_28058;
wire n_28059;
wire n_2806;
wire n_28060;
wire n_28061;
wire n_28062;
wire n_28063;
wire n_28064;
wire n_28065;
wire n_28066;
wire n_28067;
wire n_28068;
wire n_28069;
wire n_2807;
wire n_28070;
wire n_28071;
wire n_28072;
wire n_28073;
wire n_28074;
wire n_28075;
wire n_28076;
wire n_28077;
wire n_28078;
wire n_28079;
wire n_2808;
wire n_28080;
wire n_28081;
wire n_28082;
wire n_28083;
wire n_28085;
wire n_28086;
wire n_28087;
wire n_28088;
wire n_28089;
wire n_2809;
wire n_28090;
wire n_28091;
wire n_28092;
wire n_28093;
wire n_28094;
wire n_28095;
wire n_28096;
wire n_28097;
wire n_28098;
wire n_28099;
wire n_281;
wire n_2810;
wire n_28100;
wire n_28101;
wire n_28102;
wire n_28103;
wire n_28104;
wire n_28105;
wire n_28107;
wire n_28108;
wire n_28109;
wire n_2811;
wire n_28110;
wire n_28111;
wire n_28112;
wire n_28113;
wire n_28114;
wire n_28115;
wire n_28116;
wire n_28117;
wire n_28118;
wire n_28119;
wire n_2812;
wire n_28120;
wire n_28121;
wire n_28122;
wire n_28123;
wire n_28124;
wire n_28125;
wire n_28126;
wire n_28127;
wire n_28128;
wire n_28129;
wire n_2813;
wire n_28130;
wire n_28131;
wire n_28132;
wire n_28133;
wire n_28134;
wire n_28135;
wire n_28136;
wire n_28137;
wire n_28138;
wire n_28139;
wire n_28140;
wire n_28141;
wire n_28142;
wire n_28144;
wire n_28145;
wire n_28146;
wire n_28147;
wire n_28148;
wire n_28149;
wire n_2815;
wire n_28150;
wire n_28151;
wire n_28152;
wire n_28153;
wire n_28154;
wire n_28155;
wire n_28156;
wire n_28157;
wire n_28158;
wire n_28159;
wire n_2816;
wire n_28160;
wire n_28161;
wire n_28162;
wire n_28163;
wire n_28164;
wire n_28165;
wire n_28166;
wire n_28167;
wire n_28168;
wire n_28169;
wire n_2817;
wire n_28170;
wire n_28171;
wire n_28172;
wire n_28173;
wire n_28174;
wire n_28175;
wire n_28176;
wire n_28177;
wire n_28178;
wire n_28179;
wire n_2818;
wire n_28180;
wire n_28181;
wire n_28182;
wire n_28183;
wire n_28184;
wire n_28185;
wire n_28186;
wire n_28187;
wire n_28188;
wire n_28189;
wire n_2819;
wire n_28190;
wire n_28191;
wire n_28192;
wire n_28193;
wire n_28194;
wire n_28195;
wire n_28196;
wire n_28197;
wire n_28198;
wire n_28199;
wire n_282;
wire n_2820;
wire n_28200;
wire n_28201;
wire n_28202;
wire n_28203;
wire n_28204;
wire n_28205;
wire n_28206;
wire n_28207;
wire n_28208;
wire n_28209;
wire n_2821;
wire n_28210;
wire n_28212;
wire n_28213;
wire n_28214;
wire n_28215;
wire n_28216;
wire n_28217;
wire n_28218;
wire n_28219;
wire n_2822;
wire n_28220;
wire n_28221;
wire n_28222;
wire n_28223;
wire n_28224;
wire n_28225;
wire n_28226;
wire n_28227;
wire n_28228;
wire n_28229;
wire n_2823;
wire n_28230;
wire n_28231;
wire n_28232;
wire n_28233;
wire n_28234;
wire n_28235;
wire n_28236;
wire n_28237;
wire n_28238;
wire n_28239;
wire n_2824;
wire n_28240;
wire n_28241;
wire n_28242;
wire n_28243;
wire n_28244;
wire n_28245;
wire n_28246;
wire n_28247;
wire n_28248;
wire n_28249;
wire n_2825;
wire n_28250;
wire n_28251;
wire n_28252;
wire n_28253;
wire n_28254;
wire n_28255;
wire n_28256;
wire n_28257;
wire n_28258;
wire n_2826;
wire n_28260;
wire n_28261;
wire n_28263;
wire n_28264;
wire n_28265;
wire n_28266;
wire n_28267;
wire n_28268;
wire n_28269;
wire n_2827;
wire n_28270;
wire n_28271;
wire n_28272;
wire n_28273;
wire n_28274;
wire n_28275;
wire n_28276;
wire n_28277;
wire n_28278;
wire n_28279;
wire n_2828;
wire n_28280;
wire n_28281;
wire n_28282;
wire n_28283;
wire n_28284;
wire n_28285;
wire n_28286;
wire n_28287;
wire n_28288;
wire n_28289;
wire n_2829;
wire n_28290;
wire n_28291;
wire n_28294;
wire n_28295;
wire n_28297;
wire n_28298;
wire n_28299;
wire n_283;
wire n_2830;
wire n_28301;
wire n_28302;
wire n_28303;
wire n_28304;
wire n_28306;
wire n_28308;
wire n_2831;
wire n_28310;
wire n_28312;
wire n_28314;
wire n_28315;
wire n_28316;
wire n_28317;
wire n_28318;
wire n_28319;
wire n_2832;
wire n_28320;
wire n_28321;
wire n_28322;
wire n_28323;
wire n_28324;
wire n_28325;
wire n_28326;
wire n_28327;
wire n_28328;
wire n_28329;
wire n_2833;
wire n_28330;
wire n_28331;
wire n_28332;
wire n_28333;
wire n_28334;
wire n_28335;
wire n_28336;
wire n_28337;
wire n_28338;
wire n_28339;
wire n_2834;
wire n_28340;
wire n_28341;
wire n_28342;
wire n_28343;
wire n_28344;
wire n_28345;
wire n_28346;
wire n_28347;
wire n_28348;
wire n_28349;
wire n_2835;
wire n_28350;
wire n_28351;
wire n_28352;
wire n_28353;
wire n_28354;
wire n_28355;
wire n_28356;
wire n_28357;
wire n_28359;
wire n_2836;
wire n_28360;
wire n_28361;
wire n_28362;
wire n_28363;
wire n_28365;
wire n_28366;
wire n_28367;
wire n_28368;
wire n_28369;
wire n_2837;
wire n_28370;
wire n_28371;
wire n_28372;
wire n_28373;
wire n_28374;
wire n_28375;
wire n_28376;
wire n_28377;
wire n_28378;
wire n_28379;
wire n_2838;
wire n_28380;
wire n_28381;
wire n_28382;
wire n_28383;
wire n_28384;
wire n_28385;
wire n_28386;
wire n_28387;
wire n_28388;
wire n_28389;
wire n_2839;
wire n_28390;
wire n_28391;
wire n_28392;
wire n_28393;
wire n_28394;
wire n_28396;
wire n_28397;
wire n_28398;
wire n_28399;
wire n_284;
wire n_2840;
wire n_28400;
wire n_28401;
wire n_28402;
wire n_28403;
wire n_28404;
wire n_28405;
wire n_28406;
wire n_28407;
wire n_28408;
wire n_28409;
wire n_2841;
wire n_28410;
wire n_28411;
wire n_28412;
wire n_28413;
wire n_28414;
wire n_28415;
wire n_28416;
wire n_28417;
wire n_28418;
wire n_28419;
wire n_2842;
wire n_28420;
wire n_28421;
wire n_28422;
wire n_28424;
wire n_28425;
wire n_28427;
wire n_28429;
wire n_2843;
wire n_28430;
wire n_28431;
wire n_28432;
wire n_28433;
wire n_28434;
wire n_28435;
wire n_28436;
wire n_28437;
wire n_28438;
wire n_28439;
wire n_2844;
wire n_28440;
wire n_28441;
wire n_28442;
wire n_28443;
wire n_28444;
wire n_28445;
wire n_28446;
wire n_28447;
wire n_28448;
wire n_28449;
wire n_2845;
wire n_28450;
wire n_28451;
wire n_28452;
wire n_28453;
wire n_28454;
wire n_28455;
wire n_28456;
wire n_28457;
wire n_28458;
wire n_28459;
wire n_2846;
wire n_28460;
wire n_28461;
wire n_28462;
wire n_28463;
wire n_28464;
wire n_28465;
wire n_28466;
wire n_28467;
wire n_28468;
wire n_28469;
wire n_2847;
wire n_28470;
wire n_28471;
wire n_28472;
wire n_28473;
wire n_28474;
wire n_28475;
wire n_28476;
wire n_28477;
wire n_28478;
wire n_2848;
wire n_28480;
wire n_28481;
wire n_28482;
wire n_28484;
wire n_28485;
wire n_28486;
wire n_28487;
wire n_28488;
wire n_28489;
wire n_2849;
wire n_28490;
wire n_28491;
wire n_28492;
wire n_28493;
wire n_28494;
wire n_28495;
wire n_28496;
wire n_28497;
wire n_28498;
wire n_28499;
wire n_285;
wire n_2850;
wire n_28500;
wire n_28501;
wire n_28502;
wire n_28503;
wire n_28504;
wire n_28505;
wire n_28506;
wire n_28507;
wire n_28508;
wire n_28509;
wire n_2851;
wire n_28510;
wire n_28511;
wire n_28513;
wire n_28515;
wire n_28516;
wire n_28517;
wire n_28518;
wire n_28519;
wire n_2852;
wire n_28520;
wire n_28521;
wire n_28522;
wire n_28523;
wire n_28524;
wire n_28525;
wire n_28527;
wire n_28528;
wire n_28529;
wire n_2853;
wire n_28530;
wire n_28531;
wire n_28532;
wire n_28533;
wire n_28534;
wire n_28535;
wire n_28536;
wire n_28537;
wire n_28538;
wire n_28539;
wire n_2854;
wire n_28540;
wire n_28541;
wire n_28542;
wire n_28543;
wire n_28544;
wire n_28545;
wire n_28546;
wire n_28547;
wire n_28548;
wire n_28549;
wire n_2855;
wire n_28550;
wire n_28551;
wire n_28552;
wire n_28553;
wire n_28554;
wire n_28555;
wire n_28556;
wire n_28557;
wire n_28558;
wire n_28559;
wire n_2856;
wire n_28560;
wire n_28561;
wire n_28562;
wire n_28563;
wire n_28564;
wire n_28565;
wire n_28566;
wire n_28567;
wire n_28568;
wire n_28569;
wire n_2857;
wire n_28570;
wire n_28571;
wire n_28572;
wire n_28573;
wire n_28574;
wire n_28575;
wire n_28576;
wire n_28577;
wire n_28578;
wire n_28579;
wire n_28580;
wire n_28581;
wire n_28582;
wire n_28583;
wire n_28584;
wire n_28585;
wire n_28586;
wire n_28587;
wire n_28588;
wire n_28589;
wire n_2859;
wire n_28590;
wire n_28591;
wire n_28592;
wire n_28593;
wire n_28594;
wire n_28595;
wire n_28597;
wire n_28598;
wire n_28599;
wire n_286;
wire n_2860;
wire n_28601;
wire n_28602;
wire n_28603;
wire n_28604;
wire n_28606;
wire n_28607;
wire n_28608;
wire n_28609;
wire n_2861;
wire n_28611;
wire n_28612;
wire n_28613;
wire n_28614;
wire n_28616;
wire n_28617;
wire n_28619;
wire n_2862;
wire n_28622;
wire n_28623;
wire n_28624;
wire n_28625;
wire n_28626;
wire n_28627;
wire n_28628;
wire n_28629;
wire n_2863;
wire n_28630;
wire n_28631;
wire n_28632;
wire n_28633;
wire n_28634;
wire n_28635;
wire n_28636;
wire n_28637;
wire n_28638;
wire n_28639;
wire n_2864;
wire n_28640;
wire n_28641;
wire n_28642;
wire n_28643;
wire n_28644;
wire n_28645;
wire n_28646;
wire n_28647;
wire n_28648;
wire n_28649;
wire n_2865;
wire n_28650;
wire n_28652;
wire n_28653;
wire n_28654;
wire n_28655;
wire n_28656;
wire n_28657;
wire n_28658;
wire n_28659;
wire n_2866;
wire n_28660;
wire n_28661;
wire n_28662;
wire n_28663;
wire n_28664;
wire n_28665;
wire n_28666;
wire n_28668;
wire n_28669;
wire n_2867;
wire n_28670;
wire n_28672;
wire n_28673;
wire n_28674;
wire n_28677;
wire n_28678;
wire n_28679;
wire n_2868;
wire n_28680;
wire n_28681;
wire n_28682;
wire n_28683;
wire n_28684;
wire n_28686;
wire n_28687;
wire n_28689;
wire n_2869;
wire n_28690;
wire n_28691;
wire n_28693;
wire n_28694;
wire n_28695;
wire n_28696;
wire n_28697;
wire n_28698;
wire n_28699;
wire n_287;
wire n_2870;
wire n_28700;
wire n_28701;
wire n_28702;
wire n_28703;
wire n_28704;
wire n_28705;
wire n_28706;
wire n_28707;
wire n_28708;
wire n_28709;
wire n_2871;
wire n_28710;
wire n_28712;
wire n_28713;
wire n_28714;
wire n_28715;
wire n_28716;
wire n_28717;
wire n_28718;
wire n_28719;
wire n_2872;
wire n_28720;
wire n_28721;
wire n_28722;
wire n_28723;
wire n_28724;
wire n_28725;
wire n_28726;
wire n_28727;
wire n_28728;
wire n_28729;
wire n_2873;
wire n_28730;
wire n_28731;
wire n_28732;
wire n_28733;
wire n_28734;
wire n_28735;
wire n_28736;
wire n_28737;
wire n_28738;
wire n_28739;
wire n_2874;
wire n_28740;
wire n_28741;
wire n_28742;
wire n_28743;
wire n_28744;
wire n_28745;
wire n_28746;
wire n_28747;
wire n_28748;
wire n_28749;
wire n_2875;
wire n_28750;
wire n_28751;
wire n_28752;
wire n_28753;
wire n_28754;
wire n_28755;
wire n_28756;
wire n_28757;
wire n_28758;
wire n_28759;
wire n_2876;
wire n_28760;
wire n_28761;
wire n_28762;
wire n_28763;
wire n_28764;
wire n_28765;
wire n_28766;
wire n_28767;
wire n_28769;
wire n_2877;
wire n_28770;
wire n_28771;
wire n_28772;
wire n_28773;
wire n_28774;
wire n_28775;
wire n_28776;
wire n_28777;
wire n_28778;
wire n_28779;
wire n_2878;
wire n_28780;
wire n_28781;
wire n_28782;
wire n_28783;
wire n_28784;
wire n_28785;
wire n_28786;
wire n_28787;
wire n_28788;
wire n_28789;
wire n_2879;
wire n_28790;
wire n_28791;
wire n_28792;
wire n_28793;
wire n_28794;
wire n_28795;
wire n_28796;
wire n_28797;
wire n_28798;
wire n_28799;
wire n_288;
wire n_2880;
wire n_28800;
wire n_28801;
wire n_28802;
wire n_28803;
wire n_28804;
wire n_28805;
wire n_28806;
wire n_28807;
wire n_28808;
wire n_28809;
wire n_2881;
wire n_28810;
wire n_28811;
wire n_28812;
wire n_28813;
wire n_28814;
wire n_28815;
wire n_28816;
wire n_28817;
wire n_28818;
wire n_28819;
wire n_2882;
wire n_28821;
wire n_28822;
wire n_28823;
wire n_28824;
wire n_28825;
wire n_28826;
wire n_28827;
wire n_28828;
wire n_28829;
wire n_2883;
wire n_28830;
wire n_28831;
wire n_28832;
wire n_28833;
wire n_28834;
wire n_28835;
wire n_28836;
wire n_28837;
wire n_28838;
wire n_28839;
wire n_2884;
wire n_28840;
wire n_28841;
wire n_28842;
wire n_28843;
wire n_28844;
wire n_28845;
wire n_28846;
wire n_28847;
wire n_28848;
wire n_28849;
wire n_2885;
wire n_28850;
wire n_28851;
wire n_28853;
wire n_28854;
wire n_28855;
wire n_28856;
wire n_28857;
wire n_28858;
wire n_28859;
wire n_2886;
wire n_28860;
wire n_28861;
wire n_28862;
wire n_28863;
wire n_28864;
wire n_28865;
wire n_28866;
wire n_28867;
wire n_28868;
wire n_2887;
wire n_28870;
wire n_28871;
wire n_28872;
wire n_28873;
wire n_28874;
wire n_28875;
wire n_28876;
wire n_28877;
wire n_28878;
wire n_28879;
wire n_2888;
wire n_28880;
wire n_28881;
wire n_28882;
wire n_28883;
wire n_28884;
wire n_28885;
wire n_28886;
wire n_28887;
wire n_28888;
wire n_28889;
wire n_2889;
wire n_28890;
wire n_28891;
wire n_28892;
wire n_28893;
wire n_28894;
wire n_28895;
wire n_28896;
wire n_28897;
wire n_28898;
wire n_28899;
wire n_289;
wire n_2890;
wire n_28900;
wire n_28901;
wire n_28902;
wire n_28903;
wire n_28904;
wire n_28905;
wire n_28906;
wire n_28907;
wire n_28908;
wire n_28909;
wire n_2891;
wire n_28910;
wire n_28911;
wire n_28912;
wire n_28913;
wire n_28914;
wire n_28915;
wire n_28917;
wire n_28919;
wire n_2892;
wire n_28920;
wire n_28921;
wire n_28923;
wire n_28925;
wire n_28926;
wire n_28927;
wire n_28928;
wire n_28929;
wire n_2893;
wire n_28931;
wire n_28932;
wire n_28933;
wire n_28934;
wire n_28935;
wire n_28936;
wire n_28937;
wire n_28938;
wire n_28939;
wire n_2894;
wire n_28940;
wire n_28941;
wire n_28942;
wire n_28943;
wire n_28944;
wire n_28945;
wire n_28948;
wire n_28949;
wire n_2895;
wire n_28950;
wire n_28951;
wire n_28952;
wire n_28953;
wire n_28954;
wire n_28955;
wire n_28956;
wire n_28957;
wire n_28958;
wire n_28959;
wire n_2896;
wire n_28960;
wire n_28961;
wire n_28962;
wire n_28963;
wire n_28964;
wire n_28965;
wire n_28966;
wire n_28967;
wire n_28968;
wire n_28969;
wire n_2897;
wire n_28970;
wire n_28971;
wire n_28972;
wire n_28973;
wire n_28974;
wire n_28975;
wire n_28976;
wire n_28977;
wire n_28978;
wire n_28979;
wire n_2898;
wire n_28980;
wire n_28981;
wire n_28982;
wire n_28983;
wire n_28984;
wire n_28985;
wire n_28986;
wire n_28987;
wire n_28988;
wire n_28989;
wire n_2899;
wire n_28990;
wire n_28991;
wire n_28992;
wire n_28993;
wire n_28994;
wire n_28995;
wire n_28996;
wire n_28997;
wire n_28998;
wire n_28999;
wire n_29;
wire n_290;
wire n_2900;
wire n_29000;
wire n_29001;
wire n_29002;
wire n_29003;
wire n_29004;
wire n_29005;
wire n_29006;
wire n_29007;
wire n_29008;
wire n_29009;
wire n_2901;
wire n_29010;
wire n_29011;
wire n_29012;
wire n_29013;
wire n_29014;
wire n_29015;
wire n_29016;
wire n_29017;
wire n_29018;
wire n_29019;
wire n_2902;
wire n_29020;
wire n_29021;
wire n_29023;
wire n_29024;
wire n_29026;
wire n_29027;
wire n_29029;
wire n_2903;
wire n_29030;
wire n_29031;
wire n_29033;
wire n_29034;
wire n_29035;
wire n_29036;
wire n_29037;
wire n_29038;
wire n_29039;
wire n_2904;
wire n_29040;
wire n_29042;
wire n_29043;
wire n_29045;
wire n_29046;
wire n_29047;
wire n_29049;
wire n_2905;
wire n_29050;
wire n_29051;
wire n_29052;
wire n_29053;
wire n_29054;
wire n_29055;
wire n_29056;
wire n_29057;
wire n_29058;
wire n_29059;
wire n_2906;
wire n_29060;
wire n_29061;
wire n_29062;
wire n_29063;
wire n_29064;
wire n_29065;
wire n_29066;
wire n_29067;
wire n_29068;
wire n_29069;
wire n_2907;
wire n_29070;
wire n_29071;
wire n_29072;
wire n_29073;
wire n_29074;
wire n_29075;
wire n_29076;
wire n_29077;
wire n_29078;
wire n_29079;
wire n_2908;
wire n_29080;
wire n_29081;
wire n_29082;
wire n_29083;
wire n_29084;
wire n_29085;
wire n_29086;
wire n_29087;
wire n_29088;
wire n_29089;
wire n_2909;
wire n_29090;
wire n_29091;
wire n_29092;
wire n_29093;
wire n_29094;
wire n_29095;
wire n_29096;
wire n_29097;
wire n_29098;
wire n_291;
wire n_2910;
wire n_29100;
wire n_29101;
wire n_29103;
wire n_29104;
wire n_29105;
wire n_29106;
wire n_29108;
wire n_29109;
wire n_2911;
wire n_29110;
wire n_29111;
wire n_29112;
wire n_29113;
wire n_29114;
wire n_29115;
wire n_29116;
wire n_29117;
wire n_29118;
wire n_29119;
wire n_2912;
wire n_29120;
wire n_29121;
wire n_29122;
wire n_29123;
wire n_29124;
wire n_29125;
wire n_29126;
wire n_29127;
wire n_29128;
wire n_29129;
wire n_2913;
wire n_29130;
wire n_29131;
wire n_29132;
wire n_29133;
wire n_29134;
wire n_29135;
wire n_29136;
wire n_29137;
wire n_29138;
wire n_29139;
wire n_2914;
wire n_29140;
wire n_29141;
wire n_29142;
wire n_29143;
wire n_29144;
wire n_29145;
wire n_29146;
wire n_29147;
wire n_29148;
wire n_29149;
wire n_2915;
wire n_29150;
wire n_29151;
wire n_29152;
wire n_29153;
wire n_29154;
wire n_29155;
wire n_29156;
wire n_29157;
wire n_29158;
wire n_29159;
wire n_2916;
wire n_29160;
wire n_29161;
wire n_29162;
wire n_29163;
wire n_29164;
wire n_29165;
wire n_29166;
wire n_29167;
wire n_29168;
wire n_29169;
wire n_2917;
wire n_29170;
wire n_29171;
wire n_29174;
wire n_29175;
wire n_29176;
wire n_29178;
wire n_29179;
wire n_2918;
wire n_29180;
wire n_29181;
wire n_29182;
wire n_29183;
wire n_29184;
wire n_29185;
wire n_29186;
wire n_29187;
wire n_29188;
wire n_29189;
wire n_2919;
wire n_29190;
wire n_29191;
wire n_29192;
wire n_29193;
wire n_29194;
wire n_29195;
wire n_29196;
wire n_29197;
wire n_29198;
wire n_29199;
wire n_292;
wire n_2920;
wire n_29200;
wire n_29201;
wire n_29202;
wire n_29203;
wire n_29204;
wire n_29205;
wire n_29206;
wire n_29207;
wire n_29208;
wire n_2921;
wire n_29210;
wire n_29211;
wire n_29212;
wire n_29213;
wire n_29214;
wire n_29215;
wire n_29216;
wire n_29217;
wire n_29218;
wire n_29219;
wire n_2922;
wire n_29220;
wire n_29221;
wire n_29222;
wire n_29223;
wire n_29224;
wire n_29225;
wire n_29226;
wire n_29227;
wire n_29228;
wire n_29229;
wire n_2923;
wire n_29230;
wire n_29231;
wire n_29232;
wire n_29233;
wire n_29234;
wire n_29235;
wire n_29236;
wire n_29237;
wire n_29238;
wire n_29239;
wire n_2924;
wire n_29240;
wire n_29241;
wire n_29242;
wire n_29243;
wire n_29244;
wire n_29245;
wire n_29246;
wire n_29247;
wire n_29248;
wire n_29249;
wire n_2925;
wire n_29250;
wire n_29251;
wire n_29252;
wire n_29253;
wire n_29254;
wire n_29256;
wire n_29257;
wire n_29258;
wire n_2926;
wire n_29260;
wire n_29261;
wire n_29263;
wire n_29264;
wire n_29265;
wire n_29266;
wire n_29268;
wire n_29269;
wire n_2927;
wire n_29270;
wire n_29271;
wire n_29272;
wire n_29273;
wire n_29274;
wire n_29275;
wire n_29276;
wire n_29277;
wire n_29278;
wire n_29279;
wire n_2928;
wire n_29280;
wire n_29281;
wire n_29282;
wire n_29283;
wire n_29284;
wire n_29285;
wire n_29286;
wire n_29287;
wire n_29288;
wire n_29289;
wire n_2929;
wire n_29290;
wire n_29291;
wire n_29292;
wire n_29293;
wire n_29294;
wire n_29295;
wire n_29296;
wire n_29297;
wire n_29298;
wire n_29299;
wire n_293;
wire n_2930;
wire n_29300;
wire n_29302;
wire n_29304;
wire n_29305;
wire n_29306;
wire n_29307;
wire n_29308;
wire n_29309;
wire n_2931;
wire n_29310;
wire n_29311;
wire n_29312;
wire n_29313;
wire n_29314;
wire n_29315;
wire n_29316;
wire n_29317;
wire n_29318;
wire n_29319;
wire n_2932;
wire n_29320;
wire n_29321;
wire n_29322;
wire n_29323;
wire n_29324;
wire n_29325;
wire n_29326;
wire n_29327;
wire n_29328;
wire n_29329;
wire n_2933;
wire n_29330;
wire n_29331;
wire n_29332;
wire n_29333;
wire n_29334;
wire n_29335;
wire n_29336;
wire n_29337;
wire n_29338;
wire n_2934;
wire n_29340;
wire n_29341;
wire n_29342;
wire n_29343;
wire n_29344;
wire n_29346;
wire n_29347;
wire n_29349;
wire n_2935;
wire n_29350;
wire n_29351;
wire n_29353;
wire n_29354;
wire n_29355;
wire n_29356;
wire n_29357;
wire n_29358;
wire n_29359;
wire n_2936;
wire n_29360;
wire n_29361;
wire n_29362;
wire n_29363;
wire n_29364;
wire n_29365;
wire n_29366;
wire n_29367;
wire n_29368;
wire n_29369;
wire n_2937;
wire n_29370;
wire n_29371;
wire n_29372;
wire n_29373;
wire n_29374;
wire n_29375;
wire n_29376;
wire n_29377;
wire n_29378;
wire n_29379;
wire n_2938;
wire n_29380;
wire n_29381;
wire n_29382;
wire n_29383;
wire n_29384;
wire n_29385;
wire n_29386;
wire n_29387;
wire n_29388;
wire n_29389;
wire n_2939;
wire n_29390;
wire n_29391;
wire n_29392;
wire n_29393;
wire n_29394;
wire n_29396;
wire n_29398;
wire n_29399;
wire n_294;
wire n_2940;
wire n_29400;
wire n_29401;
wire n_29403;
wire n_29404;
wire n_29406;
wire n_29408;
wire n_29409;
wire n_2941;
wire n_29410;
wire n_29411;
wire n_29412;
wire n_29413;
wire n_29415;
wire n_29416;
wire n_29417;
wire n_29418;
wire n_29419;
wire n_2942;
wire n_29420;
wire n_29421;
wire n_29422;
wire n_29423;
wire n_29424;
wire n_29425;
wire n_29426;
wire n_29427;
wire n_29428;
wire n_29429;
wire n_2943;
wire n_29430;
wire n_29431;
wire n_29432;
wire n_29433;
wire n_29434;
wire n_29435;
wire n_29437;
wire n_29438;
wire n_29439;
wire n_2944;
wire n_29440;
wire n_29441;
wire n_29442;
wire n_29443;
wire n_29444;
wire n_29446;
wire n_29447;
wire n_29448;
wire n_29449;
wire n_2945;
wire n_29450;
wire n_29451;
wire n_29452;
wire n_29454;
wire n_29455;
wire n_29456;
wire n_29457;
wire n_29458;
wire n_29459;
wire n_2946;
wire n_29460;
wire n_29462;
wire n_29463;
wire n_29464;
wire n_29465;
wire n_29466;
wire n_29467;
wire n_29468;
wire n_29469;
wire n_2947;
wire n_29470;
wire n_29471;
wire n_29472;
wire n_29473;
wire n_29474;
wire n_29475;
wire n_29476;
wire n_29477;
wire n_29478;
wire n_29479;
wire n_2948;
wire n_29480;
wire n_29481;
wire n_29482;
wire n_29483;
wire n_29484;
wire n_29485;
wire n_29486;
wire n_29487;
wire n_29488;
wire n_29489;
wire n_2949;
wire n_29490;
wire n_29491;
wire n_29492;
wire n_29493;
wire n_29494;
wire n_29495;
wire n_29496;
wire n_29497;
wire n_29498;
wire n_295;
wire n_2950;
wire n_29500;
wire n_29501;
wire n_29502;
wire n_29503;
wire n_29504;
wire n_29505;
wire n_29506;
wire n_29507;
wire n_29508;
wire n_29509;
wire n_2951;
wire n_29510;
wire n_29511;
wire n_29512;
wire n_29513;
wire n_29514;
wire n_29515;
wire n_29516;
wire n_29517;
wire n_29518;
wire n_29519;
wire n_2952;
wire n_29520;
wire n_29521;
wire n_29522;
wire n_29524;
wire n_29525;
wire n_29526;
wire n_29528;
wire n_2953;
wire n_29530;
wire n_29532;
wire n_29533;
wire n_29534;
wire n_29535;
wire n_29536;
wire n_29537;
wire n_29538;
wire n_29539;
wire n_2954;
wire n_29540;
wire n_29541;
wire n_29542;
wire n_29543;
wire n_29544;
wire n_29545;
wire n_29546;
wire n_29547;
wire n_29548;
wire n_29549;
wire n_2955;
wire n_29550;
wire n_29551;
wire n_29552;
wire n_29553;
wire n_29556;
wire n_29557;
wire n_29559;
wire n_2956;
wire n_29561;
wire n_29562;
wire n_29563;
wire n_29564;
wire n_29566;
wire n_29567;
wire n_29569;
wire n_2957;
wire n_29570;
wire n_29572;
wire n_29573;
wire n_29574;
wire n_29575;
wire n_29576;
wire n_29577;
wire n_29578;
wire n_29579;
wire n_2958;
wire n_29580;
wire n_29581;
wire n_29583;
wire n_29584;
wire n_29585;
wire n_29587;
wire n_29588;
wire n_29589;
wire n_2959;
wire n_29592;
wire n_29593;
wire n_29594;
wire n_29596;
wire n_29598;
wire n_296;
wire n_2960;
wire n_29600;
wire n_29601;
wire n_29602;
wire n_29603;
wire n_29604;
wire n_29605;
wire n_29606;
wire n_29607;
wire n_29608;
wire n_29609;
wire n_2961;
wire n_29611;
wire n_29612;
wire n_29613;
wire n_29614;
wire n_29616;
wire n_29617;
wire n_29618;
wire n_29619;
wire n_2962;
wire n_29620;
wire n_29622;
wire n_29623;
wire n_29624;
wire n_29625;
wire n_29626;
wire n_29627;
wire n_29629;
wire n_2963;
wire n_29630;
wire n_29631;
wire n_29632;
wire n_29633;
wire n_29634;
wire n_29635;
wire n_29636;
wire n_29638;
wire n_29639;
wire n_2964;
wire n_29640;
wire n_29641;
wire n_29642;
wire n_29643;
wire n_29644;
wire n_29646;
wire n_29647;
wire n_29649;
wire n_2965;
wire n_29650;
wire n_29651;
wire n_29652;
wire n_29653;
wire n_29654;
wire n_29656;
wire n_29657;
wire n_29658;
wire n_29659;
wire n_2966;
wire n_29660;
wire n_29662;
wire n_29664;
wire n_29665;
wire n_29667;
wire n_29668;
wire n_29669;
wire n_29670;
wire n_29672;
wire n_29673;
wire n_29674;
wire n_29675;
wire n_29676;
wire n_29677;
wire n_29678;
wire n_2968;
wire n_29680;
wire n_29681;
wire n_29682;
wire n_29683;
wire n_29684;
wire n_29685;
wire n_29686;
wire n_29687;
wire n_29688;
wire n_29689;
wire n_2969;
wire n_29691;
wire n_29692;
wire n_29693;
wire n_29694;
wire n_29695;
wire n_29696;
wire n_29698;
wire n_29699;
wire n_297;
wire n_2970;
wire n_29700;
wire n_29701;
wire n_29702;
wire n_29703;
wire n_29705;
wire n_29706;
wire n_29707;
wire n_29708;
wire n_29709;
wire n_2971;
wire n_29710;
wire n_2972;
wire n_2973;
wire n_2974;
wire n_2975;
wire n_2976;
wire n_2977;
wire n_2978;
wire n_2979;
wire n_298;
wire n_2980;
wire n_2981;
wire n_2982;
wire n_2983;
wire n_2984;
wire n_2985;
wire n_2986;
wire n_2987;
wire n_2988;
wire n_2989;
wire n_299;
wire n_2990;
wire n_2991;
wire n_2992;
wire n_2993;
wire n_2994;
wire n_2995;
wire n_2996;
wire n_2997;
wire n_2998;
wire n_2999;
wire n_3;
wire n_30;
wire n_300;
wire n_3000;
wire n_3001;
wire n_3002;
wire n_3003;
wire n_3004;
wire n_3005;
wire n_3006;
wire n_3007;
wire n_3008;
wire n_3009;
wire n_301;
wire n_3010;
wire n_3011;
wire n_3012;
wire n_3013;
wire n_3014;
wire n_3015;
wire n_3016;
wire n_3017;
wire n_3018;
wire n_3019;
wire n_302;
wire n_3020;
wire n_3021;
wire n_3022;
wire n_3023;
wire n_3024;
wire n_3025;
wire n_3026;
wire n_3027;
wire n_3028;
wire n_3029;
wire n_303;
wire n_3030;
wire n_3031;
wire n_3032;
wire n_3033;
wire n_3034;
wire n_3035;
wire n_3036;
wire n_3037;
wire n_3038;
wire n_3039;
wire n_304;
wire n_3040;
wire n_3041;
wire n_3042;
wire n_3043;
wire n_3044;
wire n_3045;
wire n_3046;
wire n_3047;
wire n_3048;
wire n_3049;
wire n_305;
wire n_3050;
wire n_3051;
wire n_3052;
wire n_3053;
wire n_3054;
wire n_3055;
wire n_3056;
wire n_3057;
wire n_3058;
wire n_3059;
wire n_306;
wire n_3060;
wire n_3061;
wire n_3062;
wire n_3063;
wire n_3064;
wire n_3065;
wire n_3066;
wire n_3067;
wire n_3068;
wire n_307;
wire n_3070;
wire n_3071;
wire n_3072;
wire n_3073;
wire n_3074;
wire n_3075;
wire n_3076;
wire n_3077;
wire n_3078;
wire n_3079;
wire n_308;
wire n_3080;
wire n_3081;
wire n_3082;
wire n_3083;
wire n_3084;
wire n_3085;
wire n_3086;
wire n_3087;
wire n_3088;
wire n_3089;
wire n_309;
wire n_3090;
wire n_3091;
wire n_3092;
wire n_3093;
wire n_3094;
wire n_3095;
wire n_3096;
wire n_3097;
wire n_3098;
wire n_3099;
wire n_31;
wire n_310;
wire n_3100;
wire n_3101;
wire n_3102;
wire n_3103;
wire n_3104;
wire n_3105;
wire n_3106;
wire n_3107;
wire n_3108;
wire n_3109;
wire n_311;
wire n_3110;
wire n_3111;
wire n_3112;
wire n_3113;
wire n_3114;
wire n_3115;
wire n_3116;
wire n_3117;
wire n_3118;
wire n_3119;
wire n_312;
wire n_3120;
wire n_3121;
wire n_3122;
wire n_3123;
wire n_3124;
wire n_3125;
wire n_3126;
wire n_3127;
wire n_3128;
wire n_3129;
wire n_313;
wire n_3130;
wire n_3131;
wire n_3132;
wire n_3133;
wire n_3134;
wire n_3135;
wire n_3136;
wire n_3137;
wire n_3138;
wire n_3139;
wire n_314;
wire n_3140;
wire n_3141;
wire n_3142;
wire n_3143;
wire n_3144;
wire n_3145;
wire n_3146;
wire n_3147;
wire n_3148;
wire n_3149;
wire n_315;
wire n_3150;
wire n_3151;
wire n_3152;
wire n_3153;
wire n_3154;
wire n_3155;
wire n_3156;
wire n_3157;
wire n_3158;
wire n_3159;
wire n_316;
wire n_3160;
wire n_3161;
wire n_3162;
wire n_3163;
wire n_3164;
wire n_3165;
wire n_3166;
wire n_3167;
wire n_3168;
wire n_3169;
wire n_317;
wire n_3170;
wire n_3171;
wire n_3172;
wire n_3173;
wire n_3174;
wire n_3175;
wire n_3176;
wire n_3177;
wire n_3178;
wire n_3179;
wire n_318;
wire n_3180;
wire n_3181;
wire n_3182;
wire n_3183;
wire n_3184;
wire n_3185;
wire n_3186;
wire n_3187;
wire n_3188;
wire n_3189;
wire n_319;
wire n_3190;
wire n_3191;
wire n_3192;
wire n_3193;
wire n_3194;
wire n_3195;
wire n_3196;
wire n_3197;
wire n_3198;
wire n_3199;
wire n_32;
wire n_320;
wire n_3200;
wire n_3201;
wire n_3202;
wire n_3203;
wire n_3204;
wire n_3205;
wire n_3206;
wire n_3207;
wire n_3208;
wire n_3209;
wire n_321;
wire n_3210;
wire n_3211;
wire n_3212;
wire n_3213;
wire n_3214;
wire n_3215;
wire n_3216;
wire n_3217;
wire n_3218;
wire n_3219;
wire n_322;
wire n_3220;
wire n_3221;
wire n_3222;
wire n_3223;
wire n_3224;
wire n_3225;
wire n_3226;
wire n_3227;
wire n_3228;
wire n_3229;
wire n_323;
wire n_3230;
wire n_3231;
wire n_3232;
wire n_3233;
wire n_3234;
wire n_3235;
wire n_3236;
wire n_3237;
wire n_3238;
wire n_3239;
wire n_324;
wire n_3240;
wire n_3241;
wire n_3242;
wire n_3243;
wire n_3244;
wire n_3245;
wire n_3246;
wire n_3247;
wire n_3248;
wire n_3249;
wire n_325;
wire n_3250;
wire n_3251;
wire n_3252;
wire n_3253;
wire n_3254;
wire n_3255;
wire n_3256;
wire n_3257;
wire n_3258;
wire n_3259;
wire n_326;
wire n_3260;
wire n_3261;
wire n_3262;
wire n_3263;
wire n_3264;
wire n_3266;
wire n_3267;
wire n_3268;
wire n_3269;
wire n_327;
wire n_3270;
wire n_3271;
wire n_3272;
wire n_32729;
wire n_3273;
wire n_32730;
wire n_32731;
wire n_32732;
wire n_32733;
wire n_32734;
wire n_32735;
wire n_32736;
wire n_32737;
wire n_32738;
wire n_32739;
wire n_3274;
wire n_32740;
wire n_32741;
wire n_32742;
wire n_32743;
wire n_32744;
wire n_3275;
wire n_3276;
wire n_3277;
wire n_3278;
wire n_3279;
wire n_328;
wire n_3280;
wire n_3281;
wire n_3282;
wire n_3283;
wire n_3284;
wire n_3285;
wire n_3286;
wire n_3287;
wire n_3288;
wire n_3289;
wire n_329;
wire n_3290;
wire n_3291;
wire n_3292;
wire n_3293;
wire n_3294;
wire n_3295;
wire n_3296;
wire n_3297;
wire n_3298;
wire n_3299;
wire n_33;
wire n_330;
wire n_3300;
wire n_3301;
wire n_3302;
wire n_3303;
wire n_3304;
wire n_3305;
wire n_3306;
wire n_3307;
wire n_3308;
wire n_3309;
wire n_331;
wire n_3310;
wire n_3311;
wire n_3312;
wire n_3313;
wire n_3314;
wire n_3315;
wire n_3316;
wire n_3317;
wire n_3318;
wire n_3319;
wire n_332;
wire n_3320;
wire n_3321;
wire n_3322;
wire n_3323;
wire n_3324;
wire n_3325;
wire n_3326;
wire n_3327;
wire n_3328;
wire n_3329;
wire n_333;
wire n_3330;
wire n_3331;
wire n_3332;
wire n_3333;
wire n_3334;
wire n_3335;
wire n_3336;
wire n_3337;
wire n_3338;
wire n_3339;
wire n_334;
wire n_3340;
wire n_3341;
wire n_3342;
wire n_3343;
wire n_3344;
wire n_3345;
wire n_3346;
wire n_3347;
wire n_3348;
wire n_3349;
wire n_335;
wire n_3350;
wire n_3351;
wire n_3352;
wire n_3353;
wire n_3354;
wire n_3355;
wire n_3356;
wire n_3357;
wire n_3358;
wire n_3359;
wire n_336;
wire n_3360;
wire n_3361;
wire n_3362;
wire n_3363;
wire n_3364;
wire n_3365;
wire n_3366;
wire n_3367;
wire n_3368;
wire n_3369;
wire n_337;
wire n_3370;
wire n_3371;
wire n_3372;
wire n_3373;
wire n_3374;
wire n_3375;
wire n_3376;
wire n_3377;
wire n_3378;
wire n_3379;
wire n_338;
wire n_3380;
wire n_3381;
wire n_3382;
wire n_3383;
wire n_3384;
wire n_3385;
wire n_3386;
wire n_3387;
wire n_3388;
wire n_3389;
wire n_339;
wire n_3390;
wire n_3391;
wire n_3392;
wire n_3393;
wire n_3394;
wire n_3395;
wire n_3396;
wire n_3397;
wire n_3398;
wire n_3399;
wire n_34;
wire n_340;
wire n_3400;
wire n_3401;
wire n_3403;
wire n_3404;
wire n_3406;
wire n_3407;
wire n_3409;
wire n_341;
wire n_3410;
wire n_3414;
wire n_3415;
wire n_3416;
wire n_3417;
wire n_3418;
wire n_3419;
wire n_342;
wire n_3420;
wire n_3421;
wire n_3422;
wire n_3423;
wire n_3424;
wire n_3425;
wire n_3426;
wire n_3427;
wire n_343;
wire n_3430;
wire n_3431;
wire n_3432;
wire n_3433;
wire n_3434;
wire n_3435;
wire n_3436;
wire n_3437;
wire n_3438;
wire n_3439;
wire n_344;
wire n_3440;
wire n_3441;
wire n_3445;
wire n_3446;
wire n_3447;
wire n_3448;
wire n_3449;
wire n_345;
wire n_3450;
wire n_3451;
wire n_3452;
wire n_3453;
wire n_3455;
wire n_3456;
wire n_3457;
wire n_3458;
wire n_3459;
wire n_346;
wire n_3460;
wire n_3461;
wire n_3462;
wire n_3464;
wire n_3465;
wire n_3466;
wire n_3467;
wire n_3468;
wire n_3469;
wire n_347;
wire n_3470;
wire n_3471;
wire n_3472;
wire n_3473;
wire n_3474;
wire n_3475;
wire n_3476;
wire n_3477;
wire n_3478;
wire n_348;
wire n_3481;
wire n_3482;
wire n_3483;
wire n_3484;
wire n_3485;
wire n_3486;
wire n_3487;
wire n_3488;
wire n_3489;
wire n_349;
wire n_3490;
wire n_3491;
wire n_3492;
wire n_3493;
wire n_3494;
wire n_3495;
wire n_3496;
wire n_3498;
wire n_3499;
wire n_35;
wire n_350;
wire n_3500;
wire n_3501;
wire n_3502;
wire n_3503;
wire n_3504;
wire n_3505;
wire n_3506;
wire n_3507;
wire n_3508;
wire n_3509;
wire n_351;
wire n_3510;
wire n_3511;
wire n_3512;
wire n_3513;
wire n_3514;
wire n_3515;
wire n_3516;
wire n_3517;
wire n_3518;
wire n_3519;
wire n_352;
wire n_3520;
wire n_3521;
wire n_3522;
wire n_3523;
wire n_3524;
wire n_3525;
wire n_3526;
wire n_3527;
wire n_3528;
wire n_3529;
wire n_353;
wire n_3530;
wire n_3531;
wire n_3532;
wire n_3533;
wire n_3534;
wire n_3535;
wire n_3536;
wire n_3537;
wire n_3538;
wire n_3539;
wire n_354;
wire n_3540;
wire n_3541;
wire n_3542;
wire n_3543;
wire n_3544;
wire n_3545;
wire n_3546;
wire n_3547;
wire n_3548;
wire n_3549;
wire n_355;
wire n_3550;
wire n_3551;
wire n_3552;
wire n_3553;
wire n_3554;
wire n_3555;
wire n_3557;
wire n_3558;
wire n_3559;
wire n_356;
wire n_3560;
wire n_3561;
wire n_3562;
wire n_3563;
wire n_3564;
wire n_3565;
wire n_3566;
wire n_3568;
wire n_3569;
wire n_357;
wire n_3570;
wire n_3571;
wire n_3572;
wire n_3573;
wire n_3574;
wire n_3575;
wire n_3576;
wire n_3577;
wire n_3578;
wire n_3579;
wire n_358;
wire n_3580;
wire n_3581;
wire n_3582;
wire n_3583;
wire n_3584;
wire n_3585;
wire n_3586;
wire n_3587;
wire n_3588;
wire n_3589;
wire n_359;
wire n_3590;
wire n_3591;
wire n_3592;
wire n_3593;
wire n_3594;
wire n_3595;
wire n_3596;
wire n_3597;
wire n_3598;
wire n_3599;
wire n_36;
wire n_360;
wire n_3600;
wire n_3601;
wire n_3602;
wire n_3603;
wire n_3604;
wire n_3605;
wire n_3606;
wire n_3607;
wire n_3608;
wire n_3609;
wire n_361;
wire n_3611;
wire n_3612;
wire n_3613;
wire n_3614;
wire n_3615;
wire n_3616;
wire n_3617;
wire n_3618;
wire n_3619;
wire n_362;
wire n_3620;
wire n_3621;
wire n_3622;
wire n_3623;
wire n_3624;
wire n_3625;
wire n_3626;
wire n_3627;
wire n_3628;
wire n_3629;
wire n_363;
wire n_3630;
wire n_3631;
wire n_3632;
wire n_3633;
wire n_3634;
wire n_3635;
wire n_3636;
wire n_3637;
wire n_3638;
wire n_3639;
wire n_364;
wire n_3640;
wire n_3641;
wire n_3642;
wire n_3643;
wire n_3644;
wire n_3645;
wire n_3646;
wire n_3647;
wire n_3648;
wire n_3649;
wire n_365;
wire n_3650;
wire n_3651;
wire n_3652;
wire n_3653;
wire n_3654;
wire n_3655;
wire n_3656;
wire n_3657;
wire n_3658;
wire n_3659;
wire n_366;
wire n_3660;
wire n_3661;
wire n_3662;
wire n_3663;
wire n_3664;
wire n_3665;
wire n_3666;
wire n_3667;
wire n_3668;
wire n_3669;
wire n_367;
wire n_3670;
wire n_3671;
wire n_3672;
wire n_3673;
wire n_3674;
wire n_3675;
wire n_3676;
wire n_3677;
wire n_3678;
wire n_3679;
wire n_368;
wire n_3680;
wire n_3681;
wire n_3682;
wire n_3683;
wire n_3684;
wire n_3685;
wire n_3686;
wire n_3687;
wire n_3688;
wire n_3689;
wire n_369;
wire n_3690;
wire n_3691;
wire n_3692;
wire n_3693;
wire n_3694;
wire n_3695;
wire n_3696;
wire n_3697;
wire n_3698;
wire n_3699;
wire n_37;
wire n_370;
wire n_3700;
wire n_3701;
wire n_3702;
wire n_3703;
wire n_3704;
wire n_3705;
wire n_3706;
wire n_3707;
wire n_3708;
wire n_3709;
wire n_371;
wire n_3710;
wire n_3711;
wire n_3712;
wire n_3713;
wire n_3714;
wire n_3715;
wire n_3716;
wire n_3717;
wire n_3718;
wire n_3719;
wire n_372;
wire n_3720;
wire n_3721;
wire n_3722;
wire n_3723;
wire n_3724;
wire n_3725;
wire n_3726;
wire n_3727;
wire n_3728;
wire n_3729;
wire n_373;
wire n_3730;
wire n_3731;
wire n_3732;
wire n_3733;
wire n_3734;
wire n_3735;
wire n_3736;
wire n_3737;
wire n_3738;
wire n_3739;
wire n_374;
wire n_3740;
wire n_3741;
wire n_3742;
wire n_3743;
wire n_3744;
wire n_3745;
wire n_3746;
wire n_3747;
wire n_3748;
wire n_3749;
wire n_375;
wire n_3750;
wire n_3751;
wire n_3752;
wire n_3753;
wire n_3754;
wire n_3755;
wire n_3756;
wire n_3757;
wire n_3758;
wire n_3759;
wire n_376;
wire n_3760;
wire n_3761;
wire n_3762;
wire n_3763;
wire n_3764;
wire n_3765;
wire n_3766;
wire n_3767;
wire n_3768;
wire n_3769;
wire n_377;
wire n_3770;
wire n_3771;
wire n_3772;
wire n_3773;
wire n_3774;
wire n_3775;
wire n_3776;
wire n_3777;
wire n_3778;
wire n_3779;
wire n_378;
wire n_3780;
wire n_3781;
wire n_3782;
wire n_3783;
wire n_3784;
wire n_3785;
wire n_3786;
wire n_3787;
wire n_3788;
wire n_3789;
wire n_379;
wire n_3790;
wire n_3791;
wire n_3792;
wire n_3793;
wire n_3795;
wire n_3796;
wire n_3797;
wire n_3798;
wire n_3799;
wire n_38;
wire n_380;
wire n_3800;
wire n_3801;
wire n_3802;
wire n_3803;
wire n_3804;
wire n_3805;
wire n_3806;
wire n_3807;
wire n_3808;
wire n_3809;
wire n_381;
wire n_3811;
wire n_3812;
wire n_3813;
wire n_3814;
wire n_3815;
wire n_3816;
wire n_3817;
wire n_3818;
wire n_3819;
wire n_382;
wire n_3820;
wire n_3821;
wire n_3822;
wire n_3823;
wire n_3824;
wire n_3825;
wire n_3826;
wire n_3827;
wire n_3828;
wire n_3829;
wire n_383;
wire n_3830;
wire n_3831;
wire n_3832;
wire n_3833;
wire n_3834;
wire n_3835;
wire n_3836;
wire n_3837;
wire n_3838;
wire n_3839;
wire n_384;
wire n_3840;
wire n_3841;
wire n_3842;
wire n_3843;
wire n_3844;
wire n_3845;
wire n_3846;
wire n_3847;
wire n_3848;
wire n_3849;
wire n_385;
wire n_3850;
wire n_3851;
wire n_3852;
wire n_3853;
wire n_3854;
wire n_3855;
wire n_3856;
wire n_3857;
wire n_3858;
wire n_3859;
wire n_386;
wire n_3860;
wire n_3861;
wire n_3862;
wire n_3863;
wire n_3864;
wire n_3865;
wire n_3866;
wire n_3867;
wire n_3868;
wire n_3869;
wire n_387;
wire n_3870;
wire n_3871;
wire n_3872;
wire n_3873;
wire n_3874;
wire n_3875;
wire n_3876;
wire n_3877;
wire n_3878;
wire n_3879;
wire n_388;
wire n_3880;
wire n_3881;
wire n_3882;
wire n_3883;
wire n_3884;
wire n_3885;
wire n_3886;
wire n_3887;
wire n_3888;
wire n_3889;
wire n_389;
wire n_3890;
wire n_3891;
wire n_3892;
wire n_3893;
wire n_3894;
wire n_3895;
wire n_3896;
wire n_3897;
wire n_3898;
wire n_3899;
wire n_39;
wire n_390;
wire n_3900;
wire n_3901;
wire n_3902;
wire n_3903;
wire n_3904;
wire n_3905;
wire n_3906;
wire n_3907;
wire n_3908;
wire n_3909;
wire n_391;
wire n_3910;
wire n_3911;
wire n_3912;
wire n_3913;
wire n_3914;
wire n_3915;
wire n_3916;
wire n_3917;
wire n_3918;
wire n_392;
wire n_3920;
wire n_3921;
wire n_3922;
wire n_3923;
wire n_3924;
wire n_3925;
wire n_3926;
wire n_3927;
wire n_3928;
wire n_3929;
wire n_393;
wire n_3930;
wire n_3931;
wire n_3932;
wire n_3933;
wire n_3934;
wire n_3935;
wire n_3936;
wire n_3937;
wire n_3938;
wire n_3939;
wire n_394;
wire n_3940;
wire n_3941;
wire n_3942;
wire n_3943;
wire n_3944;
wire n_3945;
wire n_3946;
wire n_3947;
wire n_3948;
wire n_3949;
wire n_395;
wire n_3950;
wire n_3951;
wire n_3952;
wire n_3953;
wire n_3954;
wire n_3955;
wire n_3956;
wire n_3957;
wire n_3958;
wire n_3959;
wire n_396;
wire n_3960;
wire n_3961;
wire n_3962;
wire n_3963;
wire n_3964;
wire n_3965;
wire n_3966;
wire n_3967;
wire n_3968;
wire n_3969;
wire n_397;
wire n_3970;
wire n_3971;
wire n_3972;
wire n_3973;
wire n_3974;
wire n_3975;
wire n_3976;
wire n_3977;
wire n_3978;
wire n_3979;
wire n_398;
wire n_3980;
wire n_3981;
wire n_3982;
wire n_3983;
wire n_3984;
wire n_3985;
wire n_3986;
wire n_3987;
wire n_3988;
wire n_3989;
wire n_399;
wire n_3990;
wire n_3991;
wire n_3992;
wire n_3993;
wire n_3994;
wire n_3995;
wire n_3996;
wire n_3997;
wire n_3998;
wire n_3999;
wire n_4;
wire n_40;
wire n_400;
wire n_4000;
wire n_4001;
wire n_4002;
wire n_4003;
wire n_4004;
wire n_4005;
wire n_4006;
wire n_4007;
wire n_4008;
wire n_4009;
wire n_401;
wire n_4010;
wire n_4011;
wire n_4012;
wire n_4013;
wire n_4014;
wire n_4015;
wire n_4016;
wire n_4017;
wire n_4018;
wire n_4019;
wire n_402;
wire n_4020;
wire n_4021;
wire n_4022;
wire n_4023;
wire n_4024;
wire n_4025;
wire n_4026;
wire n_4027;
wire n_4028;
wire n_4029;
wire n_403;
wire n_4030;
wire n_4031;
wire n_4032;
wire n_4033;
wire n_4034;
wire n_4035;
wire n_4036;
wire n_4037;
wire n_4039;
wire n_404;
wire n_4040;
wire n_4041;
wire n_4042;
wire n_4043;
wire n_4044;
wire n_4045;
wire n_4046;
wire n_4047;
wire n_4048;
wire n_4049;
wire n_405;
wire n_4050;
wire n_4051;
wire n_4052;
wire n_4053;
wire n_4054;
wire n_4055;
wire n_4056;
wire n_4057;
wire n_4058;
wire n_4059;
wire n_406;
wire n_4060;
wire n_4061;
wire n_4062;
wire n_4063;
wire n_4064;
wire n_4065;
wire n_4066;
wire n_4067;
wire n_4068;
wire n_4069;
wire n_407;
wire n_4070;
wire n_4071;
wire n_4072;
wire n_4074;
wire n_4075;
wire n_4076;
wire n_4077;
wire n_4078;
wire n_408;
wire n_4080;
wire n_4081;
wire n_4082;
wire n_4083;
wire n_4084;
wire n_4085;
wire n_4086;
wire n_4087;
wire n_4088;
wire n_4089;
wire n_409;
wire n_4090;
wire n_4091;
wire n_4092;
wire n_4093;
wire n_4094;
wire n_4095;
wire n_4097;
wire n_4098;
wire n_4099;
wire n_41;
wire n_410;
wire n_4100;
wire n_4101;
wire n_4102;
wire n_4103;
wire n_4104;
wire n_4105;
wire n_4106;
wire n_4107;
wire n_4108;
wire n_4109;
wire n_411;
wire n_4110;
wire n_4111;
wire n_4112;
wire n_4114;
wire n_4115;
wire n_4116;
wire n_4117;
wire n_4118;
wire n_4119;
wire n_412;
wire n_4120;
wire n_4121;
wire n_4122;
wire n_4123;
wire n_4124;
wire n_4126;
wire n_4127;
wire n_4128;
wire n_4129;
wire n_413;
wire n_4130;
wire n_4131;
wire n_4132;
wire n_4133;
wire n_4134;
wire n_4135;
wire n_4136;
wire n_4137;
wire n_4138;
wire n_4139;
wire n_414;
wire n_4140;
wire n_4141;
wire n_4142;
wire n_4143;
wire n_4144;
wire n_4145;
wire n_4146;
wire n_4147;
wire n_4148;
wire n_4149;
wire n_415;
wire n_4150;
wire n_4151;
wire n_4152;
wire n_4153;
wire n_4154;
wire n_4155;
wire n_4156;
wire n_4158;
wire n_4159;
wire n_416;
wire n_4160;
wire n_4161;
wire n_4162;
wire n_4163;
wire n_4164;
wire n_4165;
wire n_4166;
wire n_4167;
wire n_4168;
wire n_4169;
wire n_417;
wire n_4170;
wire n_4171;
wire n_4172;
wire n_4173;
wire n_4174;
wire n_4175;
wire n_4176;
wire n_4177;
wire n_418;
wire n_4180;
wire n_4181;
wire n_4182;
wire n_4183;
wire n_4185;
wire n_4186;
wire n_419;
wire n_4190;
wire n_4192;
wire n_4193;
wire n_4194;
wire n_4195;
wire n_4196;
wire n_4197;
wire n_4198;
wire n_4199;
wire n_42;
wire n_420;
wire n_4201;
wire n_4202;
wire n_4203;
wire n_4204;
wire n_4205;
wire n_4206;
wire n_4207;
wire n_4208;
wire n_4209;
wire n_421;
wire n_4210;
wire n_4211;
wire n_4212;
wire n_4213;
wire n_4214;
wire n_4215;
wire n_4217;
wire n_4218;
wire n_4219;
wire n_422;
wire n_4220;
wire n_4221;
wire n_4222;
wire n_4223;
wire n_4224;
wire n_4225;
wire n_4226;
wire n_4227;
wire n_4228;
wire n_4229;
wire n_423;
wire n_4230;
wire n_4231;
wire n_4232;
wire n_4233;
wire n_4234;
wire n_4235;
wire n_4236;
wire n_4239;
wire n_424;
wire n_4240;
wire n_4241;
wire n_4247;
wire n_4248;
wire n_4249;
wire n_425;
wire n_4250;
wire n_4251;
wire n_4252;
wire n_4253;
wire n_4254;
wire n_4256;
wire n_4257;
wire n_4258;
wire n_4259;
wire n_426;
wire n_4260;
wire n_4262;
wire n_4263;
wire n_4264;
wire n_4265;
wire n_4266;
wire n_4267;
wire n_427;
wire n_4270;
wire n_4276;
wire n_428;
wire n_4280;
wire n_4288;
wire n_4289;
wire n_429;
wire n_4290;
wire n_4291;
wire n_4292;
wire n_4293;
wire n_4294;
wire n_4295;
wire n_4296;
wire n_4297;
wire n_4298;
wire n_4299;
wire n_43;
wire n_430;
wire n_4300;
wire n_4301;
wire n_4302;
wire n_4303;
wire n_4304;
wire n_4305;
wire n_4306;
wire n_4307;
wire n_4308;
wire n_4309;
wire n_431;
wire n_4310;
wire n_4311;
wire n_4312;
wire n_4315;
wire n_4316;
wire n_4317;
wire n_4318;
wire n_4319;
wire n_432;
wire n_4320;
wire n_4322;
wire n_4323;
wire n_4324;
wire n_4325;
wire n_4326;
wire n_4327;
wire n_4328;
wire n_4329;
wire n_433;
wire n_4331;
wire n_4332;
wire n_4334;
wire n_4335;
wire n_4336;
wire n_4337;
wire n_4338;
wire n_434;
wire n_4340;
wire n_4341;
wire n_4342;
wire n_4343;
wire n_4344;
wire n_4345;
wire n_4346;
wire n_4347;
wire n_4349;
wire n_435;
wire n_4350;
wire n_4352;
wire n_4353;
wire n_4354;
wire n_4355;
wire n_4356;
wire n_4357;
wire n_4358;
wire n_4359;
wire n_436;
wire n_4360;
wire n_4362;
wire n_4364;
wire n_4365;
wire n_4366;
wire n_4367;
wire n_4368;
wire n_4369;
wire n_437;
wire n_4370;
wire n_4371;
wire n_4373;
wire n_4374;
wire n_4376;
wire n_4377;
wire n_4378;
wire n_4379;
wire n_438;
wire n_4380;
wire n_4381;
wire n_4382;
wire n_4383;
wire n_4385;
wire n_4386;
wire n_4387;
wire n_4388;
wire n_4389;
wire n_439;
wire n_4390;
wire n_4391;
wire n_4392;
wire n_4393;
wire n_4394;
wire n_4395;
wire n_4396;
wire n_4397;
wire n_4398;
wire n_4399;
wire n_44;
wire n_440;
wire n_4400;
wire n_4401;
wire n_4402;
wire n_4403;
wire n_4404;
wire n_4405;
wire n_4406;
wire n_4407;
wire n_4408;
wire n_4409;
wire n_441;
wire n_4410;
wire n_4411;
wire n_4412;
wire n_4413;
wire n_4414;
wire n_4415;
wire n_4416;
wire n_4417;
wire n_4418;
wire n_4419;
wire n_442;
wire n_4420;
wire n_4421;
wire n_4422;
wire n_4423;
wire n_4424;
wire n_4425;
wire n_4426;
wire n_4427;
wire n_4428;
wire n_4429;
wire n_443;
wire n_4430;
wire n_4431;
wire n_4432;
wire n_4433;
wire n_4434;
wire n_4435;
wire n_4436;
wire n_4437;
wire n_4438;
wire n_4439;
wire n_444;
wire n_4440;
wire n_4441;
wire n_4442;
wire n_4443;
wire n_4444;
wire n_4445;
wire n_4446;
wire n_4447;
wire n_4448;
wire n_4449;
wire n_445;
wire n_4450;
wire n_4451;
wire n_4452;
wire n_4453;
wire n_4454;
wire n_4455;
wire n_4456;
wire n_4457;
wire n_4458;
wire n_4459;
wire n_446;
wire n_4460;
wire n_4461;
wire n_4462;
wire n_4463;
wire n_4464;
wire n_4465;
wire n_4466;
wire n_4467;
wire n_4468;
wire n_4469;
wire n_447;
wire n_4470;
wire n_4471;
wire n_4472;
wire n_4473;
wire n_4474;
wire n_4475;
wire n_4476;
wire n_4477;
wire n_4478;
wire n_4479;
wire n_448;
wire n_4480;
wire n_4481;
wire n_4482;
wire n_4483;
wire n_4484;
wire n_4485;
wire n_4486;
wire n_4487;
wire n_4488;
wire n_4489;
wire n_449;
wire n_4490;
wire n_4491;
wire n_4492;
wire n_4493;
wire n_4494;
wire n_4495;
wire n_4496;
wire n_4497;
wire n_4498;
wire n_4499;
wire n_45;
wire n_450;
wire n_4500;
wire n_4501;
wire n_4502;
wire n_4503;
wire n_4504;
wire n_4505;
wire n_4506;
wire n_4507;
wire n_4508;
wire n_4509;
wire n_451;
wire n_4510;
wire n_4511;
wire n_4512;
wire n_4513;
wire n_4514;
wire n_4515;
wire n_4516;
wire n_4517;
wire n_4518;
wire n_4519;
wire n_452;
wire n_4520;
wire n_4521;
wire n_4522;
wire n_4523;
wire n_4524;
wire n_4525;
wire n_4526;
wire n_4527;
wire n_4528;
wire n_4529;
wire n_453;
wire n_4530;
wire n_4531;
wire n_4532;
wire n_4533;
wire n_4534;
wire n_4535;
wire n_4536;
wire n_4537;
wire n_4538;
wire n_4539;
wire n_454;
wire n_4540;
wire n_4541;
wire n_4542;
wire n_4543;
wire n_4544;
wire n_4545;
wire n_4546;
wire n_4547;
wire n_4548;
wire n_4549;
wire n_455;
wire n_4550;
wire n_4551;
wire n_4552;
wire n_4553;
wire n_4554;
wire n_4555;
wire n_4556;
wire n_4557;
wire n_4558;
wire n_4559;
wire n_456;
wire n_4560;
wire n_4561;
wire n_4562;
wire n_4563;
wire n_4564;
wire n_4565;
wire n_4566;
wire n_4567;
wire n_4568;
wire n_4569;
wire n_457;
wire n_4570;
wire n_4571;
wire n_4572;
wire n_4573;
wire n_4574;
wire n_4575;
wire n_4576;
wire n_4577;
wire n_4578;
wire n_4579;
wire n_458;
wire n_4580;
wire n_4581;
wire n_4582;
wire n_4583;
wire n_4584;
wire n_4585;
wire n_4586;
wire n_4587;
wire n_4588;
wire n_4589;
wire n_459;
wire n_4590;
wire n_4591;
wire n_4592;
wire n_4593;
wire n_4594;
wire n_4595;
wire n_4596;
wire n_4597;
wire n_4598;
wire n_4599;
wire n_46;
wire n_460;
wire n_4600;
wire n_4601;
wire n_4602;
wire n_4603;
wire n_4604;
wire n_4605;
wire n_4606;
wire n_4607;
wire n_4608;
wire n_4609;
wire n_461;
wire n_4610;
wire n_4611;
wire n_4612;
wire n_4613;
wire n_4614;
wire n_4615;
wire n_4616;
wire n_4617;
wire n_4618;
wire n_4619;
wire n_462;
wire n_4620;
wire n_4621;
wire n_4622;
wire n_4623;
wire n_4624;
wire n_4625;
wire n_4626;
wire n_4627;
wire n_4628;
wire n_4629;
wire n_463;
wire n_4630;
wire n_4631;
wire n_4632;
wire n_4633;
wire n_4634;
wire n_4635;
wire n_4636;
wire n_4637;
wire n_4638;
wire n_4639;
wire n_464;
wire n_4640;
wire n_4641;
wire n_4642;
wire n_4643;
wire n_4644;
wire n_4645;
wire n_4646;
wire n_4647;
wire n_4648;
wire n_4649;
wire n_465;
wire n_4650;
wire n_4651;
wire n_4652;
wire n_4653;
wire n_4654;
wire n_4655;
wire n_4656;
wire n_4657;
wire n_4658;
wire n_4659;
wire n_466;
wire n_4660;
wire n_4661;
wire n_4662;
wire n_4663;
wire n_4664;
wire n_4665;
wire n_4666;
wire n_4667;
wire n_4668;
wire n_4669;
wire n_467;
wire n_4670;
wire n_4671;
wire n_4672;
wire n_4673;
wire n_4674;
wire n_4675;
wire n_4676;
wire n_4677;
wire n_4678;
wire n_4679;
wire n_468;
wire n_4680;
wire n_4681;
wire n_4682;
wire n_4683;
wire n_4684;
wire n_4685;
wire n_4686;
wire n_4687;
wire n_4688;
wire n_4689;
wire n_469;
wire n_4690;
wire n_4691;
wire n_4692;
wire n_4693;
wire n_4694;
wire n_4695;
wire n_4696;
wire n_4697;
wire n_4698;
wire n_4699;
wire n_47;
wire n_470;
wire n_4700;
wire n_4701;
wire n_4702;
wire n_4703;
wire n_4704;
wire n_4705;
wire n_4706;
wire n_4707;
wire n_4708;
wire n_4709;
wire n_471;
wire n_4710;
wire n_4711;
wire n_4712;
wire n_4713;
wire n_4714;
wire n_4715;
wire n_4716;
wire n_4717;
wire n_4718;
wire n_4719;
wire n_472;
wire n_4720;
wire n_4722;
wire n_4723;
wire n_4724;
wire n_4725;
wire n_4726;
wire n_4727;
wire n_4728;
wire n_4729;
wire n_473;
wire n_4730;
wire n_4731;
wire n_4732;
wire n_4733;
wire n_4734;
wire n_4735;
wire n_4736;
wire n_4737;
wire n_4738;
wire n_4739;
wire n_474;
wire n_4740;
wire n_4741;
wire n_4742;
wire n_4743;
wire n_4744;
wire n_4745;
wire n_4746;
wire n_4747;
wire n_4748;
wire n_4749;
wire n_475;
wire n_4750;
wire n_4751;
wire n_4752;
wire n_4753;
wire n_4754;
wire n_4755;
wire n_4756;
wire n_4757;
wire n_4758;
wire n_4759;
wire n_476;
wire n_4760;
wire n_4761;
wire n_4762;
wire n_4763;
wire n_4764;
wire n_4765;
wire n_4766;
wire n_4767;
wire n_4768;
wire n_4769;
wire n_477;
wire n_4770;
wire n_4771;
wire n_4772;
wire n_4773;
wire n_4774;
wire n_4775;
wire n_4776;
wire n_4777;
wire n_4778;
wire n_4779;
wire n_478;
wire n_4780;
wire n_4781;
wire n_4782;
wire n_4783;
wire n_4784;
wire n_4785;
wire n_4786;
wire n_4787;
wire n_4788;
wire n_4789;
wire n_479;
wire n_4790;
wire n_4791;
wire n_4793;
wire n_4794;
wire n_4796;
wire n_4797;
wire n_4798;
wire n_4799;
wire n_48;
wire n_480;
wire n_4800;
wire n_4801;
wire n_4802;
wire n_4804;
wire n_4805;
wire n_4806;
wire n_4807;
wire n_4808;
wire n_4809;
wire n_481;
wire n_4810;
wire n_4811;
wire n_4812;
wire n_4813;
wire n_4814;
wire n_4815;
wire n_4816;
wire n_4817;
wire n_4818;
wire n_4819;
wire n_482;
wire n_4820;
wire n_4821;
wire n_4822;
wire n_4823;
wire n_4824;
wire n_4825;
wire n_4826;
wire n_4827;
wire n_4828;
wire n_4829;
wire n_483;
wire n_4830;
wire n_4831;
wire n_4832;
wire n_4833;
wire n_4834;
wire n_4835;
wire n_4836;
wire n_4837;
wire n_4838;
wire n_4839;
wire n_484;
wire n_4840;
wire n_4841;
wire n_4842;
wire n_4843;
wire n_4844;
wire n_4845;
wire n_4846;
wire n_4847;
wire n_4848;
wire n_4849;
wire n_485;
wire n_4850;
wire n_4851;
wire n_4852;
wire n_4853;
wire n_4854;
wire n_4855;
wire n_4856;
wire n_4857;
wire n_4858;
wire n_4859;
wire n_486;
wire n_4860;
wire n_4861;
wire n_4862;
wire n_4863;
wire n_4864;
wire n_4865;
wire n_4866;
wire n_4867;
wire n_4868;
wire n_4869;
wire n_487;
wire n_4870;
wire n_4871;
wire n_4872;
wire n_4873;
wire n_4874;
wire n_4876;
wire n_4878;
wire n_4879;
wire n_488;
wire n_4880;
wire n_4881;
wire n_4882;
wire n_4883;
wire n_4884;
wire n_4885;
wire n_4886;
wire n_4887;
wire n_4888;
wire n_4889;
wire n_489;
wire n_4890;
wire n_4891;
wire n_4892;
wire n_4893;
wire n_4894;
wire n_4895;
wire n_4896;
wire n_4898;
wire n_4899;
wire n_49;
wire n_490;
wire n_4900;
wire n_4901;
wire n_4902;
wire n_4903;
wire n_4905;
wire n_4906;
wire n_4907;
wire n_4908;
wire n_4909;
wire n_491;
wire n_4911;
wire n_4912;
wire n_4913;
wire n_4914;
wire n_4915;
wire n_4916;
wire n_4917;
wire n_4918;
wire n_4919;
wire n_492;
wire n_4920;
wire n_4921;
wire n_4922;
wire n_4923;
wire n_4924;
wire n_4925;
wire n_4927;
wire n_4928;
wire n_4929;
wire n_493;
wire n_4931;
wire n_4932;
wire n_4933;
wire n_4934;
wire n_4935;
wire n_4936;
wire n_4937;
wire n_4938;
wire n_4939;
wire n_494;
wire n_4940;
wire n_4941;
wire n_4942;
wire n_4943;
wire n_4944;
wire n_4945;
wire n_4946;
wire n_4947;
wire n_4948;
wire n_4949;
wire n_495;
wire n_4950;
wire n_4951;
wire n_4952;
wire n_4953;
wire n_4954;
wire n_4955;
wire n_4956;
wire n_4957;
wire n_4958;
wire n_4959;
wire n_496;
wire n_4960;
wire n_4961;
wire n_4962;
wire n_4963;
wire n_4964;
wire n_4965;
wire n_4966;
wire n_4967;
wire n_4968;
wire n_4969;
wire n_497;
wire n_4970;
wire n_4971;
wire n_4972;
wire n_4973;
wire n_4974;
wire n_4975;
wire n_4976;
wire n_4977;
wire n_4978;
wire n_4979;
wire n_498;
wire n_4980;
wire n_4981;
wire n_4982;
wire n_4983;
wire n_4984;
wire n_4985;
wire n_4986;
wire n_4987;
wire n_4988;
wire n_4989;
wire n_499;
wire n_4990;
wire n_4991;
wire n_4992;
wire n_4993;
wire n_4994;
wire n_4995;
wire n_4996;
wire n_4997;
wire n_4998;
wire n_4999;
wire n_5;
wire n_50;
wire n_500;
wire n_5000;
wire n_5001;
wire n_5003;
wire n_5006;
wire n_501;
wire n_502;
wire n_5022;
wire n_5023;
wire n_5024;
wire n_5025;
wire n_5026;
wire n_5027;
wire n_5028;
wire n_503;
wire n_5031;
wire n_5032;
wire n_5034;
wire n_5035;
wire n_5036;
wire n_5038;
wire n_5039;
wire n_504;
wire n_5041;
wire n_5042;
wire n_5043;
wire n_5045;
wire n_5046;
wire n_5048;
wire n_5049;
wire n_505;
wire n_5050;
wire n_5054;
wire n_5055;
wire n_5056;
wire n_5057;
wire n_506;
wire n_5062;
wire n_5063;
wire n_5064;
wire n_5065;
wire n_5067;
wire n_5068;
wire n_5069;
wire n_507;
wire n_5071;
wire n_5072;
wire n_5073;
wire n_5074;
wire n_5075;
wire n_5076;
wire n_5078;
wire n_5079;
wire n_508;
wire n_5080;
wire n_5081;
wire n_5084;
wire n_5085;
wire n_5087;
wire n_5088;
wire n_5089;
wire n_509;
wire n_5090;
wire n_5091;
wire n_5092;
wire n_5093;
wire n_5094;
wire n_5095;
wire n_5096;
wire n_5097;
wire n_5098;
wire n_5099;
wire n_51;
wire n_510;
wire n_5100;
wire n_5101;
wire n_5102;
wire n_5103;
wire n_5104;
wire n_5105;
wire n_5106;
wire n_5107;
wire n_5108;
wire n_5109;
wire n_511;
wire n_5110;
wire n_5111;
wire n_5112;
wire n_5113;
wire n_5114;
wire n_5115;
wire n_5116;
wire n_5117;
wire n_5118;
wire n_5119;
wire n_512;
wire n_5120;
wire n_5121;
wire n_5122;
wire n_5123;
wire n_5124;
wire n_5125;
wire n_5126;
wire n_5127;
wire n_5128;
wire n_5129;
wire n_513;
wire n_5130;
wire n_5131;
wire n_5132;
wire n_5133;
wire n_5134;
wire n_5135;
wire n_5136;
wire n_5137;
wire n_5138;
wire n_5139;
wire n_514;
wire n_5140;
wire n_5141;
wire n_5142;
wire n_5143;
wire n_5144;
wire n_5145;
wire n_5146;
wire n_5147;
wire n_5148;
wire n_5149;
wire n_515;
wire n_5150;
wire n_5151;
wire n_5152;
wire n_5153;
wire n_5154;
wire n_5156;
wire n_5157;
wire n_5158;
wire n_5159;
wire n_516;
wire n_5160;
wire n_5161;
wire n_5162;
wire n_5163;
wire n_5164;
wire n_5165;
wire n_5166;
wire n_5167;
wire n_5168;
wire n_5169;
wire n_517;
wire n_5170;
wire n_5171;
wire n_5172;
wire n_5173;
wire n_5174;
wire n_5175;
wire n_5176;
wire n_5177;
wire n_5178;
wire n_5179;
wire n_518;
wire n_5180;
wire n_5181;
wire n_5182;
wire n_5183;
wire n_5185;
wire n_5186;
wire n_5187;
wire n_5188;
wire n_5189;
wire n_519;
wire n_5190;
wire n_5191;
wire n_5192;
wire n_5193;
wire n_5194;
wire n_5195;
wire n_5196;
wire n_5197;
wire n_5198;
wire n_5199;
wire n_52;
wire n_520;
wire n_5200;
wire n_5201;
wire n_5202;
wire n_5203;
wire n_5204;
wire n_5205;
wire n_5206;
wire n_5207;
wire n_5208;
wire n_5209;
wire n_521;
wire n_5210;
wire n_5211;
wire n_5212;
wire n_5213;
wire n_5214;
wire n_5215;
wire n_5216;
wire n_5217;
wire n_5218;
wire n_5219;
wire n_522;
wire n_5220;
wire n_5221;
wire n_5222;
wire n_5223;
wire n_5224;
wire n_5225;
wire n_5226;
wire n_5227;
wire n_5228;
wire n_5229;
wire n_523;
wire n_5230;
wire n_5231;
wire n_5232;
wire n_5233;
wire n_5234;
wire n_5235;
wire n_5236;
wire n_5237;
wire n_5238;
wire n_5239;
wire n_524;
wire n_5240;
wire n_5241;
wire n_5242;
wire n_5243;
wire n_5244;
wire n_5245;
wire n_5246;
wire n_5247;
wire n_5248;
wire n_5249;
wire n_525;
wire n_5250;
wire n_5251;
wire n_5252;
wire n_5253;
wire n_5254;
wire n_5255;
wire n_5256;
wire n_5257;
wire n_5258;
wire n_5259;
wire n_526;
wire n_5260;
wire n_5261;
wire n_5262;
wire n_5263;
wire n_5264;
wire n_5265;
wire n_5266;
wire n_5267;
wire n_5268;
wire n_5269;
wire n_527;
wire n_5270;
wire n_5271;
wire n_5272;
wire n_5273;
wire n_5274;
wire n_5275;
wire n_5276;
wire n_5277;
wire n_5278;
wire n_5279;
wire n_528;
wire n_5280;
wire n_5281;
wire n_5282;
wire n_5283;
wire n_5284;
wire n_5285;
wire n_5286;
wire n_5287;
wire n_5288;
wire n_5289;
wire n_529;
wire n_5290;
wire n_5291;
wire n_5292;
wire n_5293;
wire n_5294;
wire n_5295;
wire n_5296;
wire n_5297;
wire n_5298;
wire n_5299;
wire n_53;
wire n_530;
wire n_5300;
wire n_5301;
wire n_5302;
wire n_5303;
wire n_5304;
wire n_5305;
wire n_5306;
wire n_5307;
wire n_5308;
wire n_5309;
wire n_531;
wire n_5310;
wire n_5311;
wire n_5312;
wire n_5313;
wire n_5314;
wire n_5315;
wire n_5316;
wire n_5317;
wire n_5318;
wire n_5319;
wire n_532;
wire n_5320;
wire n_5321;
wire n_5322;
wire n_5323;
wire n_5324;
wire n_5325;
wire n_5326;
wire n_5327;
wire n_5328;
wire n_5329;
wire n_533;
wire n_5330;
wire n_5331;
wire n_5332;
wire n_5333;
wire n_5334;
wire n_5335;
wire n_5336;
wire n_5337;
wire n_5338;
wire n_5339;
wire n_534;
wire n_5340;
wire n_5341;
wire n_5342;
wire n_5343;
wire n_5344;
wire n_5345;
wire n_5346;
wire n_5347;
wire n_5348;
wire n_5349;
wire n_535;
wire n_5350;
wire n_5351;
wire n_5352;
wire n_5353;
wire n_5354;
wire n_5355;
wire n_5356;
wire n_5357;
wire n_5358;
wire n_5359;
wire n_536;
wire n_5360;
wire n_5361;
wire n_5362;
wire n_5363;
wire n_5364;
wire n_5365;
wire n_5366;
wire n_5367;
wire n_5368;
wire n_5369;
wire n_537;
wire n_5370;
wire n_5371;
wire n_5372;
wire n_5373;
wire n_5374;
wire n_5375;
wire n_5376;
wire n_5377;
wire n_5378;
wire n_538;
wire n_5380;
wire n_5381;
wire n_5382;
wire n_5383;
wire n_5384;
wire n_5385;
wire n_5386;
wire n_5387;
wire n_5388;
wire n_5389;
wire n_539;
wire n_5390;
wire n_5391;
wire n_5392;
wire n_5393;
wire n_5394;
wire n_5395;
wire n_5396;
wire n_5397;
wire n_5398;
wire n_5399;
wire n_54;
wire n_540;
wire n_5400;
wire n_5401;
wire n_5402;
wire n_5403;
wire n_5404;
wire n_5405;
wire n_5406;
wire n_5407;
wire n_5408;
wire n_5409;
wire n_541;
wire n_5410;
wire n_5411;
wire n_5412;
wire n_5414;
wire n_5415;
wire n_5416;
wire n_5417;
wire n_5418;
wire n_5419;
wire n_542;
wire n_5420;
wire n_5421;
wire n_5422;
wire n_5423;
wire n_5424;
wire n_5425;
wire n_5426;
wire n_5427;
wire n_5428;
wire n_5429;
wire n_543;
wire n_5430;
wire n_5431;
wire n_5432;
wire n_5433;
wire n_5434;
wire n_5435;
wire n_5436;
wire n_5437;
wire n_5438;
wire n_5439;
wire n_544;
wire n_5440;
wire n_5441;
wire n_5442;
wire n_5443;
wire n_5444;
wire n_5445;
wire n_5446;
wire n_5447;
wire n_5448;
wire n_5449;
wire n_545;
wire n_5450;
wire n_5451;
wire n_5452;
wire n_5453;
wire n_5454;
wire n_5455;
wire n_5456;
wire n_5457;
wire n_5458;
wire n_5459;
wire n_546;
wire n_5460;
wire n_5461;
wire n_5462;
wire n_5463;
wire n_5464;
wire n_5465;
wire n_5466;
wire n_5467;
wire n_5468;
wire n_5469;
wire n_547;
wire n_5470;
wire n_5471;
wire n_5472;
wire n_5473;
wire n_5474;
wire n_5475;
wire n_5476;
wire n_5477;
wire n_5478;
wire n_5479;
wire n_548;
wire n_5480;
wire n_5481;
wire n_5482;
wire n_5483;
wire n_5484;
wire n_5485;
wire n_5486;
wire n_5487;
wire n_5488;
wire n_5489;
wire n_549;
wire n_5490;
wire n_5491;
wire n_5492;
wire n_5493;
wire n_5494;
wire n_5495;
wire n_5496;
wire n_5497;
wire n_5498;
wire n_5499;
wire n_55;
wire n_550;
wire n_5500;
wire n_5501;
wire n_5502;
wire n_5503;
wire n_5504;
wire n_5505;
wire n_5506;
wire n_5507;
wire n_5508;
wire n_5509;
wire n_551;
wire n_5510;
wire n_5511;
wire n_5512;
wire n_5513;
wire n_5514;
wire n_5515;
wire n_5516;
wire n_5517;
wire n_5518;
wire n_5519;
wire n_552;
wire n_5520;
wire n_5521;
wire n_5522;
wire n_5523;
wire n_5524;
wire n_5525;
wire n_5526;
wire n_5527;
wire n_5528;
wire n_5529;
wire n_553;
wire n_5530;
wire n_5531;
wire n_5532;
wire n_5533;
wire n_5534;
wire n_5535;
wire n_5536;
wire n_5537;
wire n_5538;
wire n_5539;
wire n_554;
wire n_5540;
wire n_5541;
wire n_5542;
wire n_5543;
wire n_5544;
wire n_5545;
wire n_5546;
wire n_5547;
wire n_5548;
wire n_5549;
wire n_555;
wire n_5550;
wire n_5551;
wire n_5552;
wire n_5553;
wire n_5554;
wire n_5555;
wire n_5556;
wire n_5557;
wire n_5558;
wire n_5559;
wire n_556;
wire n_5560;
wire n_5561;
wire n_5562;
wire n_5563;
wire n_5564;
wire n_5565;
wire n_5566;
wire n_5567;
wire n_5568;
wire n_5569;
wire n_557;
wire n_5570;
wire n_5571;
wire n_5572;
wire n_5573;
wire n_5574;
wire n_5575;
wire n_5576;
wire n_5577;
wire n_5578;
wire n_5579;
wire n_558;
wire n_5580;
wire n_5581;
wire n_5582;
wire n_5583;
wire n_5584;
wire n_5585;
wire n_5586;
wire n_5587;
wire n_5588;
wire n_5589;
wire n_559;
wire n_5590;
wire n_5591;
wire n_5592;
wire n_5593;
wire n_5594;
wire n_5595;
wire n_5596;
wire n_5597;
wire n_5598;
wire n_56;
wire n_560;
wire n_5600;
wire n_5601;
wire n_5602;
wire n_5603;
wire n_5604;
wire n_5605;
wire n_5606;
wire n_5607;
wire n_5608;
wire n_5609;
wire n_561;
wire n_5610;
wire n_5611;
wire n_5612;
wire n_5613;
wire n_5614;
wire n_5615;
wire n_5616;
wire n_5617;
wire n_5618;
wire n_5619;
wire n_562;
wire n_5620;
wire n_5621;
wire n_5622;
wire n_5623;
wire n_5624;
wire n_5625;
wire n_5626;
wire n_5627;
wire n_5628;
wire n_5629;
wire n_563;
wire n_5630;
wire n_5631;
wire n_5632;
wire n_5633;
wire n_5634;
wire n_5635;
wire n_5636;
wire n_5637;
wire n_5638;
wire n_5639;
wire n_564;
wire n_5640;
wire n_5641;
wire n_5642;
wire n_5643;
wire n_5644;
wire n_5645;
wire n_5646;
wire n_5647;
wire n_5648;
wire n_5649;
wire n_565;
wire n_5650;
wire n_5651;
wire n_5652;
wire n_5653;
wire n_5654;
wire n_5655;
wire n_5656;
wire n_5657;
wire n_5658;
wire n_5659;
wire n_566;
wire n_5660;
wire n_5661;
wire n_5662;
wire n_5663;
wire n_5664;
wire n_5665;
wire n_5666;
wire n_5667;
wire n_5668;
wire n_5669;
wire n_567;
wire n_5670;
wire n_5671;
wire n_5672;
wire n_5673;
wire n_5674;
wire n_5675;
wire n_5676;
wire n_5677;
wire n_5678;
wire n_5679;
wire n_568;
wire n_5680;
wire n_5681;
wire n_5682;
wire n_5683;
wire n_5684;
wire n_5685;
wire n_5686;
wire n_5687;
wire n_5688;
wire n_5689;
wire n_569;
wire n_5690;
wire n_5691;
wire n_5692;
wire n_5693;
wire n_5694;
wire n_5695;
wire n_5696;
wire n_5697;
wire n_5698;
wire n_5699;
wire n_57;
wire n_570;
wire n_5700;
wire n_5701;
wire n_5702;
wire n_5703;
wire n_5704;
wire n_5705;
wire n_5706;
wire n_5707;
wire n_5708;
wire n_5709;
wire n_571;
wire n_5710;
wire n_5711;
wire n_5712;
wire n_5713;
wire n_5714;
wire n_5715;
wire n_5716;
wire n_5717;
wire n_5718;
wire n_5719;
wire n_572;
wire n_5720;
wire n_5721;
wire n_5722;
wire n_5723;
wire n_5724;
wire n_5725;
wire n_5726;
wire n_5727;
wire n_5728;
wire n_5729;
wire n_573;
wire n_5730;
wire n_5731;
wire n_5732;
wire n_5733;
wire n_5734;
wire n_5735;
wire n_5736;
wire n_5737;
wire n_5738;
wire n_5739;
wire n_574;
wire n_5740;
wire n_5741;
wire n_5742;
wire n_5743;
wire n_5744;
wire n_5745;
wire n_5746;
wire n_5747;
wire n_5748;
wire n_5749;
wire n_575;
wire n_5750;
wire n_5751;
wire n_5752;
wire n_5753;
wire n_5754;
wire n_5755;
wire n_5756;
wire n_5757;
wire n_5758;
wire n_5759;
wire n_576;
wire n_5760;
wire n_5761;
wire n_5762;
wire n_5763;
wire n_5764;
wire n_5765;
wire n_5766;
wire n_5767;
wire n_5768;
wire n_5769;
wire n_577;
wire n_5770;
wire n_5771;
wire n_5772;
wire n_5773;
wire n_5774;
wire n_5775;
wire n_5776;
wire n_5777;
wire n_5778;
wire n_5779;
wire n_578;
wire n_5780;
wire n_5781;
wire n_5782;
wire n_5783;
wire n_5784;
wire n_5785;
wire n_5786;
wire n_5787;
wire n_5788;
wire n_5789;
wire n_579;
wire n_5790;
wire n_5791;
wire n_5792;
wire n_5793;
wire n_5794;
wire n_5795;
wire n_5796;
wire n_5797;
wire n_5798;
wire n_5799;
wire n_58;
wire n_580;
wire n_5800;
wire n_5801;
wire n_5802;
wire n_5803;
wire n_5804;
wire n_5805;
wire n_5806;
wire n_5807;
wire n_5808;
wire n_5809;
wire n_581;
wire n_5810;
wire n_5811;
wire n_5812;
wire n_5813;
wire n_5814;
wire n_5815;
wire n_5816;
wire n_5817;
wire n_5818;
wire n_5819;
wire n_582;
wire n_5820;
wire n_5821;
wire n_5822;
wire n_5823;
wire n_5824;
wire n_5825;
wire n_5826;
wire n_5827;
wire n_5828;
wire n_5829;
wire n_583;
wire n_5830;
wire n_5831;
wire n_5832;
wire n_5833;
wire n_5834;
wire n_5835;
wire n_5836;
wire n_5837;
wire n_5838;
wire n_5839;
wire n_584;
wire n_5840;
wire n_5841;
wire n_5842;
wire n_5843;
wire n_5844;
wire n_5845;
wire n_5846;
wire n_5847;
wire n_5848;
wire n_5849;
wire n_585;
wire n_5850;
wire n_5851;
wire n_5852;
wire n_5853;
wire n_5854;
wire n_5855;
wire n_5856;
wire n_5857;
wire n_5858;
wire n_5859;
wire n_586;
wire n_5860;
wire n_5861;
wire n_5862;
wire n_5863;
wire n_5864;
wire n_5865;
wire n_5866;
wire n_5867;
wire n_5868;
wire n_5869;
wire n_587;
wire n_5870;
wire n_5871;
wire n_5872;
wire n_5873;
wire n_5874;
wire n_5875;
wire n_5876;
wire n_5877;
wire n_5878;
wire n_5879;
wire n_588;
wire n_5880;
wire n_5881;
wire n_5882;
wire n_5883;
wire n_5884;
wire n_5885;
wire n_5886;
wire n_5887;
wire n_5888;
wire n_5889;
wire n_589;
wire n_5890;
wire n_5891;
wire n_5892;
wire n_5893;
wire n_5894;
wire n_5895;
wire n_5896;
wire n_5897;
wire n_5898;
wire n_5899;
wire n_59;
wire n_590;
wire n_5900;
wire n_5901;
wire n_5902;
wire n_5903;
wire n_5904;
wire n_5905;
wire n_5906;
wire n_5907;
wire n_5908;
wire n_5909;
wire n_591;
wire n_5910;
wire n_5911;
wire n_5912;
wire n_5913;
wire n_5914;
wire n_5915;
wire n_5916;
wire n_5917;
wire n_5918;
wire n_5919;
wire n_592;
wire n_5920;
wire n_5921;
wire n_5922;
wire n_5923;
wire n_5924;
wire n_5925;
wire n_5926;
wire n_5927;
wire n_5928;
wire n_5929;
wire n_593;
wire n_5930;
wire n_5931;
wire n_5932;
wire n_5933;
wire n_5934;
wire n_5935;
wire n_5936;
wire n_5937;
wire n_5938;
wire n_5939;
wire n_594;
wire n_5940;
wire n_5941;
wire n_5942;
wire n_5943;
wire n_5944;
wire n_5945;
wire n_5946;
wire n_5947;
wire n_5948;
wire n_5949;
wire n_595;
wire n_5950;
wire n_5951;
wire n_5952;
wire n_5953;
wire n_5954;
wire n_5955;
wire n_5956;
wire n_5957;
wire n_5958;
wire n_5959;
wire n_596;
wire n_5960;
wire n_5961;
wire n_5962;
wire n_5963;
wire n_5964;
wire n_5965;
wire n_5966;
wire n_5967;
wire n_5968;
wire n_5969;
wire n_597;
wire n_5970;
wire n_5971;
wire n_5972;
wire n_5973;
wire n_5974;
wire n_5975;
wire n_5976;
wire n_5977;
wire n_5978;
wire n_5979;
wire n_598;
wire n_5980;
wire n_5981;
wire n_5983;
wire n_5984;
wire n_5985;
wire n_5986;
wire n_5987;
wire n_5988;
wire n_5989;
wire n_599;
wire n_5990;
wire n_5991;
wire n_5992;
wire n_5993;
wire n_5994;
wire n_5995;
wire n_5996;
wire n_5997;
wire n_5998;
wire n_5999;
wire n_6;
wire n_60;
wire n_600;
wire n_6000;
wire n_6001;
wire n_6002;
wire n_6003;
wire n_6004;
wire n_6005;
wire n_6006;
wire n_6007;
wire n_6008;
wire n_6009;
wire n_601;
wire n_6010;
wire n_6011;
wire n_6012;
wire n_6013;
wire n_6014;
wire n_6015;
wire n_6016;
wire n_6017;
wire n_6018;
wire n_6019;
wire n_602;
wire n_6020;
wire n_6021;
wire n_6022;
wire n_6023;
wire n_6024;
wire n_6025;
wire n_6026;
wire n_6027;
wire n_6028;
wire n_6029;
wire n_603;
wire n_6030;
wire n_6031;
wire n_6032;
wire n_6033;
wire n_6034;
wire n_6035;
wire n_6036;
wire n_6037;
wire n_6038;
wire n_604;
wire n_6040;
wire n_6041;
wire n_6042;
wire n_6043;
wire n_6044;
wire n_6045;
wire n_6046;
wire n_6047;
wire n_6048;
wire n_6049;
wire n_605;
wire n_6050;
wire n_6051;
wire n_6052;
wire n_6053;
wire n_6054;
wire n_6055;
wire n_6056;
wire n_6057;
wire n_6058;
wire n_6059;
wire n_606;
wire n_6060;
wire n_6061;
wire n_6062;
wire n_6063;
wire n_6064;
wire n_6065;
wire n_6066;
wire n_6067;
wire n_6068;
wire n_6069;
wire n_607;
wire n_6070;
wire n_6071;
wire n_6072;
wire n_6073;
wire n_6074;
wire n_6075;
wire n_6076;
wire n_6077;
wire n_6078;
wire n_6079;
wire n_608;
wire n_6080;
wire n_6081;
wire n_6082;
wire n_6083;
wire n_6084;
wire n_6085;
wire n_6086;
wire n_6087;
wire n_6088;
wire n_6089;
wire n_609;
wire n_6090;
wire n_6091;
wire n_6092;
wire n_6093;
wire n_6094;
wire n_6095;
wire n_6096;
wire n_6097;
wire n_6098;
wire n_6099;
wire n_61;
wire n_610;
wire n_6100;
wire n_6101;
wire n_6102;
wire n_6103;
wire n_6104;
wire n_6105;
wire n_6106;
wire n_6107;
wire n_6108;
wire n_6109;
wire n_611;
wire n_6110;
wire n_6111;
wire n_6112;
wire n_6113;
wire n_6114;
wire n_6115;
wire n_6116;
wire n_6117;
wire n_6118;
wire n_6119;
wire n_612;
wire n_6120;
wire n_6121;
wire n_6122;
wire n_6123;
wire n_6124;
wire n_6125;
wire n_6126;
wire n_6127;
wire n_6128;
wire n_6129;
wire n_613;
wire n_6130;
wire n_6131;
wire n_6132;
wire n_6133;
wire n_6134;
wire n_6135;
wire n_6136;
wire n_6137;
wire n_6138;
wire n_6139;
wire n_614;
wire n_6140;
wire n_6141;
wire n_6142;
wire n_6143;
wire n_6144;
wire n_6145;
wire n_6146;
wire n_6147;
wire n_6148;
wire n_6149;
wire n_615;
wire n_6150;
wire n_6151;
wire n_6152;
wire n_6153;
wire n_6154;
wire n_6155;
wire n_6156;
wire n_6157;
wire n_6158;
wire n_6159;
wire n_616;
wire n_6160;
wire n_6161;
wire n_6162;
wire n_6163;
wire n_6164;
wire n_6165;
wire n_6166;
wire n_6167;
wire n_6168;
wire n_6169;
wire n_617;
wire n_6170;
wire n_6171;
wire n_6172;
wire n_6173;
wire n_6174;
wire n_6175;
wire n_6176;
wire n_6177;
wire n_6178;
wire n_6179;
wire n_618;
wire n_6180;
wire n_6181;
wire n_6182;
wire n_6183;
wire n_6184;
wire n_6185;
wire n_6186;
wire n_6187;
wire n_6188;
wire n_6189;
wire n_619;
wire n_6190;
wire n_6191;
wire n_6192;
wire n_6193;
wire n_6194;
wire n_6195;
wire n_6196;
wire n_6197;
wire n_6198;
wire n_6199;
wire n_62;
wire n_620;
wire n_6200;
wire n_6201;
wire n_6202;
wire n_6203;
wire n_6204;
wire n_6205;
wire n_6206;
wire n_6207;
wire n_6208;
wire n_6209;
wire n_621;
wire n_6210;
wire n_6211;
wire n_6212;
wire n_6213;
wire n_6214;
wire n_6215;
wire n_6216;
wire n_6217;
wire n_6218;
wire n_6219;
wire n_622;
wire n_6220;
wire n_6221;
wire n_6222;
wire n_6223;
wire n_6224;
wire n_6225;
wire n_6226;
wire n_6227;
wire n_6228;
wire n_6229;
wire n_623;
wire n_6230;
wire n_6231;
wire n_6232;
wire n_6233;
wire n_6234;
wire n_6235;
wire n_6236;
wire n_6237;
wire n_6238;
wire n_6239;
wire n_624;
wire n_6240;
wire n_6241;
wire n_6242;
wire n_6243;
wire n_6244;
wire n_6245;
wire n_6246;
wire n_6247;
wire n_6248;
wire n_6249;
wire n_625;
wire n_6250;
wire n_6251;
wire n_6252;
wire n_6253;
wire n_6254;
wire n_6255;
wire n_6256;
wire n_6257;
wire n_6258;
wire n_6259;
wire n_626;
wire n_6260;
wire n_6261;
wire n_6262;
wire n_6263;
wire n_6264;
wire n_6265;
wire n_6266;
wire n_6267;
wire n_6268;
wire n_6269;
wire n_627;
wire n_6270;
wire n_6271;
wire n_6272;
wire n_6273;
wire n_6274;
wire n_6275;
wire n_6276;
wire n_6277;
wire n_6278;
wire n_6279;
wire n_628;
wire n_6280;
wire n_6281;
wire n_6282;
wire n_6283;
wire n_6284;
wire n_6285;
wire n_6286;
wire n_6287;
wire n_6288;
wire n_6289;
wire n_629;
wire n_6290;
wire n_6291;
wire n_6292;
wire n_6293;
wire n_6294;
wire n_6295;
wire n_6296;
wire n_6297;
wire n_6298;
wire n_6299;
wire n_63;
wire n_630;
wire n_6300;
wire n_6301;
wire n_6302;
wire n_6303;
wire n_6304;
wire n_6305;
wire n_6306;
wire n_6307;
wire n_6308;
wire n_6309;
wire n_631;
wire n_6310;
wire n_6311;
wire n_6312;
wire n_6313;
wire n_6314;
wire n_6315;
wire n_6316;
wire n_6317;
wire n_6318;
wire n_6319;
wire n_632;
wire n_6320;
wire n_6321;
wire n_6322;
wire n_6323;
wire n_6324;
wire n_6325;
wire n_6326;
wire n_6327;
wire n_6328;
wire n_6329;
wire n_633;
wire n_6330;
wire n_6331;
wire n_6332;
wire n_6333;
wire n_6334;
wire n_6335;
wire n_6336;
wire n_6337;
wire n_6338;
wire n_6339;
wire n_634;
wire n_6340;
wire n_6341;
wire n_6342;
wire n_6343;
wire n_6344;
wire n_6345;
wire n_6346;
wire n_6347;
wire n_6348;
wire n_6349;
wire n_635;
wire n_6350;
wire n_6351;
wire n_6352;
wire n_6353;
wire n_6354;
wire n_6355;
wire n_6356;
wire n_6357;
wire n_6358;
wire n_6359;
wire n_636;
wire n_6360;
wire n_6361;
wire n_6362;
wire n_6363;
wire n_6364;
wire n_6365;
wire n_6366;
wire n_6367;
wire n_6368;
wire n_6369;
wire n_637;
wire n_6370;
wire n_6371;
wire n_6372;
wire n_6373;
wire n_6374;
wire n_6375;
wire n_6376;
wire n_6377;
wire n_6378;
wire n_6379;
wire n_638;
wire n_6380;
wire n_6381;
wire n_6382;
wire n_6383;
wire n_6384;
wire n_6385;
wire n_6386;
wire n_6387;
wire n_6388;
wire n_6389;
wire n_639;
wire n_6390;
wire n_6391;
wire n_6392;
wire n_6393;
wire n_6394;
wire n_6395;
wire n_6396;
wire n_6397;
wire n_6398;
wire n_6399;
wire n_64;
wire n_640;
wire n_6400;
wire n_6401;
wire n_6402;
wire n_6403;
wire n_6404;
wire n_6405;
wire n_6406;
wire n_6407;
wire n_6408;
wire n_6409;
wire n_641;
wire n_6410;
wire n_6411;
wire n_6412;
wire n_6413;
wire n_6414;
wire n_6415;
wire n_6416;
wire n_6417;
wire n_6418;
wire n_6419;
wire n_642;
wire n_6420;
wire n_6421;
wire n_6422;
wire n_6423;
wire n_6424;
wire n_6425;
wire n_6426;
wire n_6427;
wire n_6428;
wire n_6429;
wire n_643;
wire n_6430;
wire n_6431;
wire n_6432;
wire n_6433;
wire n_6434;
wire n_6435;
wire n_6436;
wire n_6437;
wire n_6438;
wire n_6439;
wire n_644;
wire n_6440;
wire n_6441;
wire n_6442;
wire n_6443;
wire n_6444;
wire n_6445;
wire n_6446;
wire n_6447;
wire n_6448;
wire n_6449;
wire n_645;
wire n_6450;
wire n_6451;
wire n_6452;
wire n_6453;
wire n_6454;
wire n_6455;
wire n_6456;
wire n_6457;
wire n_6458;
wire n_6459;
wire n_646;
wire n_6460;
wire n_6461;
wire n_6462;
wire n_6463;
wire n_6464;
wire n_6465;
wire n_6466;
wire n_6467;
wire n_6468;
wire n_6469;
wire n_647;
wire n_6470;
wire n_6471;
wire n_6472;
wire n_6473;
wire n_6474;
wire n_6475;
wire n_6476;
wire n_6477;
wire n_6478;
wire n_6479;
wire n_648;
wire n_6480;
wire n_6481;
wire n_6482;
wire n_6483;
wire n_6484;
wire n_6485;
wire n_6486;
wire n_6487;
wire n_6488;
wire n_6489;
wire n_649;
wire n_6490;
wire n_6491;
wire n_6492;
wire n_6493;
wire n_6494;
wire n_6495;
wire n_6496;
wire n_6497;
wire n_6498;
wire n_6499;
wire n_65;
wire n_650;
wire n_6500;
wire n_6501;
wire n_6502;
wire n_6503;
wire n_6504;
wire n_6505;
wire n_6506;
wire n_6507;
wire n_6508;
wire n_6509;
wire n_651;
wire n_6510;
wire n_6511;
wire n_6512;
wire n_6513;
wire n_6514;
wire n_6515;
wire n_6516;
wire n_6517;
wire n_6518;
wire n_6519;
wire n_652;
wire n_6520;
wire n_6521;
wire n_6522;
wire n_6523;
wire n_6524;
wire n_6525;
wire n_6526;
wire n_6527;
wire n_6528;
wire n_6529;
wire n_653;
wire n_6530;
wire n_6531;
wire n_6532;
wire n_6533;
wire n_6534;
wire n_6535;
wire n_6536;
wire n_6537;
wire n_6538;
wire n_6539;
wire n_654;
wire n_6540;
wire n_6541;
wire n_6542;
wire n_6543;
wire n_6544;
wire n_6545;
wire n_6546;
wire n_6547;
wire n_6548;
wire n_6549;
wire n_655;
wire n_6550;
wire n_6551;
wire n_6552;
wire n_6553;
wire n_6554;
wire n_6555;
wire n_6556;
wire n_6557;
wire n_6558;
wire n_6559;
wire n_656;
wire n_6560;
wire n_6561;
wire n_6562;
wire n_6563;
wire n_6564;
wire n_6565;
wire n_6566;
wire n_6567;
wire n_6568;
wire n_6569;
wire n_657;
wire n_6570;
wire n_6571;
wire n_6572;
wire n_6573;
wire n_6574;
wire n_6575;
wire n_6576;
wire n_6577;
wire n_6578;
wire n_6579;
wire n_658;
wire n_6580;
wire n_6581;
wire n_6582;
wire n_6583;
wire n_6584;
wire n_6585;
wire n_6586;
wire n_6587;
wire n_6588;
wire n_6589;
wire n_659;
wire n_6590;
wire n_6591;
wire n_6592;
wire n_6593;
wire n_6594;
wire n_6595;
wire n_6596;
wire n_6597;
wire n_6598;
wire n_6599;
wire n_66;
wire n_660;
wire n_6600;
wire n_6601;
wire n_6602;
wire n_6603;
wire n_6604;
wire n_6605;
wire n_6606;
wire n_6607;
wire n_6608;
wire n_6609;
wire n_661;
wire n_6610;
wire n_6611;
wire n_6612;
wire n_6613;
wire n_6614;
wire n_6615;
wire n_6616;
wire n_6617;
wire n_6618;
wire n_6619;
wire n_662;
wire n_6620;
wire n_6621;
wire n_6622;
wire n_6623;
wire n_6624;
wire n_6625;
wire n_6626;
wire n_6627;
wire n_6628;
wire n_6629;
wire n_663;
wire n_6630;
wire n_6631;
wire n_6632;
wire n_6633;
wire n_6634;
wire n_6635;
wire n_6636;
wire n_6637;
wire n_6638;
wire n_6639;
wire n_664;
wire n_6640;
wire n_6641;
wire n_6642;
wire n_6643;
wire n_6644;
wire n_6645;
wire n_6646;
wire n_6647;
wire n_6648;
wire n_6649;
wire n_665;
wire n_6650;
wire n_6651;
wire n_6652;
wire n_6653;
wire n_6654;
wire n_6655;
wire n_6656;
wire n_6657;
wire n_6658;
wire n_6659;
wire n_666;
wire n_6660;
wire n_6661;
wire n_6662;
wire n_6663;
wire n_6664;
wire n_6665;
wire n_6666;
wire n_6667;
wire n_6668;
wire n_6669;
wire n_667;
wire n_6670;
wire n_6671;
wire n_6672;
wire n_6673;
wire n_6674;
wire n_6675;
wire n_6676;
wire n_6677;
wire n_6678;
wire n_6679;
wire n_668;
wire n_6680;
wire n_6681;
wire n_6682;
wire n_6683;
wire n_6684;
wire n_6685;
wire n_6686;
wire n_6687;
wire n_6688;
wire n_6689;
wire n_669;
wire n_6690;
wire n_6691;
wire n_6692;
wire n_6693;
wire n_6694;
wire n_6695;
wire n_6696;
wire n_6697;
wire n_6698;
wire n_6699;
wire n_67;
wire n_670;
wire n_6700;
wire n_6701;
wire n_6702;
wire n_6703;
wire n_6704;
wire n_6705;
wire n_6706;
wire n_6707;
wire n_6708;
wire n_6709;
wire n_671;
wire n_6710;
wire n_6711;
wire n_6712;
wire n_6713;
wire n_6714;
wire n_6715;
wire n_6716;
wire n_6717;
wire n_6718;
wire n_6719;
wire n_672;
wire n_6720;
wire n_6721;
wire n_6722;
wire n_6723;
wire n_6724;
wire n_6725;
wire n_6726;
wire n_6727;
wire n_6728;
wire n_6729;
wire n_673;
wire n_6730;
wire n_6731;
wire n_6732;
wire n_6733;
wire n_6734;
wire n_6735;
wire n_6736;
wire n_6737;
wire n_6738;
wire n_6739;
wire n_674;
wire n_6740;
wire n_6741;
wire n_6742;
wire n_6743;
wire n_6744;
wire n_6745;
wire n_6746;
wire n_6747;
wire n_6748;
wire n_6749;
wire n_675;
wire n_6750;
wire n_6751;
wire n_6752;
wire n_6753;
wire n_6754;
wire n_6755;
wire n_6756;
wire n_6757;
wire n_6758;
wire n_6759;
wire n_676;
wire n_6760;
wire n_6761;
wire n_6762;
wire n_6763;
wire n_6764;
wire n_6765;
wire n_6766;
wire n_6767;
wire n_6768;
wire n_6769;
wire n_677;
wire n_6770;
wire n_6771;
wire n_6772;
wire n_6773;
wire n_6774;
wire n_6775;
wire n_6776;
wire n_6777;
wire n_6778;
wire n_6779;
wire n_678;
wire n_6780;
wire n_6781;
wire n_6782;
wire n_6783;
wire n_6784;
wire n_6785;
wire n_6786;
wire n_6787;
wire n_6788;
wire n_6789;
wire n_679;
wire n_6790;
wire n_6791;
wire n_6792;
wire n_6793;
wire n_6794;
wire n_6795;
wire n_6796;
wire n_6797;
wire n_6798;
wire n_6799;
wire n_68;
wire n_680;
wire n_6800;
wire n_6801;
wire n_6802;
wire n_6803;
wire n_6804;
wire n_6805;
wire n_6806;
wire n_6807;
wire n_6808;
wire n_6809;
wire n_681;
wire n_6810;
wire n_6811;
wire n_6812;
wire n_6813;
wire n_6814;
wire n_6815;
wire n_6816;
wire n_6817;
wire n_6818;
wire n_6819;
wire n_682;
wire n_6820;
wire n_6821;
wire n_6822;
wire n_6823;
wire n_6824;
wire n_6825;
wire n_6826;
wire n_6827;
wire n_6828;
wire n_6829;
wire n_683;
wire n_6830;
wire n_6831;
wire n_6832;
wire n_6833;
wire n_6834;
wire n_6835;
wire n_6836;
wire n_6837;
wire n_6838;
wire n_6839;
wire n_684;
wire n_6840;
wire n_6841;
wire n_6842;
wire n_6843;
wire n_6844;
wire n_6845;
wire n_6846;
wire n_6847;
wire n_6848;
wire n_6849;
wire n_685;
wire n_6850;
wire n_6851;
wire n_6852;
wire n_6853;
wire n_6854;
wire n_6855;
wire n_6856;
wire n_6857;
wire n_6858;
wire n_6859;
wire n_686;
wire n_6860;
wire n_6861;
wire n_6862;
wire n_6863;
wire n_6864;
wire n_6865;
wire n_6866;
wire n_6867;
wire n_6868;
wire n_6869;
wire n_687;
wire n_6870;
wire n_6871;
wire n_6872;
wire n_6873;
wire n_6874;
wire n_6875;
wire n_6876;
wire n_6877;
wire n_6878;
wire n_6879;
wire n_688;
wire n_6880;
wire n_6881;
wire n_6882;
wire n_6883;
wire n_6884;
wire n_6885;
wire n_6886;
wire n_6887;
wire n_6888;
wire n_6889;
wire n_689;
wire n_6890;
wire n_6891;
wire n_6892;
wire n_6893;
wire n_6894;
wire n_6895;
wire n_6896;
wire n_6897;
wire n_6898;
wire n_6899;
wire n_69;
wire n_690;
wire n_6900;
wire n_6901;
wire n_6902;
wire n_6903;
wire n_6904;
wire n_6905;
wire n_6906;
wire n_6907;
wire n_6908;
wire n_6909;
wire n_691;
wire n_6910;
wire n_6911;
wire n_6912;
wire n_6913;
wire n_6914;
wire n_6915;
wire n_6916;
wire n_6917;
wire n_6918;
wire n_6919;
wire n_692;
wire n_6920;
wire n_6921;
wire n_6922;
wire n_6923;
wire n_6924;
wire n_6925;
wire n_6926;
wire n_6927;
wire n_6928;
wire n_6929;
wire n_693;
wire n_6930;
wire n_6931;
wire n_6932;
wire n_6933;
wire n_6934;
wire n_6935;
wire n_6936;
wire n_6937;
wire n_6938;
wire n_6939;
wire n_694;
wire n_6940;
wire n_6941;
wire n_6942;
wire n_6943;
wire n_6944;
wire n_6945;
wire n_6946;
wire n_6947;
wire n_6948;
wire n_6949;
wire n_695;
wire n_6950;
wire n_6951;
wire n_6952;
wire n_6953;
wire n_6954;
wire n_6955;
wire n_6956;
wire n_6957;
wire n_6958;
wire n_6959;
wire n_696;
wire n_6960;
wire n_6961;
wire n_6962;
wire n_6963;
wire n_6964;
wire n_6965;
wire n_6966;
wire n_6967;
wire n_6968;
wire n_6969;
wire n_697;
wire n_6970;
wire n_6971;
wire n_6972;
wire n_6973;
wire n_6974;
wire n_6975;
wire n_6976;
wire n_6977;
wire n_6978;
wire n_6979;
wire n_698;
wire n_6980;
wire n_6981;
wire n_6982;
wire n_6983;
wire n_6984;
wire n_6985;
wire n_6986;
wire n_6987;
wire n_6988;
wire n_6989;
wire n_699;
wire n_6990;
wire n_6991;
wire n_6992;
wire n_6993;
wire n_6994;
wire n_6995;
wire n_6996;
wire n_6997;
wire n_6998;
wire n_6999;
wire n_7;
wire n_70;
wire n_700;
wire n_7000;
wire n_7001;
wire n_7002;
wire n_7003;
wire n_7004;
wire n_7005;
wire n_7006;
wire n_7007;
wire n_7008;
wire n_7009;
wire n_701;
wire n_7010;
wire n_7011;
wire n_7012;
wire n_7013;
wire n_7014;
wire n_7015;
wire n_7016;
wire n_7017;
wire n_7018;
wire n_7019;
wire n_702;
wire n_7020;
wire n_7021;
wire n_7022;
wire n_7023;
wire n_7024;
wire n_7025;
wire n_7026;
wire n_7027;
wire n_7028;
wire n_7029;
wire n_703;
wire n_7030;
wire n_7031;
wire n_7032;
wire n_7033;
wire n_7034;
wire n_7035;
wire n_7036;
wire n_7037;
wire n_7038;
wire n_7039;
wire n_704;
wire n_7040;
wire n_7041;
wire n_7042;
wire n_7043;
wire n_7044;
wire n_7045;
wire n_7046;
wire n_7047;
wire n_7048;
wire n_7049;
wire n_705;
wire n_7050;
wire n_7051;
wire n_7052;
wire n_7053;
wire n_7054;
wire n_7055;
wire n_7056;
wire n_7057;
wire n_7058;
wire n_7059;
wire n_706;
wire n_7060;
wire n_7061;
wire n_7062;
wire n_7063;
wire n_7064;
wire n_7065;
wire n_7066;
wire n_7067;
wire n_7068;
wire n_7069;
wire n_707;
wire n_7070;
wire n_7071;
wire n_7072;
wire n_7073;
wire n_7074;
wire n_7075;
wire n_7076;
wire n_7077;
wire n_7078;
wire n_7079;
wire n_708;
wire n_7080;
wire n_7081;
wire n_7082;
wire n_7083;
wire n_7084;
wire n_7085;
wire n_7086;
wire n_7087;
wire n_7088;
wire n_7089;
wire n_709;
wire n_7090;
wire n_7091;
wire n_7092;
wire n_7093;
wire n_7094;
wire n_7095;
wire n_7096;
wire n_7097;
wire n_7098;
wire n_7099;
wire n_71;
wire n_710;
wire n_7100;
wire n_7101;
wire n_7102;
wire n_7103;
wire n_7104;
wire n_7105;
wire n_7106;
wire n_7107;
wire n_7108;
wire n_7109;
wire n_711;
wire n_7110;
wire n_7111;
wire n_7112;
wire n_7113;
wire n_7114;
wire n_7115;
wire n_7116;
wire n_7117;
wire n_7118;
wire n_7119;
wire n_712;
wire n_7120;
wire n_7121;
wire n_7122;
wire n_7123;
wire n_7124;
wire n_7125;
wire n_7126;
wire n_7127;
wire n_7128;
wire n_7129;
wire n_713;
wire n_7130;
wire n_7131;
wire n_7132;
wire n_7133;
wire n_7134;
wire n_7135;
wire n_7136;
wire n_7137;
wire n_7138;
wire n_7139;
wire n_714;
wire n_7140;
wire n_7141;
wire n_7142;
wire n_7143;
wire n_7144;
wire n_7145;
wire n_7146;
wire n_7147;
wire n_7148;
wire n_7149;
wire n_715;
wire n_7150;
wire n_7151;
wire n_7152;
wire n_7153;
wire n_7154;
wire n_7155;
wire n_7156;
wire n_7157;
wire n_7158;
wire n_7159;
wire n_716;
wire n_7160;
wire n_7161;
wire n_7162;
wire n_7163;
wire n_7164;
wire n_7165;
wire n_7166;
wire n_7167;
wire n_7168;
wire n_7169;
wire n_717;
wire n_7170;
wire n_7171;
wire n_7172;
wire n_7173;
wire n_7174;
wire n_7175;
wire n_7176;
wire n_7177;
wire n_7178;
wire n_7179;
wire n_718;
wire n_7180;
wire n_7181;
wire n_7182;
wire n_7183;
wire n_7184;
wire n_7185;
wire n_7186;
wire n_7187;
wire n_7188;
wire n_7189;
wire n_719;
wire n_7190;
wire n_7191;
wire n_7192;
wire n_7193;
wire n_7194;
wire n_7195;
wire n_7196;
wire n_7197;
wire n_7198;
wire n_7199;
wire n_72;
wire n_720;
wire n_7200;
wire n_7201;
wire n_7202;
wire n_7203;
wire n_7204;
wire n_7205;
wire n_7206;
wire n_7207;
wire n_7208;
wire n_7209;
wire n_721;
wire n_7210;
wire n_7211;
wire n_7212;
wire n_7213;
wire n_7214;
wire n_7215;
wire n_7216;
wire n_7217;
wire n_7218;
wire n_7219;
wire n_722;
wire n_7220;
wire n_7221;
wire n_7222;
wire n_7223;
wire n_7224;
wire n_7225;
wire n_7226;
wire n_7227;
wire n_7228;
wire n_7229;
wire n_723;
wire n_7230;
wire n_7231;
wire n_7232;
wire n_7233;
wire n_7234;
wire n_7235;
wire n_7236;
wire n_7237;
wire n_7238;
wire n_7239;
wire n_724;
wire n_7240;
wire n_7241;
wire n_7242;
wire n_7243;
wire n_7244;
wire n_7245;
wire n_7246;
wire n_7247;
wire n_7248;
wire n_7249;
wire n_725;
wire n_7250;
wire n_7251;
wire n_7252;
wire n_7253;
wire n_7254;
wire n_7255;
wire n_7256;
wire n_7257;
wire n_7258;
wire n_7259;
wire n_726;
wire n_7260;
wire n_7261;
wire n_7262;
wire n_7263;
wire n_7264;
wire n_7265;
wire n_7266;
wire n_7267;
wire n_7268;
wire n_7269;
wire n_727;
wire n_7270;
wire n_7271;
wire n_7272;
wire n_7273;
wire n_7274;
wire n_7275;
wire n_7276;
wire n_7277;
wire n_7278;
wire n_7279;
wire n_728;
wire n_7280;
wire n_7281;
wire n_7282;
wire n_7283;
wire n_7284;
wire n_7285;
wire n_7286;
wire n_7287;
wire n_7288;
wire n_7289;
wire n_729;
wire n_7290;
wire n_7291;
wire n_7292;
wire n_7293;
wire n_7294;
wire n_7295;
wire n_7296;
wire n_7297;
wire n_7298;
wire n_7299;
wire n_73;
wire n_730;
wire n_7300;
wire n_7301;
wire n_7302;
wire n_7303;
wire n_7304;
wire n_7305;
wire n_7306;
wire n_7307;
wire n_7308;
wire n_7309;
wire n_731;
wire n_7310;
wire n_7311;
wire n_7312;
wire n_7313;
wire n_7314;
wire n_7315;
wire n_7316;
wire n_7317;
wire n_7318;
wire n_7319;
wire n_732;
wire n_7320;
wire n_7321;
wire n_7322;
wire n_7323;
wire n_7324;
wire n_7325;
wire n_7326;
wire n_7327;
wire n_7328;
wire n_7329;
wire n_733;
wire n_7330;
wire n_7331;
wire n_7332;
wire n_7333;
wire n_7334;
wire n_7335;
wire n_7336;
wire n_7337;
wire n_7338;
wire n_7339;
wire n_734;
wire n_7340;
wire n_7341;
wire n_7342;
wire n_7343;
wire n_7344;
wire n_7345;
wire n_7346;
wire n_7347;
wire n_7348;
wire n_7349;
wire n_735;
wire n_7350;
wire n_7351;
wire n_7352;
wire n_7353;
wire n_7354;
wire n_7355;
wire n_7356;
wire n_7357;
wire n_7358;
wire n_7359;
wire n_736;
wire n_7360;
wire n_7361;
wire n_7362;
wire n_7363;
wire n_7364;
wire n_7365;
wire n_7366;
wire n_7367;
wire n_7368;
wire n_7369;
wire n_737;
wire n_7370;
wire n_7371;
wire n_7372;
wire n_7373;
wire n_7374;
wire n_7375;
wire n_7376;
wire n_7377;
wire n_7378;
wire n_7379;
wire n_738;
wire n_7380;
wire n_7381;
wire n_7382;
wire n_7383;
wire n_7384;
wire n_7385;
wire n_7386;
wire n_7387;
wire n_7388;
wire n_7389;
wire n_739;
wire n_7390;
wire n_7391;
wire n_7392;
wire n_7393;
wire n_7394;
wire n_7395;
wire n_7396;
wire n_7397;
wire n_7398;
wire n_7399;
wire n_74;
wire n_740;
wire n_7400;
wire n_7401;
wire n_7402;
wire n_7403;
wire n_7404;
wire n_7405;
wire n_7406;
wire n_7407;
wire n_7408;
wire n_7409;
wire n_741;
wire n_7410;
wire n_7411;
wire n_7412;
wire n_7413;
wire n_7414;
wire n_7415;
wire n_7416;
wire n_7417;
wire n_7418;
wire n_7419;
wire n_742;
wire n_7420;
wire n_7421;
wire n_7422;
wire n_7423;
wire n_7424;
wire n_7425;
wire n_7426;
wire n_7427;
wire n_7428;
wire n_7429;
wire n_743;
wire n_7430;
wire n_7431;
wire n_7432;
wire n_7433;
wire n_7434;
wire n_7435;
wire n_7436;
wire n_7437;
wire n_7438;
wire n_7439;
wire n_744;
wire n_7440;
wire n_7441;
wire n_7442;
wire n_7443;
wire n_7444;
wire n_7445;
wire n_7446;
wire n_7447;
wire n_7448;
wire n_7449;
wire n_745;
wire n_7450;
wire n_7451;
wire n_7452;
wire n_7453;
wire n_7454;
wire n_7455;
wire n_7456;
wire n_7457;
wire n_7458;
wire n_7459;
wire n_746;
wire n_7460;
wire n_7461;
wire n_7462;
wire n_7463;
wire n_7464;
wire n_7465;
wire n_7466;
wire n_7467;
wire n_7468;
wire n_7469;
wire n_747;
wire n_7470;
wire n_7471;
wire n_7472;
wire n_7473;
wire n_7474;
wire n_7475;
wire n_7476;
wire n_7477;
wire n_7478;
wire n_7479;
wire n_748;
wire n_7480;
wire n_7481;
wire n_7482;
wire n_7483;
wire n_7484;
wire n_7485;
wire n_7486;
wire n_7487;
wire n_7488;
wire n_7489;
wire n_749;
wire n_7490;
wire n_7491;
wire n_7492;
wire n_7493;
wire n_7494;
wire n_7495;
wire n_7496;
wire n_7497;
wire n_7498;
wire n_7499;
wire n_75;
wire n_750;
wire n_7500;
wire n_7501;
wire n_7502;
wire n_7503;
wire n_7504;
wire n_7505;
wire n_7506;
wire n_7507;
wire n_7508;
wire n_7509;
wire n_751;
wire n_7510;
wire n_7511;
wire n_7512;
wire n_7513;
wire n_7514;
wire n_7515;
wire n_7516;
wire n_7517;
wire n_7518;
wire n_7519;
wire n_752;
wire n_7520;
wire n_7521;
wire n_7522;
wire n_7523;
wire n_7524;
wire n_7525;
wire n_7526;
wire n_7527;
wire n_7528;
wire n_7529;
wire n_753;
wire n_7530;
wire n_7531;
wire n_7532;
wire n_7533;
wire n_7534;
wire n_7535;
wire n_7536;
wire n_7537;
wire n_7538;
wire n_7539;
wire n_754;
wire n_7540;
wire n_7541;
wire n_7542;
wire n_7543;
wire n_7544;
wire n_7545;
wire n_7546;
wire n_7547;
wire n_7548;
wire n_7549;
wire n_755;
wire n_7550;
wire n_7551;
wire n_7552;
wire n_7553;
wire n_7554;
wire n_7555;
wire n_7556;
wire n_7557;
wire n_7558;
wire n_7559;
wire n_756;
wire n_7560;
wire n_7561;
wire n_7562;
wire n_7563;
wire n_7564;
wire n_7565;
wire n_7566;
wire n_7567;
wire n_7568;
wire n_7569;
wire n_757;
wire n_7570;
wire n_7571;
wire n_7572;
wire n_7573;
wire n_7574;
wire n_7575;
wire n_7576;
wire n_7577;
wire n_7578;
wire n_7579;
wire n_758;
wire n_7580;
wire n_7581;
wire n_7582;
wire n_7583;
wire n_7584;
wire n_7585;
wire n_7586;
wire n_7587;
wire n_7588;
wire n_7589;
wire n_759;
wire n_7590;
wire n_7591;
wire n_7592;
wire n_7593;
wire n_7594;
wire n_7595;
wire n_7596;
wire n_7597;
wire n_7598;
wire n_7599;
wire n_76;
wire n_760;
wire n_7600;
wire n_7601;
wire n_7602;
wire n_7603;
wire n_7604;
wire n_7605;
wire n_7606;
wire n_7607;
wire n_7608;
wire n_7609;
wire n_761;
wire n_7610;
wire n_7611;
wire n_7612;
wire n_7613;
wire n_7614;
wire n_7615;
wire n_7616;
wire n_7617;
wire n_7618;
wire n_7619;
wire n_762;
wire n_7620;
wire n_7621;
wire n_7622;
wire n_7623;
wire n_7624;
wire n_7625;
wire n_7626;
wire n_7627;
wire n_7628;
wire n_7629;
wire n_763;
wire n_7630;
wire n_7631;
wire n_7632;
wire n_7633;
wire n_7634;
wire n_7635;
wire n_7636;
wire n_7637;
wire n_7638;
wire n_7639;
wire n_764;
wire n_7640;
wire n_7641;
wire n_7642;
wire n_7643;
wire n_7644;
wire n_7645;
wire n_7646;
wire n_7647;
wire n_7648;
wire n_7649;
wire n_765;
wire n_7650;
wire n_7651;
wire n_7652;
wire n_7653;
wire n_7654;
wire n_7655;
wire n_7656;
wire n_7657;
wire n_7658;
wire n_7659;
wire n_766;
wire n_7660;
wire n_7661;
wire n_7662;
wire n_7663;
wire n_7664;
wire n_7665;
wire n_7666;
wire n_7667;
wire n_7668;
wire n_7669;
wire n_767;
wire n_7670;
wire n_7671;
wire n_7672;
wire n_7673;
wire n_7674;
wire n_7675;
wire n_7676;
wire n_7677;
wire n_7678;
wire n_7679;
wire n_768;
wire n_7680;
wire n_7681;
wire n_7682;
wire n_7683;
wire n_7684;
wire n_7685;
wire n_7686;
wire n_7687;
wire n_7688;
wire n_7689;
wire n_769;
wire n_7690;
wire n_7691;
wire n_7692;
wire n_7693;
wire n_7694;
wire n_7695;
wire n_7696;
wire n_7697;
wire n_7698;
wire n_7699;
wire n_77;
wire n_770;
wire n_7700;
wire n_7701;
wire n_7702;
wire n_7703;
wire n_7704;
wire n_7705;
wire n_7706;
wire n_7707;
wire n_7708;
wire n_7709;
wire n_771;
wire n_7710;
wire n_7711;
wire n_7712;
wire n_7713;
wire n_7714;
wire n_7715;
wire n_7716;
wire n_7717;
wire n_7718;
wire n_7719;
wire n_772;
wire n_7720;
wire n_7721;
wire n_7722;
wire n_7723;
wire n_7724;
wire n_7725;
wire n_7726;
wire n_7727;
wire n_7728;
wire n_7729;
wire n_773;
wire n_7730;
wire n_7731;
wire n_7732;
wire n_7733;
wire n_7734;
wire n_7735;
wire n_7736;
wire n_7737;
wire n_7738;
wire n_7739;
wire n_774;
wire n_7740;
wire n_7741;
wire n_7742;
wire n_7743;
wire n_7744;
wire n_7745;
wire n_7746;
wire n_7747;
wire n_7748;
wire n_7749;
wire n_775;
wire n_7750;
wire n_7751;
wire n_7752;
wire n_7753;
wire n_7754;
wire n_7755;
wire n_7756;
wire n_7757;
wire n_7758;
wire n_7759;
wire n_776;
wire n_7760;
wire n_7761;
wire n_7762;
wire n_7763;
wire n_7764;
wire n_7765;
wire n_7766;
wire n_7767;
wire n_7768;
wire n_7769;
wire n_777;
wire n_7770;
wire n_7771;
wire n_7772;
wire n_7773;
wire n_7774;
wire n_7775;
wire n_7776;
wire n_7777;
wire n_7778;
wire n_7779;
wire n_778;
wire n_7780;
wire n_7781;
wire n_7782;
wire n_7783;
wire n_7784;
wire n_7785;
wire n_7786;
wire n_7787;
wire n_7788;
wire n_7789;
wire n_779;
wire n_7790;
wire n_7791;
wire n_7792;
wire n_7793;
wire n_7794;
wire n_7795;
wire n_7796;
wire n_7797;
wire n_7798;
wire n_7799;
wire n_78;
wire n_780;
wire n_7800;
wire n_7801;
wire n_7802;
wire n_7803;
wire n_7804;
wire n_7805;
wire n_7806;
wire n_7807;
wire n_7808;
wire n_7809;
wire n_781;
wire n_7810;
wire n_7811;
wire n_7812;
wire n_7813;
wire n_7814;
wire n_7815;
wire n_7816;
wire n_7817;
wire n_7818;
wire n_7819;
wire n_782;
wire n_7820;
wire n_7821;
wire n_7822;
wire n_7823;
wire n_7824;
wire n_7825;
wire n_7826;
wire n_7827;
wire n_7828;
wire n_7829;
wire n_783;
wire n_7830;
wire n_7831;
wire n_7832;
wire n_7833;
wire n_7834;
wire n_7835;
wire n_7836;
wire n_7837;
wire n_7838;
wire n_7839;
wire n_784;
wire n_7840;
wire n_7841;
wire n_7842;
wire n_7843;
wire n_7844;
wire n_7845;
wire n_7846;
wire n_7847;
wire n_7848;
wire n_7849;
wire n_785;
wire n_7850;
wire n_7851;
wire n_7852;
wire n_7853;
wire n_7854;
wire n_7855;
wire n_7856;
wire n_7857;
wire n_7858;
wire n_7859;
wire n_786;
wire n_7860;
wire n_7861;
wire n_7862;
wire n_7863;
wire n_7864;
wire n_7865;
wire n_7866;
wire n_7867;
wire n_7868;
wire n_7869;
wire n_787;
wire n_7870;
wire n_7871;
wire n_7872;
wire n_7873;
wire n_7874;
wire n_7875;
wire n_7876;
wire n_7877;
wire n_7878;
wire n_7879;
wire n_788;
wire n_7880;
wire n_7881;
wire n_7882;
wire n_7883;
wire n_7884;
wire n_7885;
wire n_7886;
wire n_7887;
wire n_7888;
wire n_7889;
wire n_789;
wire n_7890;
wire n_7891;
wire n_7892;
wire n_7893;
wire n_7894;
wire n_7895;
wire n_7896;
wire n_7897;
wire n_7898;
wire n_7899;
wire n_79;
wire n_790;
wire n_7900;
wire n_7901;
wire n_7902;
wire n_7903;
wire n_7904;
wire n_7905;
wire n_7906;
wire n_7907;
wire n_7908;
wire n_7909;
wire n_791;
wire n_7910;
wire n_7911;
wire n_7912;
wire n_7913;
wire n_7914;
wire n_7915;
wire n_7916;
wire n_7917;
wire n_7918;
wire n_7919;
wire n_792;
wire n_7920;
wire n_7921;
wire n_7922;
wire n_7923;
wire n_7924;
wire n_7925;
wire n_7926;
wire n_7927;
wire n_7928;
wire n_7929;
wire n_793;
wire n_7930;
wire n_7931;
wire n_7932;
wire n_7933;
wire n_7934;
wire n_7935;
wire n_7936;
wire n_7937;
wire n_7938;
wire n_7939;
wire n_794;
wire n_7940;
wire n_7941;
wire n_7942;
wire n_7943;
wire n_7944;
wire n_7945;
wire n_7946;
wire n_7947;
wire n_7948;
wire n_7949;
wire n_795;
wire n_7950;
wire n_7951;
wire n_7952;
wire n_7953;
wire n_7954;
wire n_7955;
wire n_7956;
wire n_7957;
wire n_7958;
wire n_7959;
wire n_796;
wire n_7960;
wire n_7961;
wire n_7962;
wire n_7963;
wire n_7964;
wire n_7965;
wire n_7966;
wire n_7967;
wire n_7968;
wire n_7969;
wire n_797;
wire n_7970;
wire n_7971;
wire n_7972;
wire n_7973;
wire n_7974;
wire n_7975;
wire n_7976;
wire n_7977;
wire n_7978;
wire n_7979;
wire n_798;
wire n_7980;
wire n_7981;
wire n_7982;
wire n_7983;
wire n_7984;
wire n_7985;
wire n_7986;
wire n_7987;
wire n_7988;
wire n_7989;
wire n_799;
wire n_7990;
wire n_7991;
wire n_7992;
wire n_7993;
wire n_7994;
wire n_7995;
wire n_7996;
wire n_7997;
wire n_7998;
wire n_7999;
wire n_8;
wire n_80;
wire n_800;
wire n_8000;
wire n_8001;
wire n_8002;
wire n_8003;
wire n_8004;
wire n_8005;
wire n_8006;
wire n_8007;
wire n_8008;
wire n_8009;
wire n_801;
wire n_8010;
wire n_8011;
wire n_8012;
wire n_8013;
wire n_8014;
wire n_8015;
wire n_8017;
wire n_8018;
wire n_8019;
wire n_802;
wire n_8020;
wire n_8021;
wire n_8022;
wire n_8023;
wire n_8024;
wire n_8025;
wire n_8026;
wire n_8027;
wire n_8028;
wire n_8029;
wire n_803;
wire n_8030;
wire n_8031;
wire n_8032;
wire n_8033;
wire n_8034;
wire n_8035;
wire n_8036;
wire n_8037;
wire n_8038;
wire n_8039;
wire n_804;
wire n_8040;
wire n_8041;
wire n_8042;
wire n_8043;
wire n_8044;
wire n_8045;
wire n_8046;
wire n_8047;
wire n_8048;
wire n_8049;
wire n_805;
wire n_8050;
wire n_8051;
wire n_8052;
wire n_8053;
wire n_8054;
wire n_8055;
wire n_8056;
wire n_8057;
wire n_8058;
wire n_8059;
wire n_806;
wire n_8060;
wire n_8061;
wire n_8062;
wire n_8063;
wire n_8064;
wire n_8065;
wire n_8066;
wire n_8067;
wire n_8068;
wire n_8069;
wire n_807;
wire n_8070;
wire n_8071;
wire n_8072;
wire n_8073;
wire n_8074;
wire n_8075;
wire n_8076;
wire n_8077;
wire n_8078;
wire n_8079;
wire n_808;
wire n_8080;
wire n_8081;
wire n_8082;
wire n_8083;
wire n_8084;
wire n_8085;
wire n_8086;
wire n_8087;
wire n_8088;
wire n_8089;
wire n_809;
wire n_8090;
wire n_8091;
wire n_8092;
wire n_8093;
wire n_8094;
wire n_8095;
wire n_8096;
wire n_8097;
wire n_8098;
wire n_8099;
wire n_81;
wire n_810;
wire n_8100;
wire n_8101;
wire n_8102;
wire n_8103;
wire n_8104;
wire n_8105;
wire n_8106;
wire n_8107;
wire n_8108;
wire n_8109;
wire n_811;
wire n_8110;
wire n_8111;
wire n_8112;
wire n_8113;
wire n_8114;
wire n_8115;
wire n_8116;
wire n_8117;
wire n_8118;
wire n_8119;
wire n_812;
wire n_8120;
wire n_8121;
wire n_8122;
wire n_8123;
wire n_8124;
wire n_8125;
wire n_8126;
wire n_8127;
wire n_8128;
wire n_8129;
wire n_813;
wire n_8130;
wire n_8131;
wire n_8132;
wire n_8133;
wire n_8134;
wire n_8135;
wire n_8136;
wire n_8137;
wire n_8138;
wire n_8139;
wire n_814;
wire n_8140;
wire n_8141;
wire n_8142;
wire n_8143;
wire n_8144;
wire n_8145;
wire n_8146;
wire n_8147;
wire n_8148;
wire n_8149;
wire n_815;
wire n_8150;
wire n_8151;
wire n_8152;
wire n_8153;
wire n_8154;
wire n_8155;
wire n_8156;
wire n_8157;
wire n_8158;
wire n_8159;
wire n_816;
wire n_8160;
wire n_8161;
wire n_8162;
wire n_8163;
wire n_8164;
wire n_8165;
wire n_8166;
wire n_8167;
wire n_8168;
wire n_8169;
wire n_817;
wire n_8170;
wire n_8171;
wire n_8172;
wire n_8173;
wire n_8174;
wire n_8175;
wire n_8176;
wire n_8177;
wire n_8178;
wire n_8179;
wire n_818;
wire n_8180;
wire n_8181;
wire n_8182;
wire n_8183;
wire n_8184;
wire n_8185;
wire n_8186;
wire n_8187;
wire n_8188;
wire n_8189;
wire n_819;
wire n_8190;
wire n_8191;
wire n_8192;
wire n_8193;
wire n_8194;
wire n_8195;
wire n_8196;
wire n_8197;
wire n_8198;
wire n_8199;
wire n_82;
wire n_820;
wire n_8200;
wire n_8201;
wire n_8202;
wire n_8203;
wire n_8204;
wire n_8205;
wire n_8206;
wire n_8207;
wire n_8208;
wire n_8209;
wire n_821;
wire n_8210;
wire n_8211;
wire n_8212;
wire n_8213;
wire n_8214;
wire n_8215;
wire n_8216;
wire n_8217;
wire n_8218;
wire n_8219;
wire n_822;
wire n_8220;
wire n_8221;
wire n_8222;
wire n_8223;
wire n_8224;
wire n_8225;
wire n_8226;
wire n_8227;
wire n_8228;
wire n_8229;
wire n_823;
wire n_8230;
wire n_8231;
wire n_8232;
wire n_8233;
wire n_8234;
wire n_8235;
wire n_8236;
wire n_8237;
wire n_8238;
wire n_8239;
wire n_824;
wire n_8240;
wire n_8241;
wire n_8242;
wire n_8243;
wire n_8244;
wire n_8245;
wire n_8246;
wire n_8247;
wire n_8248;
wire n_8249;
wire n_825;
wire n_8250;
wire n_8251;
wire n_8252;
wire n_8253;
wire n_8254;
wire n_8255;
wire n_8256;
wire n_8257;
wire n_8258;
wire n_8259;
wire n_826;
wire n_8260;
wire n_8261;
wire n_8262;
wire n_8263;
wire n_8264;
wire n_8265;
wire n_8266;
wire n_8267;
wire n_8268;
wire n_8269;
wire n_827;
wire n_8270;
wire n_8271;
wire n_8272;
wire n_8273;
wire n_8274;
wire n_8275;
wire n_8276;
wire n_8277;
wire n_8278;
wire n_8279;
wire n_828;
wire n_8280;
wire n_8281;
wire n_8282;
wire n_8283;
wire n_8284;
wire n_8285;
wire n_8286;
wire n_8287;
wire n_8288;
wire n_8289;
wire n_829;
wire n_8290;
wire n_8291;
wire n_8292;
wire n_8293;
wire n_8294;
wire n_8295;
wire n_8296;
wire n_8297;
wire n_8298;
wire n_8299;
wire n_83;
wire n_830;
wire n_8300;
wire n_8301;
wire n_8302;
wire n_8303;
wire n_8304;
wire n_8305;
wire n_8306;
wire n_8307;
wire n_8308;
wire n_8309;
wire n_831;
wire n_8310;
wire n_8311;
wire n_8312;
wire n_8313;
wire n_8314;
wire n_8315;
wire n_8316;
wire n_8317;
wire n_8318;
wire n_8319;
wire n_832;
wire n_8320;
wire n_8321;
wire n_8322;
wire n_8323;
wire n_8324;
wire n_8325;
wire n_8326;
wire n_8327;
wire n_8328;
wire n_8329;
wire n_833;
wire n_8330;
wire n_8331;
wire n_8332;
wire n_8333;
wire n_8334;
wire n_8335;
wire n_8336;
wire n_8337;
wire n_8338;
wire n_8339;
wire n_834;
wire n_8340;
wire n_8341;
wire n_8342;
wire n_8343;
wire n_8344;
wire n_8345;
wire n_8346;
wire n_8347;
wire n_8348;
wire n_8349;
wire n_835;
wire n_8350;
wire n_8351;
wire n_8352;
wire n_8353;
wire n_8354;
wire n_8355;
wire n_8356;
wire n_8357;
wire n_8358;
wire n_8359;
wire n_836;
wire n_8360;
wire n_8361;
wire n_8362;
wire n_8363;
wire n_8364;
wire n_8365;
wire n_8366;
wire n_8367;
wire n_8368;
wire n_8369;
wire n_837;
wire n_8370;
wire n_8371;
wire n_8372;
wire n_8373;
wire n_8374;
wire n_8375;
wire n_8376;
wire n_8377;
wire n_8378;
wire n_8379;
wire n_838;
wire n_8380;
wire n_8381;
wire n_8382;
wire n_8383;
wire n_8384;
wire n_8385;
wire n_8386;
wire n_8387;
wire n_8388;
wire n_8389;
wire n_839;
wire n_8390;
wire n_8391;
wire n_8392;
wire n_8393;
wire n_8394;
wire n_8395;
wire n_8396;
wire n_8397;
wire n_8398;
wire n_8399;
wire n_84;
wire n_840;
wire n_8400;
wire n_8401;
wire n_8402;
wire n_8403;
wire n_8404;
wire n_8405;
wire n_8406;
wire n_8407;
wire n_8408;
wire n_8409;
wire n_841;
wire n_8410;
wire n_8411;
wire n_8412;
wire n_8413;
wire n_8414;
wire n_8415;
wire n_8416;
wire n_8417;
wire n_8418;
wire n_8419;
wire n_842;
wire n_8420;
wire n_8421;
wire n_8422;
wire n_8423;
wire n_8424;
wire n_8425;
wire n_8426;
wire n_8427;
wire n_8428;
wire n_8429;
wire n_843;
wire n_8430;
wire n_8431;
wire n_8432;
wire n_8433;
wire n_8434;
wire n_8435;
wire n_8436;
wire n_8437;
wire n_8438;
wire n_8439;
wire n_844;
wire n_8440;
wire n_8441;
wire n_8442;
wire n_8443;
wire n_8444;
wire n_8445;
wire n_8446;
wire n_8447;
wire n_8448;
wire n_8449;
wire n_845;
wire n_8450;
wire n_8451;
wire n_8452;
wire n_8453;
wire n_8454;
wire n_8455;
wire n_8456;
wire n_8457;
wire n_8458;
wire n_8459;
wire n_846;
wire n_8460;
wire n_8461;
wire n_8462;
wire n_8463;
wire n_8464;
wire n_8465;
wire n_8466;
wire n_8467;
wire n_8468;
wire n_8469;
wire n_847;
wire n_8470;
wire n_8471;
wire n_8472;
wire n_8473;
wire n_8474;
wire n_8475;
wire n_8476;
wire n_8477;
wire n_8478;
wire n_8479;
wire n_848;
wire n_8480;
wire n_8481;
wire n_8482;
wire n_8483;
wire n_8484;
wire n_8485;
wire n_8486;
wire n_8487;
wire n_8488;
wire n_8489;
wire n_849;
wire n_8490;
wire n_8491;
wire n_8492;
wire n_8493;
wire n_8494;
wire n_8495;
wire n_8496;
wire n_8497;
wire n_8498;
wire n_8499;
wire n_85;
wire n_850;
wire n_8500;
wire n_8501;
wire n_8502;
wire n_8503;
wire n_8504;
wire n_8505;
wire n_8506;
wire n_8507;
wire n_8508;
wire n_8509;
wire n_851;
wire n_8510;
wire n_8511;
wire n_8512;
wire n_8513;
wire n_8514;
wire n_8515;
wire n_8516;
wire n_8517;
wire n_8518;
wire n_8519;
wire n_852;
wire n_8520;
wire n_8521;
wire n_8522;
wire n_8523;
wire n_8524;
wire n_8525;
wire n_8526;
wire n_8527;
wire n_8528;
wire n_8529;
wire n_853;
wire n_8530;
wire n_8531;
wire n_8532;
wire n_8533;
wire n_8534;
wire n_8535;
wire n_8536;
wire n_8537;
wire n_8538;
wire n_8539;
wire n_854;
wire n_8540;
wire n_8541;
wire n_8542;
wire n_8543;
wire n_8544;
wire n_8545;
wire n_8546;
wire n_8547;
wire n_8548;
wire n_8549;
wire n_855;
wire n_8550;
wire n_8551;
wire n_8552;
wire n_8553;
wire n_8554;
wire n_8555;
wire n_8556;
wire n_8557;
wire n_8558;
wire n_8559;
wire n_856;
wire n_8560;
wire n_8561;
wire n_8562;
wire n_8563;
wire n_8564;
wire n_8565;
wire n_8566;
wire n_8567;
wire n_8568;
wire n_8569;
wire n_857;
wire n_8570;
wire n_8571;
wire n_8572;
wire n_8573;
wire n_8574;
wire n_8575;
wire n_8576;
wire n_8577;
wire n_8578;
wire n_8579;
wire n_858;
wire n_8580;
wire n_8581;
wire n_8582;
wire n_8583;
wire n_8584;
wire n_8585;
wire n_8586;
wire n_8587;
wire n_8588;
wire n_8589;
wire n_859;
wire n_8590;
wire n_8591;
wire n_8592;
wire n_8593;
wire n_8594;
wire n_8595;
wire n_8596;
wire n_8597;
wire n_8598;
wire n_8599;
wire n_86;
wire n_860;
wire n_8600;
wire n_8601;
wire n_8602;
wire n_8603;
wire n_8604;
wire n_8605;
wire n_8606;
wire n_8607;
wire n_8608;
wire n_8609;
wire n_861;
wire n_8610;
wire n_8611;
wire n_8612;
wire n_8613;
wire n_8614;
wire n_8615;
wire n_8616;
wire n_8617;
wire n_8618;
wire n_8619;
wire n_862;
wire n_8620;
wire n_8621;
wire n_8622;
wire n_8623;
wire n_8624;
wire n_8625;
wire n_8626;
wire n_8627;
wire n_8628;
wire n_8629;
wire n_863;
wire n_8630;
wire n_8631;
wire n_8632;
wire n_8633;
wire n_8634;
wire n_8635;
wire n_8636;
wire n_8637;
wire n_8638;
wire n_8639;
wire n_864;
wire n_8640;
wire n_8641;
wire n_8642;
wire n_8643;
wire n_8644;
wire n_8645;
wire n_8646;
wire n_8647;
wire n_8648;
wire n_8649;
wire n_865;
wire n_8650;
wire n_8651;
wire n_8652;
wire n_8653;
wire n_8654;
wire n_8655;
wire n_8656;
wire n_8657;
wire n_8658;
wire n_8659;
wire n_866;
wire n_8660;
wire n_8661;
wire n_8662;
wire n_8663;
wire n_8664;
wire n_8665;
wire n_8666;
wire n_8667;
wire n_8668;
wire n_8669;
wire n_867;
wire n_8670;
wire n_8671;
wire n_8672;
wire n_8673;
wire n_8674;
wire n_8675;
wire n_8676;
wire n_8677;
wire n_8678;
wire n_8679;
wire n_868;
wire n_8680;
wire n_8681;
wire n_8682;
wire n_8683;
wire n_8684;
wire n_8685;
wire n_8686;
wire n_8687;
wire n_8688;
wire n_8689;
wire n_869;
wire n_8690;
wire n_8691;
wire n_8692;
wire n_8693;
wire n_8694;
wire n_8695;
wire n_8696;
wire n_8697;
wire n_8698;
wire n_8699;
wire n_87;
wire n_870;
wire n_8700;
wire n_8701;
wire n_8702;
wire n_8703;
wire n_8704;
wire n_8705;
wire n_8706;
wire n_8707;
wire n_8708;
wire n_8709;
wire n_871;
wire n_8710;
wire n_8711;
wire n_8712;
wire n_8713;
wire n_8714;
wire n_8715;
wire n_8716;
wire n_8717;
wire n_8718;
wire n_8719;
wire n_872;
wire n_8720;
wire n_8721;
wire n_8722;
wire n_8723;
wire n_8724;
wire n_8725;
wire n_8726;
wire n_8727;
wire n_8728;
wire n_8729;
wire n_873;
wire n_8730;
wire n_8731;
wire n_8732;
wire n_8733;
wire n_8734;
wire n_8735;
wire n_8736;
wire n_8737;
wire n_8738;
wire n_8739;
wire n_874;
wire n_8740;
wire n_8741;
wire n_8742;
wire n_8743;
wire n_8744;
wire n_8745;
wire n_8746;
wire n_8747;
wire n_8748;
wire n_8749;
wire n_875;
wire n_8750;
wire n_8751;
wire n_8752;
wire n_8753;
wire n_8754;
wire n_8755;
wire n_8756;
wire n_8757;
wire n_8758;
wire n_8759;
wire n_876;
wire n_8760;
wire n_8761;
wire n_8762;
wire n_8763;
wire n_8764;
wire n_8765;
wire n_8766;
wire n_8767;
wire n_8768;
wire n_8769;
wire n_877;
wire n_8770;
wire n_8771;
wire n_8772;
wire n_8773;
wire n_8774;
wire n_8775;
wire n_8776;
wire n_8777;
wire n_8778;
wire n_8779;
wire n_878;
wire n_8780;
wire n_8781;
wire n_8782;
wire n_8783;
wire n_8784;
wire n_8785;
wire n_8786;
wire n_8787;
wire n_8788;
wire n_8789;
wire n_879;
wire n_8790;
wire n_8791;
wire n_8792;
wire n_8793;
wire n_8794;
wire n_8795;
wire n_8796;
wire n_8797;
wire n_8798;
wire n_8799;
wire n_88;
wire n_880;
wire n_8800;
wire n_8801;
wire n_8802;
wire n_8803;
wire n_8804;
wire n_8805;
wire n_8806;
wire n_8807;
wire n_8808;
wire n_8809;
wire n_881;
wire n_8810;
wire n_8811;
wire n_8812;
wire n_8813;
wire n_8814;
wire n_8815;
wire n_8816;
wire n_8817;
wire n_8818;
wire n_8819;
wire n_882;
wire n_8820;
wire n_8821;
wire n_8822;
wire n_8823;
wire n_8824;
wire n_8825;
wire n_8826;
wire n_8827;
wire n_8828;
wire n_8829;
wire n_883;
wire n_8830;
wire n_8831;
wire n_8832;
wire n_8833;
wire n_8834;
wire n_8835;
wire n_8836;
wire n_8837;
wire n_8838;
wire n_8839;
wire n_884;
wire n_8840;
wire n_8841;
wire n_8842;
wire n_8843;
wire n_8844;
wire n_8845;
wire n_8846;
wire n_8847;
wire n_8848;
wire n_8849;
wire n_885;
wire n_8850;
wire n_8851;
wire n_8852;
wire n_8853;
wire n_8854;
wire n_8855;
wire n_8856;
wire n_8857;
wire n_8858;
wire n_8859;
wire n_886;
wire n_8860;
wire n_8861;
wire n_8862;
wire n_8863;
wire n_8864;
wire n_8865;
wire n_8866;
wire n_8867;
wire n_8868;
wire n_8869;
wire n_887;
wire n_8870;
wire n_8871;
wire n_8872;
wire n_8873;
wire n_8874;
wire n_8875;
wire n_8876;
wire n_8877;
wire n_8878;
wire n_8879;
wire n_888;
wire n_8880;
wire n_8881;
wire n_8882;
wire n_8883;
wire n_8884;
wire n_8885;
wire n_8886;
wire n_8887;
wire n_8888;
wire n_8889;
wire n_889;
wire n_8890;
wire n_8891;
wire n_8892;
wire n_8893;
wire n_8894;
wire n_8895;
wire n_8896;
wire n_8897;
wire n_8898;
wire n_8899;
wire n_89;
wire n_890;
wire n_8900;
wire n_8901;
wire n_8902;
wire n_8903;
wire n_8904;
wire n_8905;
wire n_8906;
wire n_8907;
wire n_8908;
wire n_8909;
wire n_891;
wire n_8910;
wire n_8911;
wire n_8912;
wire n_8913;
wire n_8914;
wire n_8915;
wire n_8916;
wire n_8917;
wire n_8918;
wire n_8919;
wire n_892;
wire n_8920;
wire n_8921;
wire n_8922;
wire n_8923;
wire n_8924;
wire n_8925;
wire n_8926;
wire n_8927;
wire n_8928;
wire n_8929;
wire n_893;
wire n_8930;
wire n_8931;
wire n_8932;
wire n_8933;
wire n_8934;
wire n_8935;
wire n_8936;
wire n_8937;
wire n_8938;
wire n_8939;
wire n_894;
wire n_8940;
wire n_8941;
wire n_8942;
wire n_8943;
wire n_8944;
wire n_8945;
wire n_8946;
wire n_8947;
wire n_8948;
wire n_8949;
wire n_895;
wire n_8950;
wire n_8951;
wire n_8952;
wire n_8953;
wire n_8954;
wire n_8955;
wire n_8956;
wire n_8957;
wire n_8958;
wire n_8959;
wire n_896;
wire n_8960;
wire n_8961;
wire n_8962;
wire n_8963;
wire n_8964;
wire n_8965;
wire n_8966;
wire n_8967;
wire n_8968;
wire n_8969;
wire n_897;
wire n_8970;
wire n_8971;
wire n_8972;
wire n_8973;
wire n_8974;
wire n_8975;
wire n_8976;
wire n_8977;
wire n_8978;
wire n_8979;
wire n_898;
wire n_8980;
wire n_8981;
wire n_8982;
wire n_8983;
wire n_8984;
wire n_8985;
wire n_8986;
wire n_8987;
wire n_8988;
wire n_8989;
wire n_899;
wire n_8990;
wire n_8991;
wire n_8992;
wire n_8993;
wire n_8994;
wire n_8995;
wire n_8996;
wire n_8997;
wire n_8998;
wire n_8999;
wire n_9;
wire n_90;
wire n_900;
wire n_9000;
wire n_9001;
wire n_9002;
wire n_9003;
wire n_9004;
wire n_9005;
wire n_9006;
wire n_9007;
wire n_9008;
wire n_9009;
wire n_901;
wire n_9010;
wire n_9011;
wire n_9012;
wire n_9013;
wire n_9014;
wire n_9015;
wire n_9016;
wire n_9017;
wire n_9018;
wire n_9019;
wire n_902;
wire n_9020;
wire n_9021;
wire n_9022;
wire n_9023;
wire n_9024;
wire n_9025;
wire n_9026;
wire n_9027;
wire n_9028;
wire n_9029;
wire n_903;
wire n_9030;
wire n_9031;
wire n_9032;
wire n_9033;
wire n_9034;
wire n_9035;
wire n_9036;
wire n_9037;
wire n_9038;
wire n_9039;
wire n_904;
wire n_9040;
wire n_9041;
wire n_9042;
wire n_9043;
wire n_9044;
wire n_9045;
wire n_9046;
wire n_9047;
wire n_9048;
wire n_9049;
wire n_905;
wire n_9050;
wire n_9051;
wire n_9052;
wire n_9053;
wire n_9054;
wire n_9055;
wire n_9056;
wire n_9057;
wire n_9058;
wire n_9059;
wire n_906;
wire n_9060;
wire n_9061;
wire n_9062;
wire n_9063;
wire n_9064;
wire n_9065;
wire n_9066;
wire n_9067;
wire n_9068;
wire n_9069;
wire n_907;
wire n_9070;
wire n_9071;
wire n_9072;
wire n_9073;
wire n_9074;
wire n_9075;
wire n_9076;
wire n_9077;
wire n_9078;
wire n_9079;
wire n_908;
wire n_9080;
wire n_9081;
wire n_9082;
wire n_9083;
wire n_9084;
wire n_9085;
wire n_9086;
wire n_9087;
wire n_9088;
wire n_9089;
wire n_909;
wire n_9090;
wire n_9091;
wire n_9092;
wire n_9093;
wire n_9094;
wire n_9095;
wire n_9096;
wire n_9097;
wire n_9098;
wire n_9099;
wire n_91;
wire n_910;
wire n_9100;
wire n_9101;
wire n_9102;
wire n_9103;
wire n_9104;
wire n_9105;
wire n_9106;
wire n_9107;
wire n_9108;
wire n_9109;
wire n_911;
wire n_9110;
wire n_9111;
wire n_9112;
wire n_9113;
wire n_9114;
wire n_9115;
wire n_9116;
wire n_9117;
wire n_9118;
wire n_9119;
wire n_912;
wire n_9120;
wire n_9121;
wire n_9122;
wire n_9123;
wire n_9124;
wire n_9125;
wire n_9126;
wire n_9127;
wire n_9128;
wire n_9129;
wire n_913;
wire n_9130;
wire n_9131;
wire n_9132;
wire n_9133;
wire n_9134;
wire n_9135;
wire n_9136;
wire n_9137;
wire n_9138;
wire n_9139;
wire n_914;
wire n_9140;
wire n_9141;
wire n_9142;
wire n_9143;
wire n_9144;
wire n_9145;
wire n_9146;
wire n_9147;
wire n_9148;
wire n_9149;
wire n_915;
wire n_9150;
wire n_9151;
wire n_9152;
wire n_9153;
wire n_9154;
wire n_9155;
wire n_9156;
wire n_9157;
wire n_9158;
wire n_9159;
wire n_916;
wire n_9160;
wire n_9161;
wire n_9162;
wire n_9163;
wire n_9164;
wire n_9165;
wire n_9166;
wire n_9167;
wire n_9168;
wire n_9169;
wire n_917;
wire n_9170;
wire n_9171;
wire n_9172;
wire n_9173;
wire n_9174;
wire n_9175;
wire n_9176;
wire n_9177;
wire n_9178;
wire n_9179;
wire n_918;
wire n_9180;
wire n_9181;
wire n_9182;
wire n_9183;
wire n_9184;
wire n_9185;
wire n_9186;
wire n_9187;
wire n_9188;
wire n_9189;
wire n_919;
wire n_9190;
wire n_9191;
wire n_9192;
wire n_9193;
wire n_9194;
wire n_9195;
wire n_9196;
wire n_9197;
wire n_9198;
wire n_9199;
wire n_92;
wire n_920;
wire n_9200;
wire n_9201;
wire n_9202;
wire n_9203;
wire n_9204;
wire n_9205;
wire n_9206;
wire n_9207;
wire n_9208;
wire n_9209;
wire n_921;
wire n_9210;
wire n_9211;
wire n_9212;
wire n_9213;
wire n_9214;
wire n_9215;
wire n_9216;
wire n_9217;
wire n_9218;
wire n_9219;
wire n_922;
wire n_9220;
wire n_9221;
wire n_9222;
wire n_9223;
wire n_9224;
wire n_9225;
wire n_9226;
wire n_9227;
wire n_9228;
wire n_9229;
wire n_923;
wire n_9230;
wire n_9231;
wire n_9232;
wire n_9233;
wire n_9234;
wire n_9235;
wire n_9236;
wire n_9237;
wire n_9238;
wire n_9239;
wire n_924;
wire n_9240;
wire n_9241;
wire n_9242;
wire n_9243;
wire n_9244;
wire n_9245;
wire n_9246;
wire n_9247;
wire n_9248;
wire n_9249;
wire n_925;
wire n_9250;
wire n_9251;
wire n_9252;
wire n_9253;
wire n_9254;
wire n_9255;
wire n_9256;
wire n_9257;
wire n_9258;
wire n_9259;
wire n_926;
wire n_9260;
wire n_9261;
wire n_9262;
wire n_9263;
wire n_9264;
wire n_9265;
wire n_9266;
wire n_9267;
wire n_9268;
wire n_9269;
wire n_927;
wire n_9270;
wire n_9271;
wire n_9272;
wire n_9273;
wire n_9274;
wire n_9275;
wire n_9276;
wire n_9277;
wire n_9278;
wire n_9279;
wire n_928;
wire n_9280;
wire n_9281;
wire n_9282;
wire n_9283;
wire n_9284;
wire n_9285;
wire n_9286;
wire n_9287;
wire n_9288;
wire n_9289;
wire n_929;
wire n_9290;
wire n_9291;
wire n_9292;
wire n_9293;
wire n_9294;
wire n_9295;
wire n_9296;
wire n_9297;
wire n_9298;
wire n_9299;
wire n_93;
wire n_930;
wire n_9300;
wire n_9301;
wire n_9302;
wire n_9303;
wire n_9304;
wire n_9305;
wire n_9306;
wire n_9307;
wire n_9308;
wire n_9309;
wire n_931;
wire n_9310;
wire n_9311;
wire n_9312;
wire n_9313;
wire n_9314;
wire n_9315;
wire n_9316;
wire n_9317;
wire n_9318;
wire n_9319;
wire n_932;
wire n_9320;
wire n_9321;
wire n_9322;
wire n_9323;
wire n_9324;
wire n_9325;
wire n_9326;
wire n_9327;
wire n_9328;
wire n_9329;
wire n_933;
wire n_9330;
wire n_9331;
wire n_9332;
wire n_9333;
wire n_9334;
wire n_9335;
wire n_9336;
wire n_9337;
wire n_9338;
wire n_9339;
wire n_934;
wire n_9340;
wire n_9341;
wire n_9342;
wire n_9343;
wire n_9344;
wire n_9345;
wire n_9346;
wire n_9347;
wire n_9348;
wire n_9349;
wire n_935;
wire n_9350;
wire n_9351;
wire n_9352;
wire n_9353;
wire n_9354;
wire n_9355;
wire n_9356;
wire n_9357;
wire n_9358;
wire n_9359;
wire n_936;
wire n_9360;
wire n_9361;
wire n_9362;
wire n_9363;
wire n_9364;
wire n_9365;
wire n_9366;
wire n_9368;
wire n_9369;
wire n_937;
wire n_9371;
wire n_9372;
wire n_9374;
wire n_9375;
wire n_9377;
wire n_9378;
wire n_938;
wire n_9380;
wire n_9381;
wire n_9383;
wire n_9384;
wire n_9385;
wire n_9386;
wire n_9387;
wire n_9388;
wire n_9389;
wire n_939;
wire n_9390;
wire n_9391;
wire n_9392;
wire n_9393;
wire n_9394;
wire n_9395;
wire n_9396;
wire n_9397;
wire n_9398;
wire n_9399;
wire n_94;
wire n_940;
wire n_9400;
wire n_9401;
wire n_9402;
wire n_9403;
wire n_9404;
wire n_9405;
wire n_9406;
wire n_9407;
wire n_9408;
wire n_9409;
wire n_941;
wire n_9410;
wire n_9411;
wire n_9412;
wire n_9413;
wire n_9414;
wire n_9415;
wire n_9416;
wire n_9417;
wire n_9418;
wire n_9419;
wire n_942;
wire n_9420;
wire n_9421;
wire n_9422;
wire n_9423;
wire n_9424;
wire n_9425;
wire n_9426;
wire n_9427;
wire n_9428;
wire n_9429;
wire n_943;
wire n_9430;
wire n_9431;
wire n_9432;
wire n_9433;
wire n_9434;
wire n_9435;
wire n_9436;
wire n_9437;
wire n_9438;
wire n_9439;
wire n_944;
wire n_9440;
wire n_9441;
wire n_9442;
wire n_9443;
wire n_9444;
wire n_9445;
wire n_9446;
wire n_9447;
wire n_9448;
wire n_9449;
wire n_945;
wire n_9450;
wire n_9451;
wire n_9452;
wire n_9453;
wire n_9454;
wire n_9455;
wire n_9456;
wire n_9457;
wire n_9458;
wire n_9459;
wire n_946;
wire n_9460;
wire n_9461;
wire n_9462;
wire n_9463;
wire n_9464;
wire n_9465;
wire n_9466;
wire n_9467;
wire n_9468;
wire n_9469;
wire n_947;
wire n_9470;
wire n_9471;
wire n_9472;
wire n_9473;
wire n_9474;
wire n_9475;
wire n_9476;
wire n_9477;
wire n_9478;
wire n_9479;
wire n_948;
wire n_9480;
wire n_9481;
wire n_9482;
wire n_9483;
wire n_9484;
wire n_9485;
wire n_9486;
wire n_9487;
wire n_9488;
wire n_9489;
wire n_949;
wire n_9490;
wire n_9491;
wire n_9492;
wire n_9493;
wire n_9494;
wire n_9495;
wire n_9496;
wire n_9497;
wire n_9498;
wire n_9499;
wire n_95;
wire n_950;
wire n_9500;
wire n_9501;
wire n_9502;
wire n_9503;
wire n_9504;
wire n_9505;
wire n_9506;
wire n_9507;
wire n_9508;
wire n_9509;
wire n_951;
wire n_9510;
wire n_9511;
wire n_9512;
wire n_9513;
wire n_9514;
wire n_9515;
wire n_9516;
wire n_9517;
wire n_9518;
wire n_9519;
wire n_952;
wire n_9520;
wire n_9521;
wire n_9522;
wire n_9523;
wire n_9524;
wire n_9525;
wire n_9526;
wire n_9527;
wire n_9528;
wire n_9529;
wire n_953;
wire n_9530;
wire n_9531;
wire n_9532;
wire n_9533;
wire n_9534;
wire n_9535;
wire n_9536;
wire n_9537;
wire n_9538;
wire n_9539;
wire n_954;
wire n_9540;
wire n_9541;
wire n_9542;
wire n_9543;
wire n_9544;
wire n_9545;
wire n_9546;
wire n_9547;
wire n_9548;
wire n_9549;
wire n_955;
wire n_9550;
wire n_9551;
wire n_9552;
wire n_9553;
wire n_9554;
wire n_9555;
wire n_9556;
wire n_9557;
wire n_9558;
wire n_9559;
wire n_956;
wire n_9560;
wire n_9561;
wire n_9562;
wire n_9563;
wire n_9564;
wire n_9565;
wire n_9566;
wire n_9567;
wire n_9568;
wire n_9569;
wire n_957;
wire n_9570;
wire n_9571;
wire n_9572;
wire n_9573;
wire n_9574;
wire n_9575;
wire n_9576;
wire n_9577;
wire n_9578;
wire n_9579;
wire n_958;
wire n_9580;
wire n_9581;
wire n_9582;
wire n_9583;
wire n_9584;
wire n_9585;
wire n_9586;
wire n_9587;
wire n_9588;
wire n_9589;
wire n_959;
wire n_9590;
wire n_9591;
wire n_9592;
wire n_9593;
wire n_9594;
wire n_9595;
wire n_9596;
wire n_9597;
wire n_9598;
wire n_9599;
wire n_96;
wire n_960;
wire n_9600;
wire n_9601;
wire n_9602;
wire n_9603;
wire n_9604;
wire n_9605;
wire n_9606;
wire n_9607;
wire n_9608;
wire n_9609;
wire n_961;
wire n_9610;
wire n_9611;
wire n_9612;
wire n_9613;
wire n_9614;
wire n_9615;
wire n_9616;
wire n_9617;
wire n_9618;
wire n_9619;
wire n_962;
wire n_9620;
wire n_9621;
wire n_9622;
wire n_9623;
wire n_9624;
wire n_9625;
wire n_9626;
wire n_9627;
wire n_9628;
wire n_9629;
wire n_963;
wire n_9630;
wire n_9631;
wire n_9632;
wire n_9633;
wire n_9634;
wire n_9635;
wire n_9636;
wire n_9637;
wire n_9638;
wire n_9639;
wire n_964;
wire n_9640;
wire n_9641;
wire n_9642;
wire n_9643;
wire n_9644;
wire n_9645;
wire n_9646;
wire n_9647;
wire n_9648;
wire n_9649;
wire n_965;
wire n_9650;
wire n_9651;
wire n_9652;
wire n_9653;
wire n_9654;
wire n_9655;
wire n_9656;
wire n_9657;
wire n_9658;
wire n_9659;
wire n_966;
wire n_9660;
wire n_9661;
wire n_9662;
wire n_9663;
wire n_9664;
wire n_9665;
wire n_9666;
wire n_9667;
wire n_9668;
wire n_9669;
wire n_967;
wire n_9670;
wire n_9671;
wire n_9672;
wire n_9673;
wire n_9674;
wire n_9675;
wire n_9676;
wire n_9677;
wire n_9678;
wire n_9679;
wire n_968;
wire n_9680;
wire n_9681;
wire n_9682;
wire n_9683;
wire n_9684;
wire n_9685;
wire n_9686;
wire n_9687;
wire n_9688;
wire n_9689;
wire n_969;
wire n_9690;
wire n_9691;
wire n_9692;
wire n_9693;
wire n_9694;
wire n_9695;
wire n_9696;
wire n_9697;
wire n_9698;
wire n_9699;
wire n_97;
wire n_970;
wire n_9700;
wire n_9701;
wire n_9702;
wire n_9703;
wire n_9704;
wire n_9705;
wire n_9706;
wire n_9707;
wire n_9708;
wire n_9709;
wire n_971;
wire n_9710;
wire n_9711;
wire n_9712;
wire n_9713;
wire n_9714;
wire n_9715;
wire n_9716;
wire n_9717;
wire n_9718;
wire n_9719;
wire n_972;
wire n_9720;
wire n_9721;
wire n_9722;
wire n_9723;
wire n_9724;
wire n_9725;
wire n_9726;
wire n_9727;
wire n_9728;
wire n_9729;
wire n_973;
wire n_9730;
wire n_9731;
wire n_9732;
wire n_9733;
wire n_9734;
wire n_9735;
wire n_9736;
wire n_9737;
wire n_9738;
wire n_9739;
wire n_974;
wire n_9740;
wire n_9741;
wire n_9742;
wire n_9743;
wire n_9744;
wire n_9745;
wire n_9746;
wire n_9747;
wire n_9748;
wire n_9749;
wire n_975;
wire n_9750;
wire n_9751;
wire n_9752;
wire n_9753;
wire n_9754;
wire n_9755;
wire n_9756;
wire n_9757;
wire n_9758;
wire n_9759;
wire n_976;
wire n_9760;
wire n_9761;
wire n_9762;
wire n_9763;
wire n_9764;
wire n_9765;
wire n_9766;
wire n_9767;
wire n_9768;
wire n_9769;
wire n_977;
wire n_9770;
wire n_9771;
wire n_9772;
wire n_9773;
wire n_9774;
wire n_9775;
wire n_9776;
wire n_9777;
wire n_9778;
wire n_9779;
wire n_978;
wire n_9780;
wire n_9781;
wire n_9782;
wire n_9783;
wire n_9784;
wire n_9785;
wire n_9786;
wire n_9787;
wire n_9788;
wire n_9789;
wire n_979;
wire n_9790;
wire n_9791;
wire n_9792;
wire n_9793;
wire n_9794;
wire n_9795;
wire n_9796;
wire n_9797;
wire n_9798;
wire n_9799;
wire n_98;
wire n_980;
wire n_9800;
wire n_9801;
wire n_9802;
wire n_9803;
wire n_9804;
wire n_9805;
wire n_9806;
wire n_9807;
wire n_9808;
wire n_9809;
wire n_981;
wire n_9810;
wire n_9811;
wire n_9812;
wire n_9813;
wire n_9814;
wire n_9815;
wire n_9816;
wire n_9817;
wire n_9818;
wire n_9819;
wire n_982;
wire n_9820;
wire n_9821;
wire n_9822;
wire n_9823;
wire n_9824;
wire n_9825;
wire n_9826;
wire n_9827;
wire n_9828;
wire n_9829;
wire n_983;
wire n_9830;
wire n_9831;
wire n_9832;
wire n_9834;
wire n_9835;
wire n_9836;
wire n_9837;
wire n_9838;
wire n_9839;
wire n_984;
wire n_9840;
wire n_9841;
wire n_9842;
wire n_9843;
wire n_9844;
wire n_9845;
wire n_9846;
wire n_9847;
wire n_9848;
wire n_9849;
wire n_985;
wire n_9850;
wire n_9851;
wire n_9852;
wire n_9853;
wire n_9854;
wire n_9855;
wire n_9856;
wire n_9857;
wire n_9858;
wire n_9859;
wire n_986;
wire n_9860;
wire n_9861;
wire n_9862;
wire n_9863;
wire n_9864;
wire n_9865;
wire n_9866;
wire n_9867;
wire n_9868;
wire n_9869;
wire n_987;
wire n_9870;
wire n_9871;
wire n_9872;
wire n_9873;
wire n_9874;
wire n_9875;
wire n_9876;
wire n_9877;
wire n_9878;
wire n_9879;
wire n_988;
wire n_9880;
wire n_9881;
wire n_9882;
wire n_9883;
wire n_9884;
wire n_9885;
wire n_9886;
wire n_9887;
wire n_9888;
wire n_9889;
wire n_989;
wire n_9890;
wire n_9891;
wire n_9892;
wire n_9893;
wire n_9894;
wire n_9895;
wire n_9896;
wire n_9897;
wire n_9898;
wire n_9899;
wire n_99;
wire n_990;
wire n_9900;
wire n_9901;
wire n_9902;
wire n_9903;
wire n_9904;
wire n_9905;
wire n_9906;
wire n_9907;
wire n_9908;
wire n_9909;
wire n_991;
wire n_9910;
wire n_9911;
wire n_9912;
wire n_9913;
wire n_9914;
wire n_9915;
wire n_9916;
wire n_9917;
wire n_9918;
wire n_9919;
wire n_992;
wire n_9920;
wire n_9921;
wire n_9922;
wire n_9923;
wire n_9924;
wire n_9925;
wire n_9926;
wire n_9927;
wire n_9928;
wire n_9929;
wire n_993;
wire n_9930;
wire n_9931;
wire n_9932;
wire n_9933;
wire n_9934;
wire n_9935;
wire n_9936;
wire n_9937;
wire n_9938;
wire n_9939;
wire n_994;
wire n_9940;
wire n_9941;
wire n_9942;
wire n_9943;
wire n_9944;
wire n_9945;
wire n_9946;
wire n_9947;
wire n_9948;
wire n_9949;
wire n_995;
wire n_9950;
wire n_9951;
wire n_9952;
wire n_9953;
wire n_9954;
wire n_9955;
wire n_9956;
wire n_9957;
wire n_9958;
wire n_9959;
wire n_996;
wire n_9960;
wire n_9961;
wire n_9962;
wire n_9963;
wire n_9964;
wire n_9965;
wire n_9966;
wire n_9967;
wire n_9968;
wire n_9969;
wire n_997;
wire n_9970;
wire n_9971;
wire n_9972;
wire n_9973;
wire n_9974;
wire n_9975;
wire n_9976;
wire n_9977;
wire n_9978;
wire n_9979;
wire n_998;
wire n_9980;
wire n_9981;
wire n_9982;
wire n_9983;
wire n_9984;
wire n_9985;
wire n_9986;
wire n_9987;
wire n_9988;
wire n_9989;
wire n_999;
wire n_9990;
wire n_9991;
wire n_9992;
wire n_9993;
wire n_9994;
wire n_9995;
wire n_9996;
wire n_9997;
wire n_9998;
wire n_9999;
wire rst;
wire x_in_0_0;
wire x_in_0_1;
wire x_in_0_10;
wire x_in_0_11;
wire x_in_0_12;
wire x_in_0_13;
wire x_in_0_14;
wire x_in_0_15;
wire x_in_0_2;
wire x_in_0_3;
wire x_in_0_4;
wire x_in_0_5;
wire x_in_0_6;
wire x_in_0_7;
wire x_in_0_8;
wire x_in_0_9;
wire x_in_10_0;
wire x_in_10_1;
wire x_in_10_10;
wire x_in_10_11;
wire x_in_10_12;
wire x_in_10_13;
wire x_in_10_14;
wire x_in_10_15;
wire x_in_10_2;
wire x_in_10_3;
wire x_in_10_4;
wire x_in_10_5;
wire x_in_10_6;
wire x_in_10_7;
wire x_in_10_8;
wire x_in_10_9;
wire x_in_11_0;
wire x_in_11_1;
wire x_in_11_10;
wire x_in_11_11;
wire x_in_11_12;
wire x_in_11_13;
wire x_in_11_14;
wire x_in_11_15;
wire x_in_11_2;
wire x_in_11_3;
wire x_in_11_4;
wire x_in_11_5;
wire x_in_11_6;
wire x_in_11_7;
wire x_in_11_8;
wire x_in_11_9;
wire x_in_12_0;
wire x_in_12_1;
wire x_in_12_10;
wire x_in_12_11;
wire x_in_12_12;
wire x_in_12_13;
wire x_in_12_14;
wire x_in_12_15;
wire x_in_12_2;
wire x_in_12_3;
wire x_in_12_4;
wire x_in_12_5;
wire x_in_12_6;
wire x_in_12_7;
wire x_in_12_8;
wire x_in_12_9;
wire x_in_13_0;
wire x_in_13_1;
wire x_in_13_10;
wire x_in_13_11;
wire x_in_13_12;
wire x_in_13_13;
wire x_in_13_14;
wire x_in_13_15;
wire x_in_13_2;
wire x_in_13_3;
wire x_in_13_4;
wire x_in_13_5;
wire x_in_13_6;
wire x_in_13_7;
wire x_in_13_8;
wire x_in_13_9;
wire x_in_14_0;
wire x_in_14_1;
wire x_in_14_10;
wire x_in_14_11;
wire x_in_14_12;
wire x_in_14_13;
wire x_in_14_14;
wire x_in_14_15;
wire x_in_14_2;
wire x_in_14_3;
wire x_in_14_4;
wire x_in_14_5;
wire x_in_14_6;
wire x_in_14_7;
wire x_in_14_8;
wire x_in_14_9;
wire x_in_15_0;
wire x_in_15_1;
wire x_in_15_10;
wire x_in_15_11;
wire x_in_15_12;
wire x_in_15_13;
wire x_in_15_14;
wire x_in_15_15;
wire x_in_15_2;
wire x_in_15_3;
wire x_in_15_4;
wire x_in_15_5;
wire x_in_15_6;
wire x_in_15_7;
wire x_in_15_8;
wire x_in_15_9;
wire x_in_16_0;
wire x_in_16_1;
wire x_in_16_10;
wire x_in_16_11;
wire x_in_16_12;
wire x_in_16_13;
wire x_in_16_14;
wire x_in_16_15;
wire x_in_16_2;
wire x_in_16_3;
wire x_in_16_4;
wire x_in_16_5;
wire x_in_16_6;
wire x_in_16_7;
wire x_in_16_8;
wire x_in_16_9;
wire x_in_17_0;
wire x_in_17_1;
wire x_in_17_10;
wire x_in_17_11;
wire x_in_17_12;
wire x_in_17_13;
wire x_in_17_14;
wire x_in_17_15;
wire x_in_17_2;
wire x_in_17_3;
wire x_in_17_4;
wire x_in_17_5;
wire x_in_17_6;
wire x_in_17_7;
wire x_in_17_8;
wire x_in_17_9;
wire x_in_18_0;
wire x_in_18_1;
wire x_in_18_10;
wire x_in_18_11;
wire x_in_18_12;
wire x_in_18_13;
wire x_in_18_14;
wire x_in_18_15;
wire x_in_18_2;
wire x_in_18_3;
wire x_in_18_4;
wire x_in_18_5;
wire x_in_18_6;
wire x_in_18_7;
wire x_in_18_8;
wire x_in_18_9;
wire x_in_19_0;
wire x_in_19_1;
wire x_in_19_10;
wire x_in_19_11;
wire x_in_19_12;
wire x_in_19_13;
wire x_in_19_14;
wire x_in_19_15;
wire x_in_19_2;
wire x_in_19_3;
wire x_in_19_4;
wire x_in_19_5;
wire x_in_19_6;
wire x_in_19_7;
wire x_in_19_8;
wire x_in_19_9;
wire x_in_1_0;
wire x_in_1_1;
wire x_in_1_10;
wire x_in_1_11;
wire x_in_1_12;
wire x_in_1_13;
wire x_in_1_14;
wire x_in_1_15;
wire x_in_1_2;
wire x_in_1_3;
wire x_in_1_4;
wire x_in_1_5;
wire x_in_1_6;
wire x_in_1_7;
wire x_in_1_8;
wire x_in_1_9;
wire x_in_20_0;
wire x_in_20_1;
wire x_in_20_10;
wire x_in_20_11;
wire x_in_20_12;
wire x_in_20_13;
wire x_in_20_14;
wire x_in_20_15;
wire x_in_20_2;
wire x_in_20_3;
wire x_in_20_4;
wire x_in_20_5;
wire x_in_20_6;
wire x_in_20_7;
wire x_in_20_8;
wire x_in_20_9;
wire x_in_21_0;
wire x_in_21_1;
wire x_in_21_10;
wire x_in_21_11;
wire x_in_21_12;
wire x_in_21_13;
wire x_in_21_14;
wire x_in_21_15;
wire x_in_21_2;
wire x_in_21_3;
wire x_in_21_4;
wire x_in_21_5;
wire x_in_21_6;
wire x_in_21_7;
wire x_in_21_8;
wire x_in_21_9;
wire x_in_22_0;
wire x_in_22_1;
wire x_in_22_10;
wire x_in_22_11;
wire x_in_22_12;
wire x_in_22_13;
wire x_in_22_14;
wire x_in_22_15;
wire x_in_22_2;
wire x_in_22_3;
wire x_in_22_4;
wire x_in_22_5;
wire x_in_22_6;
wire x_in_22_7;
wire x_in_22_8;
wire x_in_22_9;
wire x_in_23_0;
wire x_in_23_1;
wire x_in_23_10;
wire x_in_23_11;
wire x_in_23_12;
wire x_in_23_13;
wire x_in_23_14;
wire x_in_23_15;
wire x_in_23_2;
wire x_in_23_3;
wire x_in_23_4;
wire x_in_23_5;
wire x_in_23_6;
wire x_in_23_7;
wire x_in_23_8;
wire x_in_23_9;
wire x_in_24_0;
wire x_in_24_1;
wire x_in_24_10;
wire x_in_24_11;
wire x_in_24_12;
wire x_in_24_13;
wire x_in_24_14;
wire x_in_24_15;
wire x_in_24_2;
wire x_in_24_3;
wire x_in_24_4;
wire x_in_24_5;
wire x_in_24_6;
wire x_in_24_7;
wire x_in_24_8;
wire x_in_24_9;
wire x_in_25_0;
wire x_in_25_1;
wire x_in_25_10;
wire x_in_25_11;
wire x_in_25_12;
wire x_in_25_13;
wire x_in_25_14;
wire x_in_25_15;
wire x_in_25_2;
wire x_in_25_3;
wire x_in_25_4;
wire x_in_25_5;
wire x_in_25_6;
wire x_in_25_7;
wire x_in_25_8;
wire x_in_25_9;
wire x_in_26_0;
wire x_in_26_1;
wire x_in_26_10;
wire x_in_26_11;
wire x_in_26_12;
wire x_in_26_13;
wire x_in_26_14;
wire x_in_26_15;
wire x_in_26_2;
wire x_in_26_3;
wire x_in_26_4;
wire x_in_26_5;
wire x_in_26_6;
wire x_in_26_7;
wire x_in_26_8;
wire x_in_26_9;
wire x_in_27_0;
wire x_in_27_1;
wire x_in_27_10;
wire x_in_27_11;
wire x_in_27_12;
wire x_in_27_13;
wire x_in_27_14;
wire x_in_27_15;
wire x_in_27_2;
wire x_in_27_3;
wire x_in_27_4;
wire x_in_27_5;
wire x_in_27_6;
wire x_in_27_7;
wire x_in_27_8;
wire x_in_27_9;
wire x_in_28_0;
wire x_in_28_1;
wire x_in_28_10;
wire x_in_28_11;
wire x_in_28_12;
wire x_in_28_13;
wire x_in_28_14;
wire x_in_28_15;
wire x_in_28_2;
wire x_in_28_3;
wire x_in_28_4;
wire x_in_28_5;
wire x_in_28_6;
wire x_in_28_7;
wire x_in_28_8;
wire x_in_28_9;
wire x_in_29_0;
wire x_in_29_1;
wire x_in_29_10;
wire x_in_29_11;
wire x_in_29_12;
wire x_in_29_13;
wire x_in_29_14;
wire x_in_29_15;
wire x_in_29_2;
wire x_in_29_3;
wire x_in_29_4;
wire x_in_29_5;
wire x_in_29_6;
wire x_in_29_7;
wire x_in_29_8;
wire x_in_29_9;
wire x_in_2_0;
wire x_in_2_1;
wire x_in_2_10;
wire x_in_2_11;
wire x_in_2_12;
wire x_in_2_13;
wire x_in_2_14;
wire x_in_2_15;
wire x_in_2_2;
wire x_in_2_3;
wire x_in_2_4;
wire x_in_2_5;
wire x_in_2_6;
wire x_in_2_7;
wire x_in_2_8;
wire x_in_2_9;
wire x_in_30_0;
wire x_in_30_1;
wire x_in_30_10;
wire x_in_30_11;
wire x_in_30_12;
wire x_in_30_13;
wire x_in_30_14;
wire x_in_30_15;
wire x_in_30_2;
wire x_in_30_3;
wire x_in_30_4;
wire x_in_30_5;
wire x_in_30_6;
wire x_in_30_7;
wire x_in_30_8;
wire x_in_30_9;
wire x_in_31_0;
wire x_in_31_1;
wire x_in_31_10;
wire x_in_31_11;
wire x_in_31_12;
wire x_in_31_13;
wire x_in_31_14;
wire x_in_31_15;
wire x_in_31_2;
wire x_in_31_3;
wire x_in_31_4;
wire x_in_31_5;
wire x_in_31_6;
wire x_in_31_7;
wire x_in_31_8;
wire x_in_31_9;
wire x_in_32_0;
wire x_in_32_1;
wire x_in_32_10;
wire x_in_32_11;
wire x_in_32_12;
wire x_in_32_13;
wire x_in_32_14;
wire x_in_32_15;
wire x_in_32_2;
wire x_in_32_3;
wire x_in_32_4;
wire x_in_32_5;
wire x_in_32_6;
wire x_in_32_7;
wire x_in_32_8;
wire x_in_32_9;
wire x_in_33_0;
wire x_in_33_1;
wire x_in_33_10;
wire x_in_33_11;
wire x_in_33_12;
wire x_in_33_13;
wire x_in_33_14;
wire x_in_33_15;
wire x_in_33_2;
wire x_in_33_3;
wire x_in_33_4;
wire x_in_33_5;
wire x_in_33_6;
wire x_in_33_7;
wire x_in_33_8;
wire x_in_33_9;
wire x_in_34_0;
wire x_in_34_1;
wire x_in_34_10;
wire x_in_34_11;
wire x_in_34_12;
wire x_in_34_13;
wire x_in_34_14;
wire x_in_34_15;
wire x_in_34_2;
wire x_in_34_3;
wire x_in_34_4;
wire x_in_34_5;
wire x_in_34_6;
wire x_in_34_7;
wire x_in_34_8;
wire x_in_34_9;
wire x_in_35_0;
wire x_in_35_1;
wire x_in_35_10;
wire x_in_35_11;
wire x_in_35_12;
wire x_in_35_13;
wire x_in_35_14;
wire x_in_35_15;
wire x_in_35_2;
wire x_in_35_3;
wire x_in_35_4;
wire x_in_35_5;
wire x_in_35_6;
wire x_in_35_7;
wire x_in_35_8;
wire x_in_35_9;
wire x_in_36_0;
wire x_in_36_1;
wire x_in_36_10;
wire x_in_36_11;
wire x_in_36_12;
wire x_in_36_13;
wire x_in_36_14;
wire x_in_36_15;
wire x_in_36_2;
wire x_in_36_3;
wire x_in_36_4;
wire x_in_36_5;
wire x_in_36_6;
wire x_in_36_7;
wire x_in_36_8;
wire x_in_36_9;
wire x_in_37_0;
wire x_in_37_1;
wire x_in_37_10;
wire x_in_37_11;
wire x_in_37_12;
wire x_in_37_13;
wire x_in_37_14;
wire x_in_37_15;
wire x_in_37_2;
wire x_in_37_3;
wire x_in_37_4;
wire x_in_37_5;
wire x_in_37_6;
wire x_in_37_7;
wire x_in_37_8;
wire x_in_37_9;
wire x_in_38_0;
wire x_in_38_1;
wire x_in_38_10;
wire x_in_38_11;
wire x_in_38_12;
wire x_in_38_13;
wire x_in_38_14;
wire x_in_38_15;
wire x_in_38_2;
wire x_in_38_3;
wire x_in_38_4;
wire x_in_38_5;
wire x_in_38_6;
wire x_in_38_7;
wire x_in_38_8;
wire x_in_38_9;
wire x_in_39_0;
wire x_in_39_1;
wire x_in_39_10;
wire x_in_39_11;
wire x_in_39_12;
wire x_in_39_13;
wire x_in_39_14;
wire x_in_39_15;
wire x_in_39_2;
wire x_in_39_3;
wire x_in_39_4;
wire x_in_39_5;
wire x_in_39_6;
wire x_in_39_7;
wire x_in_39_8;
wire x_in_39_9;
wire x_in_3_0;
wire x_in_3_1;
wire x_in_3_10;
wire x_in_3_11;
wire x_in_3_12;
wire x_in_3_13;
wire x_in_3_14;
wire x_in_3_15;
wire x_in_3_2;
wire x_in_3_3;
wire x_in_3_4;
wire x_in_3_5;
wire x_in_3_6;
wire x_in_3_7;
wire x_in_3_8;
wire x_in_3_9;
wire x_in_40_0;
wire x_in_40_1;
wire x_in_40_10;
wire x_in_40_11;
wire x_in_40_12;
wire x_in_40_13;
wire x_in_40_14;
wire x_in_40_15;
wire x_in_40_2;
wire x_in_40_3;
wire x_in_40_4;
wire x_in_40_5;
wire x_in_40_6;
wire x_in_40_7;
wire x_in_40_8;
wire x_in_40_9;
wire x_in_41_0;
wire x_in_41_1;
wire x_in_41_10;
wire x_in_41_11;
wire x_in_41_12;
wire x_in_41_13;
wire x_in_41_14;
wire x_in_41_15;
wire x_in_41_2;
wire x_in_41_3;
wire x_in_41_4;
wire x_in_41_5;
wire x_in_41_6;
wire x_in_41_7;
wire x_in_41_8;
wire x_in_41_9;
wire x_in_42_0;
wire x_in_42_1;
wire x_in_42_10;
wire x_in_42_11;
wire x_in_42_12;
wire x_in_42_13;
wire x_in_42_14;
wire x_in_42_15;
wire x_in_42_2;
wire x_in_42_3;
wire x_in_42_4;
wire x_in_42_5;
wire x_in_42_6;
wire x_in_42_7;
wire x_in_42_8;
wire x_in_42_9;
wire x_in_43_0;
wire x_in_43_1;
wire x_in_43_10;
wire x_in_43_11;
wire x_in_43_12;
wire x_in_43_13;
wire x_in_43_14;
wire x_in_43_15;
wire x_in_43_2;
wire x_in_43_3;
wire x_in_43_4;
wire x_in_43_5;
wire x_in_43_6;
wire x_in_43_7;
wire x_in_43_8;
wire x_in_43_9;
wire x_in_44_0;
wire x_in_44_1;
wire x_in_44_10;
wire x_in_44_11;
wire x_in_44_12;
wire x_in_44_13;
wire x_in_44_14;
wire x_in_44_15;
wire x_in_44_2;
wire x_in_44_3;
wire x_in_44_4;
wire x_in_44_5;
wire x_in_44_6;
wire x_in_44_7;
wire x_in_44_8;
wire x_in_44_9;
wire x_in_45_0;
wire x_in_45_1;
wire x_in_45_10;
wire x_in_45_11;
wire x_in_45_12;
wire x_in_45_13;
wire x_in_45_14;
wire x_in_45_15;
wire x_in_45_2;
wire x_in_45_3;
wire x_in_45_4;
wire x_in_45_5;
wire x_in_45_6;
wire x_in_45_7;
wire x_in_45_8;
wire x_in_45_9;
wire x_in_46_0;
wire x_in_46_1;
wire x_in_46_10;
wire x_in_46_11;
wire x_in_46_12;
wire x_in_46_13;
wire x_in_46_14;
wire x_in_46_15;
wire x_in_46_2;
wire x_in_46_3;
wire x_in_46_4;
wire x_in_46_5;
wire x_in_46_6;
wire x_in_46_7;
wire x_in_46_8;
wire x_in_46_9;
wire x_in_47_0;
wire x_in_47_1;
wire x_in_47_10;
wire x_in_47_11;
wire x_in_47_12;
wire x_in_47_13;
wire x_in_47_14;
wire x_in_47_15;
wire x_in_47_2;
wire x_in_47_3;
wire x_in_47_4;
wire x_in_47_5;
wire x_in_47_6;
wire x_in_47_7;
wire x_in_47_8;
wire x_in_47_9;
wire x_in_48_0;
wire x_in_48_1;
wire x_in_48_10;
wire x_in_48_11;
wire x_in_48_12;
wire x_in_48_13;
wire x_in_48_14;
wire x_in_48_15;
wire x_in_48_2;
wire x_in_48_3;
wire x_in_48_4;
wire x_in_48_5;
wire x_in_48_6;
wire x_in_48_7;
wire x_in_48_8;
wire x_in_48_9;
wire x_in_49_0;
wire x_in_49_1;
wire x_in_49_10;
wire x_in_49_11;
wire x_in_49_12;
wire x_in_49_13;
wire x_in_49_14;
wire x_in_49_15;
wire x_in_49_2;
wire x_in_49_3;
wire x_in_49_4;
wire x_in_49_5;
wire x_in_49_6;
wire x_in_49_7;
wire x_in_49_8;
wire x_in_49_9;
wire x_in_4_0;
wire x_in_4_1;
wire x_in_4_10;
wire x_in_4_11;
wire x_in_4_12;
wire x_in_4_13;
wire x_in_4_14;
wire x_in_4_15;
wire x_in_4_2;
wire x_in_4_3;
wire x_in_4_4;
wire x_in_4_5;
wire x_in_4_6;
wire x_in_4_7;
wire x_in_4_8;
wire x_in_4_9;
wire x_in_50_0;
wire x_in_50_1;
wire x_in_50_10;
wire x_in_50_11;
wire x_in_50_12;
wire x_in_50_13;
wire x_in_50_14;
wire x_in_50_15;
wire x_in_50_2;
wire x_in_50_3;
wire x_in_50_4;
wire x_in_50_5;
wire x_in_50_6;
wire x_in_50_7;
wire x_in_50_8;
wire x_in_50_9;
wire x_in_51_0;
wire x_in_51_1;
wire x_in_51_10;
wire x_in_51_11;
wire x_in_51_12;
wire x_in_51_13;
wire x_in_51_14;
wire x_in_51_15;
wire x_in_51_2;
wire x_in_51_3;
wire x_in_51_4;
wire x_in_51_5;
wire x_in_51_6;
wire x_in_51_7;
wire x_in_51_8;
wire x_in_51_9;
wire x_in_52_0;
wire x_in_52_1;
wire x_in_52_10;
wire x_in_52_11;
wire x_in_52_12;
wire x_in_52_13;
wire x_in_52_14;
wire x_in_52_15;
wire x_in_52_2;
wire x_in_52_3;
wire x_in_52_4;
wire x_in_52_5;
wire x_in_52_6;
wire x_in_52_7;
wire x_in_52_8;
wire x_in_52_9;
wire x_in_53_0;
wire x_in_53_1;
wire x_in_53_10;
wire x_in_53_11;
wire x_in_53_12;
wire x_in_53_13;
wire x_in_53_14;
wire x_in_53_15;
wire x_in_53_2;
wire x_in_53_3;
wire x_in_53_4;
wire x_in_53_5;
wire x_in_53_6;
wire x_in_53_7;
wire x_in_53_8;
wire x_in_53_9;
wire x_in_54_0;
wire x_in_54_1;
wire x_in_54_10;
wire x_in_54_11;
wire x_in_54_12;
wire x_in_54_13;
wire x_in_54_14;
wire x_in_54_15;
wire x_in_54_2;
wire x_in_54_3;
wire x_in_54_4;
wire x_in_54_5;
wire x_in_54_6;
wire x_in_54_7;
wire x_in_54_8;
wire x_in_54_9;
wire x_in_55_0;
wire x_in_55_1;
wire x_in_55_10;
wire x_in_55_11;
wire x_in_55_12;
wire x_in_55_13;
wire x_in_55_14;
wire x_in_55_15;
wire x_in_55_2;
wire x_in_55_3;
wire x_in_55_4;
wire x_in_55_5;
wire x_in_55_6;
wire x_in_55_7;
wire x_in_55_8;
wire x_in_55_9;
wire x_in_56_0;
wire x_in_56_1;
wire x_in_56_10;
wire x_in_56_11;
wire x_in_56_12;
wire x_in_56_13;
wire x_in_56_14;
wire x_in_56_15;
wire x_in_56_2;
wire x_in_56_3;
wire x_in_56_4;
wire x_in_56_5;
wire x_in_56_6;
wire x_in_56_7;
wire x_in_56_8;
wire x_in_56_9;
wire x_in_57_0;
wire x_in_57_1;
wire x_in_57_10;
wire x_in_57_11;
wire x_in_57_12;
wire x_in_57_13;
wire x_in_57_14;
wire x_in_57_15;
wire x_in_57_2;
wire x_in_57_3;
wire x_in_57_4;
wire x_in_57_5;
wire x_in_57_6;
wire x_in_57_7;
wire x_in_57_8;
wire x_in_57_9;
wire x_in_58_0;
wire x_in_58_1;
wire x_in_58_10;
wire x_in_58_11;
wire x_in_58_12;
wire x_in_58_13;
wire x_in_58_14;
wire x_in_58_15;
wire x_in_58_2;
wire x_in_58_3;
wire x_in_58_4;
wire x_in_58_5;
wire x_in_58_6;
wire x_in_58_7;
wire x_in_58_8;
wire x_in_58_9;
wire x_in_59_0;
wire x_in_59_1;
wire x_in_59_10;
wire x_in_59_11;
wire x_in_59_12;
wire x_in_59_13;
wire x_in_59_14;
wire x_in_59_15;
wire x_in_59_2;
wire x_in_59_3;
wire x_in_59_4;
wire x_in_59_5;
wire x_in_59_6;
wire x_in_59_7;
wire x_in_59_8;
wire x_in_59_9;
wire x_in_5_0;
wire x_in_5_1;
wire x_in_5_10;
wire x_in_5_11;
wire x_in_5_12;
wire x_in_5_13;
wire x_in_5_14;
wire x_in_5_15;
wire x_in_5_2;
wire x_in_5_3;
wire x_in_5_4;
wire x_in_5_5;
wire x_in_5_6;
wire x_in_5_7;
wire x_in_5_8;
wire x_in_5_9;
wire x_in_60_0;
wire x_in_60_1;
wire x_in_60_10;
wire x_in_60_11;
wire x_in_60_12;
wire x_in_60_13;
wire x_in_60_14;
wire x_in_60_15;
wire x_in_60_2;
wire x_in_60_3;
wire x_in_60_4;
wire x_in_60_5;
wire x_in_60_6;
wire x_in_60_7;
wire x_in_60_8;
wire x_in_60_9;
wire x_in_61_0;
wire x_in_61_1;
wire x_in_61_10;
wire x_in_61_11;
wire x_in_61_12;
wire x_in_61_13;
wire x_in_61_14;
wire x_in_61_15;
wire x_in_61_2;
wire x_in_61_3;
wire x_in_61_4;
wire x_in_61_5;
wire x_in_61_6;
wire x_in_61_7;
wire x_in_61_8;
wire x_in_61_9;
wire x_in_62_0;
wire x_in_62_1;
wire x_in_62_10;
wire x_in_62_11;
wire x_in_62_12;
wire x_in_62_13;
wire x_in_62_14;
wire x_in_62_15;
wire x_in_62_2;
wire x_in_62_3;
wire x_in_62_4;
wire x_in_62_5;
wire x_in_62_6;
wire x_in_62_7;
wire x_in_62_8;
wire x_in_62_9;
wire x_in_63_0;
wire x_in_63_1;
wire x_in_63_10;
wire x_in_63_11;
wire x_in_63_12;
wire x_in_63_13;
wire x_in_63_14;
wire x_in_63_15;
wire x_in_63_2;
wire x_in_63_3;
wire x_in_63_4;
wire x_in_63_5;
wire x_in_63_6;
wire x_in_63_7;
wire x_in_63_8;
wire x_in_63_9;
wire x_in_6_0;
wire x_in_6_1;
wire x_in_6_10;
wire x_in_6_11;
wire x_in_6_12;
wire x_in_6_13;
wire x_in_6_14;
wire x_in_6_15;
wire x_in_6_2;
wire x_in_6_3;
wire x_in_6_4;
wire x_in_6_5;
wire x_in_6_6;
wire x_in_6_7;
wire x_in_6_8;
wire x_in_6_9;
wire x_in_7_0;
wire x_in_7_1;
wire x_in_7_10;
wire x_in_7_11;
wire x_in_7_12;
wire x_in_7_13;
wire x_in_7_14;
wire x_in_7_15;
wire x_in_7_2;
wire x_in_7_3;
wire x_in_7_4;
wire x_in_7_5;
wire x_in_7_6;
wire x_in_7_7;
wire x_in_7_8;
wire x_in_7_9;
wire x_in_8_0;
wire x_in_8_1;
wire x_in_8_10;
wire x_in_8_11;
wire x_in_8_12;
wire x_in_8_13;
wire x_in_8_14;
wire x_in_8_15;
wire x_in_8_2;
wire x_in_8_3;
wire x_in_8_4;
wire x_in_8_5;
wire x_in_8_6;
wire x_in_8_7;
wire x_in_8_8;
wire x_in_8_9;
wire x_in_9_0;
wire x_in_9_1;
wire x_in_9_10;
wire x_in_9_11;
wire x_in_9_12;
wire x_in_9_13;
wire x_in_9_14;
wire x_in_9_15;
wire x_in_9_2;
wire x_in_9_3;
wire x_in_9_4;
wire x_in_9_5;
wire x_in_9_6;
wire x_in_9_7;
wire x_in_9_8;
wire x_in_9_9;
wire x_out_0_0;
wire x_out_0_1;
wire x_out_0_10;
wire x_out_0_11;
wire x_out_0_12;
wire x_out_0_13;
wire x_out_0_14;
wire x_out_0_15;
wire x_out_0_2;
wire x_out_0_3;
wire x_out_0_4;
wire x_out_0_5;
wire x_out_0_6;
wire x_out_0_7;
wire x_out_0_8;
wire x_out_0_9;
wire x_out_10_0;
wire x_out_10_1;
wire x_out_10_10;
wire x_out_10_11;
wire x_out_10_12;
wire x_out_10_13;
wire x_out_10_14;
wire x_out_10_15;
wire x_out_10_18;
wire x_out_10_19;
wire x_out_10_2;
wire x_out_10_20;
wire x_out_10_21;
wire x_out_10_22;
wire x_out_10_23;
wire x_out_10_24;
wire x_out_10_25;
wire x_out_10_26;
wire x_out_10_27;
wire x_out_10_28;
wire x_out_10_29;
wire x_out_10_3;
wire x_out_10_30;
wire x_out_10_31;
wire x_out_10_32;
wire x_out_10_33;
wire x_out_10_4;
wire x_out_10_5;
wire x_out_10_6;
wire x_out_10_7;
wire x_out_10_8;
wire x_out_10_9;
wire x_out_11_0;
wire x_out_11_1;
wire x_out_11_10;
wire x_out_11_11;
wire x_out_11_12;
wire x_out_11_13;
wire x_out_11_14;
wire x_out_11_15;
wire x_out_11_18;
wire x_out_11_19;
wire x_out_11_2;
wire x_out_11_20;
wire x_out_11_21;
wire x_out_11_22;
wire x_out_11_23;
wire x_out_11_24;
wire x_out_11_25;
wire x_out_11_26;
wire x_out_11_27;
wire x_out_11_28;
wire x_out_11_29;
wire x_out_11_3;
wire x_out_11_30;
wire x_out_11_31;
wire x_out_11_32;
wire x_out_11_33;
wire x_out_11_4;
wire x_out_11_5;
wire x_out_11_6;
wire x_out_11_7;
wire x_out_11_8;
wire x_out_11_9;
wire x_out_12_0;
wire x_out_12_1;
wire x_out_12_10;
wire x_out_12_11;
wire x_out_12_12;
wire x_out_12_13;
wire x_out_12_14;
wire x_out_12_15;
wire x_out_12_18;
wire x_out_12_19;
wire x_out_12_2;
wire x_out_12_20;
wire x_out_12_21;
wire x_out_12_22;
wire x_out_12_23;
wire x_out_12_24;
wire x_out_12_25;
wire x_out_12_26;
wire x_out_12_27;
wire x_out_12_28;
wire x_out_12_29;
wire x_out_12_3;
wire x_out_12_30;
wire x_out_12_31;
wire x_out_12_32;
wire x_out_12_33;
wire x_out_12_4;
wire x_out_12_5;
wire x_out_12_6;
wire x_out_12_7;
wire x_out_12_8;
wire x_out_12_9;
wire x_out_13_0;
wire x_out_13_1;
wire x_out_13_10;
wire x_out_13_11;
wire x_out_13_12;
wire x_out_13_13;
wire x_out_13_14;
wire x_out_13_15;
wire x_out_13_18;
wire x_out_13_19;
wire x_out_13_2;
wire x_out_13_20;
wire x_out_13_21;
wire x_out_13_22;
wire x_out_13_23;
wire x_out_13_24;
wire x_out_13_25;
wire x_out_13_26;
wire x_out_13_27;
wire x_out_13_28;
wire x_out_13_29;
wire x_out_13_3;
wire x_out_13_30;
wire x_out_13_31;
wire x_out_13_32;
wire x_out_13_33;
wire x_out_13_4;
wire x_out_13_5;
wire x_out_13_6;
wire x_out_13_7;
wire x_out_13_8;
wire x_out_13_9;
wire x_out_14_0;
wire x_out_14_1;
wire x_out_14_10;
wire x_out_14_11;
wire x_out_14_12;
wire x_out_14_13;
wire x_out_14_14;
wire x_out_14_15;
wire x_out_14_18;
wire x_out_14_19;
wire x_out_14_2;
wire x_out_14_20;
wire x_out_14_21;
wire x_out_14_22;
wire x_out_14_23;
wire x_out_14_24;
wire x_out_14_25;
wire x_out_14_26;
wire x_out_14_27;
wire x_out_14_28;
wire x_out_14_29;
wire x_out_14_3;
wire x_out_14_30;
wire x_out_14_31;
wire x_out_14_32;
wire x_out_14_33;
wire x_out_14_4;
wire x_out_14_5;
wire x_out_14_6;
wire x_out_14_7;
wire x_out_14_8;
wire x_out_14_9;
wire x_out_15_0;
wire x_out_15_1;
wire x_out_15_10;
wire x_out_15_11;
wire x_out_15_12;
wire x_out_15_13;
wire x_out_15_14;
wire x_out_15_15;
wire x_out_15_18;
wire x_out_15_19;
wire x_out_15_2;
wire x_out_15_20;
wire x_out_15_21;
wire x_out_15_22;
wire x_out_15_23;
wire x_out_15_24;
wire x_out_15_25;
wire x_out_15_26;
wire x_out_15_27;
wire x_out_15_28;
wire x_out_15_29;
wire x_out_15_3;
wire x_out_15_30;
wire x_out_15_31;
wire x_out_15_32;
wire x_out_15_33;
wire x_out_15_4;
wire x_out_15_5;
wire x_out_15_6;
wire x_out_15_7;
wire x_out_15_8;
wire x_out_15_9;
wire x_out_16_0;
wire x_out_16_1;
wire x_out_16_10;
wire x_out_16_11;
wire x_out_16_12;
wire x_out_16_13;
wire x_out_16_14;
wire x_out_16_15;
wire x_out_16_18;
wire x_out_16_19;
wire x_out_16_2;
wire x_out_16_20;
wire x_out_16_21;
wire x_out_16_22;
wire x_out_16_23;
wire x_out_16_24;
wire x_out_16_25;
wire x_out_16_26;
wire x_out_16_27;
wire x_out_16_28;
wire x_out_16_29;
wire x_out_16_3;
wire x_out_16_30;
wire x_out_16_31;
wire x_out_16_32;
wire x_out_16_33;
wire x_out_16_4;
wire x_out_16_5;
wire x_out_16_6;
wire x_out_16_7;
wire x_out_16_8;
wire x_out_16_9;
wire x_out_17_0;
wire x_out_17_1;
wire x_out_17_10;
wire x_out_17_11;
wire x_out_17_12;
wire x_out_17_13;
wire x_out_17_14;
wire x_out_17_15;
wire x_out_17_18;
wire x_out_17_19;
wire x_out_17_2;
wire x_out_17_20;
wire x_out_17_21;
wire x_out_17_22;
wire x_out_17_23;
wire x_out_17_24;
wire x_out_17_25;
wire x_out_17_26;
wire x_out_17_27;
wire x_out_17_28;
wire x_out_17_29;
wire x_out_17_3;
wire x_out_17_30;
wire x_out_17_31;
wire x_out_17_32;
wire x_out_17_33;
wire x_out_17_4;
wire x_out_17_5;
wire x_out_17_6;
wire x_out_17_7;
wire x_out_17_8;
wire x_out_17_9;
wire x_out_18_0;
wire x_out_18_1;
wire x_out_18_10;
wire x_out_18_11;
wire x_out_18_12;
wire x_out_18_13;
wire x_out_18_14;
wire x_out_18_15;
wire x_out_18_18;
wire x_out_18_19;
wire x_out_18_2;
wire x_out_18_20;
wire x_out_18_21;
wire x_out_18_22;
wire x_out_18_23;
wire x_out_18_24;
wire x_out_18_25;
wire x_out_18_26;
wire x_out_18_27;
wire x_out_18_28;
wire x_out_18_29;
wire x_out_18_3;
wire x_out_18_30;
wire x_out_18_31;
wire x_out_18_32;
wire x_out_18_33;
wire x_out_18_4;
wire x_out_18_5;
wire x_out_18_6;
wire x_out_18_7;
wire x_out_18_8;
wire x_out_18_9;
wire x_out_19_0;
wire x_out_19_1;
wire x_out_19_10;
wire x_out_19_11;
wire x_out_19_12;
wire x_out_19_13;
wire x_out_19_14;
wire x_out_19_15;
wire x_out_19_18;
wire x_out_19_19;
wire x_out_19_2;
wire x_out_19_20;
wire x_out_19_21;
wire x_out_19_22;
wire x_out_19_23;
wire x_out_19_24;
wire x_out_19_25;
wire x_out_19_26;
wire x_out_19_27;
wire x_out_19_28;
wire x_out_19_29;
wire x_out_19_3;
wire x_out_19_30;
wire x_out_19_31;
wire x_out_19_32;
wire x_out_19_33;
wire x_out_19_4;
wire x_out_19_5;
wire x_out_19_6;
wire x_out_19_7;
wire x_out_19_8;
wire x_out_19_9;
wire x_out_1_0;
wire x_out_1_1;
wire x_out_1_10;
wire x_out_1_11;
wire x_out_1_12;
wire x_out_1_13;
wire x_out_1_14;
wire x_out_1_15;
wire x_out_1_18;
wire x_out_1_19;
wire x_out_1_2;
wire x_out_1_20;
wire x_out_1_21;
wire x_out_1_22;
wire x_out_1_23;
wire x_out_1_24;
wire x_out_1_25;
wire x_out_1_26;
wire x_out_1_27;
wire x_out_1_28;
wire x_out_1_29;
wire x_out_1_3;
wire x_out_1_30;
wire x_out_1_31;
wire x_out_1_32;
wire x_out_1_33;
wire x_out_1_4;
wire x_out_1_5;
wire x_out_1_6;
wire x_out_1_7;
wire x_out_1_8;
wire x_out_1_9;
wire x_out_20_0;
wire x_out_20_1;
wire x_out_20_10;
wire x_out_20_11;
wire x_out_20_12;
wire x_out_20_13;
wire x_out_20_14;
wire x_out_20_15;
wire x_out_20_2;
wire x_out_20_3;
wire x_out_20_4;
wire x_out_20_5;
wire x_out_20_6;
wire x_out_20_7;
wire x_out_20_8;
wire x_out_20_9;
wire x_out_21_0;
wire x_out_21_1;
wire x_out_21_10;
wire x_out_21_11;
wire x_out_21_12;
wire x_out_21_13;
wire x_out_21_14;
wire x_out_21_15;
wire x_out_21_18;
wire x_out_21_19;
wire x_out_21_2;
wire x_out_21_20;
wire x_out_21_21;
wire x_out_21_22;
wire x_out_21_23;
wire x_out_21_24;
wire x_out_21_25;
wire x_out_21_26;
wire x_out_21_27;
wire x_out_21_28;
wire x_out_21_29;
wire x_out_21_3;
wire x_out_21_30;
wire x_out_21_31;
wire x_out_21_32;
wire x_out_21_33;
wire x_out_21_4;
wire x_out_21_5;
wire x_out_21_6;
wire x_out_21_7;
wire x_out_21_8;
wire x_out_21_9;
wire x_out_22_0;
wire x_out_22_1;
wire x_out_22_10;
wire x_out_22_11;
wire x_out_22_12;
wire x_out_22_13;
wire x_out_22_14;
wire x_out_22_15;
wire x_out_22_18;
wire x_out_22_19;
wire x_out_22_2;
wire x_out_22_20;
wire x_out_22_21;
wire x_out_22_22;
wire x_out_22_23;
wire x_out_22_24;
wire x_out_22_25;
wire x_out_22_26;
wire x_out_22_27;
wire x_out_22_28;
wire x_out_22_29;
wire x_out_22_3;
wire x_out_22_30;
wire x_out_22_31;
wire x_out_22_32;
wire x_out_22_33;
wire x_out_22_4;
wire x_out_22_5;
wire x_out_22_6;
wire x_out_22_7;
wire x_out_22_8;
wire x_out_22_9;
wire x_out_23_0;
wire x_out_23_1;
wire x_out_23_10;
wire x_out_23_11;
wire x_out_23_12;
wire x_out_23_13;
wire x_out_23_14;
wire x_out_23_15;
wire x_out_23_18;
wire x_out_23_19;
wire x_out_23_2;
wire x_out_23_20;
wire x_out_23_21;
wire x_out_23_22;
wire x_out_23_23;
wire x_out_23_24;
wire x_out_23_25;
wire x_out_23_26;
wire x_out_23_27;
wire x_out_23_28;
wire x_out_23_29;
wire x_out_23_3;
wire x_out_23_30;
wire x_out_23_31;
wire x_out_23_32;
wire x_out_23_33;
wire x_out_23_4;
wire x_out_23_5;
wire x_out_23_6;
wire x_out_23_7;
wire x_out_23_8;
wire x_out_23_9;
wire x_out_24_0;
wire x_out_24_1;
wire x_out_24_10;
wire x_out_24_11;
wire x_out_24_12;
wire x_out_24_13;
wire x_out_24_14;
wire x_out_24_15;
wire x_out_24_18;
wire x_out_24_19;
wire x_out_24_2;
wire x_out_24_20;
wire x_out_24_21;
wire x_out_24_22;
wire x_out_24_23;
wire x_out_24_24;
wire x_out_24_25;
wire x_out_24_26;
wire x_out_24_27;
wire x_out_24_28;
wire x_out_24_29;
wire x_out_24_3;
wire x_out_24_30;
wire x_out_24_31;
wire x_out_24_32;
wire x_out_24_33;
wire x_out_24_4;
wire x_out_24_5;
wire x_out_24_6;
wire x_out_24_7;
wire x_out_24_8;
wire x_out_24_9;
wire x_out_25_0;
wire x_out_25_1;
wire x_out_25_10;
wire x_out_25_11;
wire x_out_25_12;
wire x_out_25_13;
wire x_out_25_14;
wire x_out_25_15;
wire x_out_25_18;
wire x_out_25_19;
wire x_out_25_2;
wire x_out_25_20;
wire x_out_25_21;
wire x_out_25_22;
wire x_out_25_23;
wire x_out_25_24;
wire x_out_25_25;
wire x_out_25_26;
wire x_out_25_27;
wire x_out_25_28;
wire x_out_25_29;
wire x_out_25_3;
wire x_out_25_30;
wire x_out_25_31;
wire x_out_25_32;
wire x_out_25_33;
wire x_out_25_4;
wire x_out_25_5;
wire x_out_25_6;
wire x_out_25_7;
wire x_out_25_8;
wire x_out_25_9;
wire x_out_26_0;
wire x_out_26_1;
wire x_out_26_10;
wire x_out_26_11;
wire x_out_26_12;
wire x_out_26_13;
wire x_out_26_14;
wire x_out_26_15;
wire x_out_26_18;
wire x_out_26_19;
wire x_out_26_2;
wire x_out_26_20;
wire x_out_26_21;
wire x_out_26_22;
wire x_out_26_23;
wire x_out_26_24;
wire x_out_26_25;
wire x_out_26_26;
wire x_out_26_27;
wire x_out_26_28;
wire x_out_26_29;
wire x_out_26_3;
wire x_out_26_30;
wire x_out_26_31;
wire x_out_26_32;
wire x_out_26_33;
wire x_out_26_4;
wire x_out_26_5;
wire x_out_26_6;
wire x_out_26_7;
wire x_out_26_8;
wire x_out_26_9;
wire x_out_27_0;
wire x_out_27_1;
wire x_out_27_10;
wire x_out_27_11;
wire x_out_27_12;
wire x_out_27_13;
wire x_out_27_14;
wire x_out_27_15;
wire x_out_27_18;
wire x_out_27_19;
wire x_out_27_2;
wire x_out_27_20;
wire x_out_27_21;
wire x_out_27_22;
wire x_out_27_23;
wire x_out_27_24;
wire x_out_27_25;
wire x_out_27_26;
wire x_out_27_27;
wire x_out_27_28;
wire x_out_27_29;
wire x_out_27_3;
wire x_out_27_30;
wire x_out_27_31;
wire x_out_27_32;
wire x_out_27_33;
wire x_out_27_4;
wire x_out_27_5;
wire x_out_27_6;
wire x_out_27_7;
wire x_out_27_8;
wire x_out_27_9;
wire x_out_28_0;
wire x_out_28_1;
wire x_out_28_10;
wire x_out_28_11;
wire x_out_28_12;
wire x_out_28_13;
wire x_out_28_14;
wire x_out_28_15;
wire x_out_28_18;
wire x_out_28_19;
wire x_out_28_2;
wire x_out_28_20;
wire x_out_28_21;
wire x_out_28_22;
wire x_out_28_23;
wire x_out_28_24;
wire x_out_28_25;
wire x_out_28_26;
wire x_out_28_27;
wire x_out_28_28;
wire x_out_28_29;
wire x_out_28_3;
wire x_out_28_30;
wire x_out_28_31;
wire x_out_28_32;
wire x_out_28_33;
wire x_out_28_4;
wire x_out_28_5;
wire x_out_28_6;
wire x_out_28_7;
wire x_out_28_8;
wire x_out_28_9;
wire x_out_29_0;
wire x_out_29_1;
wire x_out_29_10;
wire x_out_29_11;
wire x_out_29_12;
wire x_out_29_13;
wire x_out_29_14;
wire x_out_29_15;
wire x_out_29_18;
wire x_out_29_19;
wire x_out_29_2;
wire x_out_29_20;
wire x_out_29_21;
wire x_out_29_22;
wire x_out_29_23;
wire x_out_29_24;
wire x_out_29_25;
wire x_out_29_26;
wire x_out_29_27;
wire x_out_29_28;
wire x_out_29_29;
wire x_out_29_3;
wire x_out_29_30;
wire x_out_29_31;
wire x_out_29_32;
wire x_out_29_33;
wire x_out_29_4;
wire x_out_29_5;
wire x_out_29_6;
wire x_out_29_7;
wire x_out_29_8;
wire x_out_29_9;
wire x_out_2_0;
wire x_out_2_1;
wire x_out_2_10;
wire x_out_2_11;
wire x_out_2_12;
wire x_out_2_13;
wire x_out_2_14;
wire x_out_2_15;
wire x_out_2_18;
wire x_out_2_19;
wire x_out_2_2;
wire x_out_2_20;
wire x_out_2_21;
wire x_out_2_22;
wire x_out_2_23;
wire x_out_2_24;
wire x_out_2_25;
wire x_out_2_26;
wire x_out_2_27;
wire x_out_2_28;
wire x_out_2_29;
wire x_out_2_3;
wire x_out_2_30;
wire x_out_2_31;
wire x_out_2_32;
wire x_out_2_33;
wire x_out_2_4;
wire x_out_2_5;
wire x_out_2_6;
wire x_out_2_7;
wire x_out_2_8;
wire x_out_2_9;
wire x_out_30_0;
wire x_out_30_1;
wire x_out_30_10;
wire x_out_30_11;
wire x_out_30_12;
wire x_out_30_13;
wire x_out_30_14;
wire x_out_30_15;
wire x_out_30_18;
wire x_out_30_19;
wire x_out_30_2;
wire x_out_30_20;
wire x_out_30_21;
wire x_out_30_22;
wire x_out_30_23;
wire x_out_30_24;
wire x_out_30_25;
wire x_out_30_26;
wire x_out_30_27;
wire x_out_30_28;
wire x_out_30_29;
wire x_out_30_3;
wire x_out_30_30;
wire x_out_30_31;
wire x_out_30_32;
wire x_out_30_33;
wire x_out_30_4;
wire x_out_30_5;
wire x_out_30_6;
wire x_out_30_7;
wire x_out_30_8;
wire x_out_30_9;
wire x_out_31_0;
wire x_out_31_1;
wire x_out_31_10;
wire x_out_31_11;
wire x_out_31_12;
wire x_out_31_13;
wire x_out_31_14;
wire x_out_31_15;
wire x_out_31_18;
wire x_out_31_19;
wire x_out_31_2;
wire x_out_31_20;
wire x_out_31_21;
wire x_out_31_22;
wire x_out_31_23;
wire x_out_31_24;
wire x_out_31_25;
wire x_out_31_26;
wire x_out_31_27;
wire x_out_31_28;
wire x_out_31_29;
wire x_out_31_3;
wire x_out_31_30;
wire x_out_31_31;
wire x_out_31_32;
wire x_out_31_33;
wire x_out_31_4;
wire x_out_31_5;
wire x_out_31_6;
wire x_out_31_7;
wire x_out_31_8;
wire x_out_31_9;
wire x_out_32_0;
wire x_out_32_1;
wire x_out_32_10;
wire x_out_32_11;
wire x_out_32_12;
wire x_out_32_13;
wire x_out_32_14;
wire x_out_32_15;
wire x_out_32_2;
wire x_out_32_3;
wire x_out_32_4;
wire x_out_32_5;
wire x_out_32_6;
wire x_out_32_7;
wire x_out_32_8;
wire x_out_32_9;
wire x_out_33_0;
wire x_out_33_1;
wire x_out_33_10;
wire x_out_33_11;
wire x_out_33_12;
wire x_out_33_13;
wire x_out_33_14;
wire x_out_33_15;
wire x_out_33_18;
wire x_out_33_19;
wire x_out_33_2;
wire x_out_33_20;
wire x_out_33_21;
wire x_out_33_22;
wire x_out_33_23;
wire x_out_33_24;
wire x_out_33_25;
wire x_out_33_26;
wire x_out_33_27;
wire x_out_33_28;
wire x_out_33_29;
wire x_out_33_3;
wire x_out_33_30;
wire x_out_33_31;
wire x_out_33_32;
wire x_out_33_33;
wire x_out_33_4;
wire x_out_33_5;
wire x_out_33_6;
wire x_out_33_7;
wire x_out_33_8;
wire x_out_33_9;
wire x_out_34_0;
wire x_out_34_1;
wire x_out_34_10;
wire x_out_34_11;
wire x_out_34_12;
wire x_out_34_13;
wire x_out_34_14;
wire x_out_34_15;
wire x_out_34_18;
wire x_out_34_19;
wire x_out_34_2;
wire x_out_34_20;
wire x_out_34_21;
wire x_out_34_22;
wire x_out_34_23;
wire x_out_34_24;
wire x_out_34_25;
wire x_out_34_26;
wire x_out_34_27;
wire x_out_34_28;
wire x_out_34_29;
wire x_out_34_3;
wire x_out_34_30;
wire x_out_34_31;
wire x_out_34_32;
wire x_out_34_33;
wire x_out_34_4;
wire x_out_34_5;
wire x_out_34_6;
wire x_out_34_7;
wire x_out_34_8;
wire x_out_34_9;
wire x_out_35_0;
wire x_out_35_1;
wire x_out_35_10;
wire x_out_35_11;
wire x_out_35_12;
wire x_out_35_13;
wire x_out_35_14;
wire x_out_35_15;
wire x_out_35_18;
wire x_out_35_19;
wire x_out_35_2;
wire x_out_35_20;
wire x_out_35_21;
wire x_out_35_22;
wire x_out_35_23;
wire x_out_35_24;
wire x_out_35_25;
wire x_out_35_26;
wire x_out_35_27;
wire x_out_35_28;
wire x_out_35_29;
wire x_out_35_3;
wire x_out_35_30;
wire x_out_35_31;
wire x_out_35_32;
wire x_out_35_33;
wire x_out_35_4;
wire x_out_35_5;
wire x_out_35_6;
wire x_out_35_7;
wire x_out_35_8;
wire x_out_35_9;
wire x_out_36_0;
wire x_out_36_1;
wire x_out_36_10;
wire x_out_36_11;
wire x_out_36_12;
wire x_out_36_13;
wire x_out_36_14;
wire x_out_36_15;
wire x_out_36_18;
wire x_out_36_19;
wire x_out_36_2;
wire x_out_36_20;
wire x_out_36_21;
wire x_out_36_22;
wire x_out_36_23;
wire x_out_36_24;
wire x_out_36_25;
wire x_out_36_26;
wire x_out_36_27;
wire x_out_36_28;
wire x_out_36_29;
wire x_out_36_3;
wire x_out_36_30;
wire x_out_36_31;
wire x_out_36_32;
wire x_out_36_33;
wire x_out_36_4;
wire x_out_36_5;
wire x_out_36_6;
wire x_out_36_7;
wire x_out_36_8;
wire x_out_36_9;
wire x_out_37_0;
wire x_out_37_1;
wire x_out_37_10;
wire x_out_37_11;
wire x_out_37_12;
wire x_out_37_13;
wire x_out_37_14;
wire x_out_37_15;
wire x_out_37_18;
wire x_out_37_19;
wire x_out_37_2;
wire x_out_37_20;
wire x_out_37_21;
wire x_out_37_22;
wire x_out_37_23;
wire x_out_37_24;
wire x_out_37_25;
wire x_out_37_26;
wire x_out_37_27;
wire x_out_37_28;
wire x_out_37_29;
wire x_out_37_3;
wire x_out_37_30;
wire x_out_37_31;
wire x_out_37_32;
wire x_out_37_33;
wire x_out_37_4;
wire x_out_37_5;
wire x_out_37_6;
wire x_out_37_7;
wire x_out_37_8;
wire x_out_37_9;
wire x_out_38_0;
wire x_out_38_1;
wire x_out_38_10;
wire x_out_38_11;
wire x_out_38_12;
wire x_out_38_13;
wire x_out_38_14;
wire x_out_38_15;
wire x_out_38_18;
wire x_out_38_19;
wire x_out_38_2;
wire x_out_38_20;
wire x_out_38_21;
wire x_out_38_22;
wire x_out_38_23;
wire x_out_38_24;
wire x_out_38_25;
wire x_out_38_26;
wire x_out_38_27;
wire x_out_38_28;
wire x_out_38_29;
wire x_out_38_3;
wire x_out_38_30;
wire x_out_38_31;
wire x_out_38_32;
wire x_out_38_33;
wire x_out_38_4;
wire x_out_38_5;
wire x_out_38_6;
wire x_out_38_7;
wire x_out_38_8;
wire x_out_38_9;
wire x_out_39_0;
wire x_out_39_1;
wire x_out_39_10;
wire x_out_39_11;
wire x_out_39_12;
wire x_out_39_13;
wire x_out_39_14;
wire x_out_39_15;
wire x_out_39_18;
wire x_out_39_19;
wire x_out_39_2;
wire x_out_39_20;
wire x_out_39_21;
wire x_out_39_22;
wire x_out_39_23;
wire x_out_39_24;
wire x_out_39_25;
wire x_out_39_26;
wire x_out_39_27;
wire x_out_39_28;
wire x_out_39_29;
wire x_out_39_3;
wire x_out_39_30;
wire x_out_39_31;
wire x_out_39_32;
wire x_out_39_33;
wire x_out_39_4;
wire x_out_39_5;
wire x_out_39_6;
wire x_out_39_7;
wire x_out_39_8;
wire x_out_39_9;
wire x_out_3_0;
wire x_out_3_1;
wire x_out_3_10;
wire x_out_3_11;
wire x_out_3_12;
wire x_out_3_13;
wire x_out_3_14;
wire x_out_3_15;
wire x_out_3_18;
wire x_out_3_19;
wire x_out_3_2;
wire x_out_3_20;
wire x_out_3_21;
wire x_out_3_22;
wire x_out_3_23;
wire x_out_3_24;
wire x_out_3_25;
wire x_out_3_26;
wire x_out_3_27;
wire x_out_3_28;
wire x_out_3_29;
wire x_out_3_3;
wire x_out_3_30;
wire x_out_3_31;
wire x_out_3_32;
wire x_out_3_33;
wire x_out_3_4;
wire x_out_3_5;
wire x_out_3_6;
wire x_out_3_7;
wire x_out_3_8;
wire x_out_3_9;
wire x_out_40_0;
wire x_out_40_1;
wire x_out_40_10;
wire x_out_40_11;
wire x_out_40_12;
wire x_out_40_13;
wire x_out_40_14;
wire x_out_40_15;
wire x_out_40_18;
wire x_out_40_19;
wire x_out_40_2;
wire x_out_40_20;
wire x_out_40_21;
wire x_out_40_22;
wire x_out_40_23;
wire x_out_40_24;
wire x_out_40_25;
wire x_out_40_26;
wire x_out_40_27;
wire x_out_40_28;
wire x_out_40_29;
wire x_out_40_3;
wire x_out_40_30;
wire x_out_40_31;
wire x_out_40_32;
wire x_out_40_33;
wire x_out_40_4;
wire x_out_40_5;
wire x_out_40_6;
wire x_out_40_7;
wire x_out_40_8;
wire x_out_40_9;
wire x_out_41_0;
wire x_out_41_1;
wire x_out_41_10;
wire x_out_41_11;
wire x_out_41_12;
wire x_out_41_13;
wire x_out_41_14;
wire x_out_41_15;
wire x_out_41_18;
wire x_out_41_19;
wire x_out_41_2;
wire x_out_41_20;
wire x_out_41_21;
wire x_out_41_22;
wire x_out_41_23;
wire x_out_41_24;
wire x_out_41_25;
wire x_out_41_26;
wire x_out_41_27;
wire x_out_41_28;
wire x_out_41_29;
wire x_out_41_3;
wire x_out_41_30;
wire x_out_41_31;
wire x_out_41_32;
wire x_out_41_33;
wire x_out_41_4;
wire x_out_41_5;
wire x_out_41_6;
wire x_out_41_7;
wire x_out_41_8;
wire x_out_41_9;
wire x_out_42_0;
wire x_out_42_1;
wire x_out_42_10;
wire x_out_42_11;
wire x_out_42_12;
wire x_out_42_13;
wire x_out_42_14;
wire x_out_42_15;
wire x_out_42_18;
wire x_out_42_19;
wire x_out_42_2;
wire x_out_42_20;
wire x_out_42_21;
wire x_out_42_22;
wire x_out_42_23;
wire x_out_42_24;
wire x_out_42_25;
wire x_out_42_26;
wire x_out_42_27;
wire x_out_42_28;
wire x_out_42_29;
wire x_out_42_3;
wire x_out_42_30;
wire x_out_42_31;
wire x_out_42_32;
wire x_out_42_33;
wire x_out_42_4;
wire x_out_42_5;
wire x_out_42_6;
wire x_out_42_7;
wire x_out_42_8;
wire x_out_42_9;
wire x_out_43_0;
wire x_out_43_1;
wire x_out_43_10;
wire x_out_43_11;
wire x_out_43_12;
wire x_out_43_13;
wire x_out_43_14;
wire x_out_43_15;
wire x_out_43_18;
wire x_out_43_19;
wire x_out_43_2;
wire x_out_43_20;
wire x_out_43_21;
wire x_out_43_22;
wire x_out_43_23;
wire x_out_43_24;
wire x_out_43_25;
wire x_out_43_26;
wire x_out_43_27;
wire x_out_43_28;
wire x_out_43_29;
wire x_out_43_3;
wire x_out_43_30;
wire x_out_43_31;
wire x_out_43_32;
wire x_out_43_33;
wire x_out_43_4;
wire x_out_43_5;
wire x_out_43_6;
wire x_out_43_7;
wire x_out_43_8;
wire x_out_43_9;
wire x_out_44_0;
wire x_out_44_1;
wire x_out_44_10;
wire x_out_44_11;
wire x_out_44_12;
wire x_out_44_13;
wire x_out_44_14;
wire x_out_44_15;
wire x_out_44_18;
wire x_out_44_19;
wire x_out_44_2;
wire x_out_44_20;
wire x_out_44_21;
wire x_out_44_22;
wire x_out_44_23;
wire x_out_44_24;
wire x_out_44_25;
wire x_out_44_26;
wire x_out_44_27;
wire x_out_44_28;
wire x_out_44_29;
wire x_out_44_3;
wire x_out_44_30;
wire x_out_44_31;
wire x_out_44_32;
wire x_out_44_33;
wire x_out_44_4;
wire x_out_44_5;
wire x_out_44_6;
wire x_out_44_7;
wire x_out_44_8;
wire x_out_44_9;
wire x_out_45_0;
wire x_out_45_1;
wire x_out_45_10;
wire x_out_45_11;
wire x_out_45_12;
wire x_out_45_13;
wire x_out_45_14;
wire x_out_45_15;
wire x_out_45_18;
wire x_out_45_19;
wire x_out_45_2;
wire x_out_45_20;
wire x_out_45_21;
wire x_out_45_22;
wire x_out_45_23;
wire x_out_45_24;
wire x_out_45_25;
wire x_out_45_26;
wire x_out_45_27;
wire x_out_45_28;
wire x_out_45_29;
wire x_out_45_3;
wire x_out_45_30;
wire x_out_45_31;
wire x_out_45_32;
wire x_out_45_33;
wire x_out_45_4;
wire x_out_45_5;
wire x_out_45_6;
wire x_out_45_7;
wire x_out_45_8;
wire x_out_45_9;
wire x_out_46_0;
wire x_out_46_1;
wire x_out_46_10;
wire x_out_46_11;
wire x_out_46_12;
wire x_out_46_13;
wire x_out_46_14;
wire x_out_46_15;
wire x_out_46_18;
wire x_out_46_19;
wire x_out_46_2;
wire x_out_46_20;
wire x_out_46_21;
wire x_out_46_22;
wire x_out_46_23;
wire x_out_46_24;
wire x_out_46_25;
wire x_out_46_26;
wire x_out_46_27;
wire x_out_46_28;
wire x_out_46_29;
wire x_out_46_3;
wire x_out_46_30;
wire x_out_46_31;
wire x_out_46_32;
wire x_out_46_33;
wire x_out_46_4;
wire x_out_46_5;
wire x_out_46_6;
wire x_out_46_7;
wire x_out_46_8;
wire x_out_46_9;
wire x_out_47_0;
wire x_out_47_1;
wire x_out_47_10;
wire x_out_47_11;
wire x_out_47_12;
wire x_out_47_13;
wire x_out_47_14;
wire x_out_47_15;
wire x_out_47_18;
wire x_out_47_19;
wire x_out_47_2;
wire x_out_47_20;
wire x_out_47_21;
wire x_out_47_22;
wire x_out_47_23;
wire x_out_47_24;
wire x_out_47_25;
wire x_out_47_26;
wire x_out_47_27;
wire x_out_47_28;
wire x_out_47_29;
wire x_out_47_3;
wire x_out_47_30;
wire x_out_47_31;
wire x_out_47_32;
wire x_out_47_33;
wire x_out_47_4;
wire x_out_47_5;
wire x_out_47_6;
wire x_out_47_7;
wire x_out_47_8;
wire x_out_47_9;
wire x_out_48_0;
wire x_out_48_1;
wire x_out_48_10;
wire x_out_48_11;
wire x_out_48_12;
wire x_out_48_13;
wire x_out_48_14;
wire x_out_48_15;
wire x_out_48_18;
wire x_out_48_19;
wire x_out_48_2;
wire x_out_48_20;
wire x_out_48_21;
wire x_out_48_22;
wire x_out_48_23;
wire x_out_48_24;
wire x_out_48_25;
wire x_out_48_26;
wire x_out_48_27;
wire x_out_48_28;
wire x_out_48_29;
wire x_out_48_3;
wire x_out_48_30;
wire x_out_48_31;
wire x_out_48_32;
wire x_out_48_33;
wire x_out_48_4;
wire x_out_48_5;
wire x_out_48_6;
wire x_out_48_7;
wire x_out_48_8;
wire x_out_48_9;
wire x_out_49_0;
wire x_out_49_1;
wire x_out_49_10;
wire x_out_49_11;
wire x_out_49_12;
wire x_out_49_13;
wire x_out_49_14;
wire x_out_49_15;
wire x_out_49_18;
wire x_out_49_19;
wire x_out_49_2;
wire x_out_49_20;
wire x_out_49_21;
wire x_out_49_22;
wire x_out_49_23;
wire x_out_49_24;
wire x_out_49_25;
wire x_out_49_26;
wire x_out_49_27;
wire x_out_49_28;
wire x_out_49_29;
wire x_out_49_3;
wire x_out_49_30;
wire x_out_49_31;
wire x_out_49_32;
wire x_out_49_33;
wire x_out_49_4;
wire x_out_49_5;
wire x_out_49_6;
wire x_out_49_7;
wire x_out_49_8;
wire x_out_49_9;
wire x_out_4_0;
wire x_out_4_1;
wire x_out_4_10;
wire x_out_4_11;
wire x_out_4_12;
wire x_out_4_13;
wire x_out_4_14;
wire x_out_4_15;
wire x_out_4_18;
wire x_out_4_19;
wire x_out_4_2;
wire x_out_4_20;
wire x_out_4_21;
wire x_out_4_22;
wire x_out_4_23;
wire x_out_4_24;
wire x_out_4_25;
wire x_out_4_26;
wire x_out_4_27;
wire x_out_4_28;
wire x_out_4_29;
wire x_out_4_3;
wire x_out_4_30;
wire x_out_4_31;
wire x_out_4_32;
wire x_out_4_33;
wire x_out_4_4;
wire x_out_4_5;
wire x_out_4_6;
wire x_out_4_7;
wire x_out_4_8;
wire x_out_4_9;
wire x_out_50_0;
wire x_out_50_1;
wire x_out_50_10;
wire x_out_50_11;
wire x_out_50_12;
wire x_out_50_13;
wire x_out_50_14;
wire x_out_50_15;
wire x_out_50_18;
wire x_out_50_19;
wire x_out_50_2;
wire x_out_50_20;
wire x_out_50_21;
wire x_out_50_22;
wire x_out_50_23;
wire x_out_50_24;
wire x_out_50_25;
wire x_out_50_26;
wire x_out_50_27;
wire x_out_50_28;
wire x_out_50_29;
wire x_out_50_3;
wire x_out_50_30;
wire x_out_50_31;
wire x_out_50_32;
wire x_out_50_33;
wire x_out_50_4;
wire x_out_50_5;
wire x_out_50_6;
wire x_out_50_7;
wire x_out_50_8;
wire x_out_50_9;
wire x_out_51_0;
wire x_out_51_1;
wire x_out_51_10;
wire x_out_51_11;
wire x_out_51_12;
wire x_out_51_13;
wire x_out_51_14;
wire x_out_51_15;
wire x_out_51_18;
wire x_out_51_19;
wire x_out_51_2;
wire x_out_51_20;
wire x_out_51_21;
wire x_out_51_22;
wire x_out_51_23;
wire x_out_51_24;
wire x_out_51_25;
wire x_out_51_26;
wire x_out_51_27;
wire x_out_51_28;
wire x_out_51_29;
wire x_out_51_3;
wire x_out_51_30;
wire x_out_51_31;
wire x_out_51_32;
wire x_out_51_33;
wire x_out_51_4;
wire x_out_51_5;
wire x_out_51_6;
wire x_out_51_7;
wire x_out_51_8;
wire x_out_51_9;
wire x_out_52_0;
wire x_out_52_1;
wire x_out_52_10;
wire x_out_52_11;
wire x_out_52_12;
wire x_out_52_13;
wire x_out_52_14;
wire x_out_52_15;
wire x_out_52_2;
wire x_out_52_3;
wire x_out_52_4;
wire x_out_52_5;
wire x_out_52_6;
wire x_out_52_7;
wire x_out_52_8;
wire x_out_52_9;
wire x_out_53_0;
wire x_out_53_1;
wire x_out_53_10;
wire x_out_53_11;
wire x_out_53_12;
wire x_out_53_13;
wire x_out_53_14;
wire x_out_53_15;
wire x_out_53_18;
wire x_out_53_19;
wire x_out_53_2;
wire x_out_53_20;
wire x_out_53_21;
wire x_out_53_22;
wire x_out_53_23;
wire x_out_53_24;
wire x_out_53_25;
wire x_out_53_26;
wire x_out_53_27;
wire x_out_53_28;
wire x_out_53_29;
wire x_out_53_3;
wire x_out_53_30;
wire x_out_53_31;
wire x_out_53_32;
wire x_out_53_33;
wire x_out_53_4;
wire x_out_53_5;
wire x_out_53_6;
wire x_out_53_7;
wire x_out_53_8;
wire x_out_53_9;
wire x_out_54_0;
wire x_out_54_1;
wire x_out_54_10;
wire x_out_54_11;
wire x_out_54_12;
wire x_out_54_13;
wire x_out_54_14;
wire x_out_54_15;
wire x_out_54_18;
wire x_out_54_19;
wire x_out_54_2;
wire x_out_54_20;
wire x_out_54_21;
wire x_out_54_22;
wire x_out_54_23;
wire x_out_54_24;
wire x_out_54_25;
wire x_out_54_26;
wire x_out_54_27;
wire x_out_54_28;
wire x_out_54_29;
wire x_out_54_3;
wire x_out_54_30;
wire x_out_54_31;
wire x_out_54_32;
wire x_out_54_33;
wire x_out_54_4;
wire x_out_54_5;
wire x_out_54_6;
wire x_out_54_7;
wire x_out_54_8;
wire x_out_54_9;
wire x_out_55_0;
wire x_out_55_1;
wire x_out_55_10;
wire x_out_55_11;
wire x_out_55_12;
wire x_out_55_13;
wire x_out_55_14;
wire x_out_55_15;
wire x_out_55_18;
wire x_out_55_19;
wire x_out_55_2;
wire x_out_55_20;
wire x_out_55_21;
wire x_out_55_22;
wire x_out_55_23;
wire x_out_55_24;
wire x_out_55_25;
wire x_out_55_26;
wire x_out_55_27;
wire x_out_55_28;
wire x_out_55_29;
wire x_out_55_3;
wire x_out_55_30;
wire x_out_55_31;
wire x_out_55_32;
wire x_out_55_33;
wire x_out_55_4;
wire x_out_55_5;
wire x_out_55_6;
wire x_out_55_7;
wire x_out_55_8;
wire x_out_55_9;
wire x_out_56_0;
wire x_out_56_1;
wire x_out_56_10;
wire x_out_56_11;
wire x_out_56_12;
wire x_out_56_13;
wire x_out_56_14;
wire x_out_56_15;
wire x_out_56_18;
wire x_out_56_19;
wire x_out_56_2;
wire x_out_56_20;
wire x_out_56_21;
wire x_out_56_22;
wire x_out_56_23;
wire x_out_56_24;
wire x_out_56_25;
wire x_out_56_26;
wire x_out_56_27;
wire x_out_56_28;
wire x_out_56_29;
wire x_out_56_3;
wire x_out_56_30;
wire x_out_56_31;
wire x_out_56_32;
wire x_out_56_33;
wire x_out_56_4;
wire x_out_56_5;
wire x_out_56_6;
wire x_out_56_7;
wire x_out_56_8;
wire x_out_56_9;
wire x_out_57_0;
wire x_out_57_1;
wire x_out_57_10;
wire x_out_57_11;
wire x_out_57_12;
wire x_out_57_13;
wire x_out_57_14;
wire x_out_57_15;
wire x_out_57_18;
wire x_out_57_19;
wire x_out_57_2;
wire x_out_57_20;
wire x_out_57_21;
wire x_out_57_22;
wire x_out_57_23;
wire x_out_57_24;
wire x_out_57_25;
wire x_out_57_26;
wire x_out_57_27;
wire x_out_57_28;
wire x_out_57_29;
wire x_out_57_3;
wire x_out_57_30;
wire x_out_57_31;
wire x_out_57_32;
wire x_out_57_33;
wire x_out_57_4;
wire x_out_57_5;
wire x_out_57_6;
wire x_out_57_7;
wire x_out_57_8;
wire x_out_57_9;
wire x_out_58_0;
wire x_out_58_1;
wire x_out_58_10;
wire x_out_58_11;
wire x_out_58_12;
wire x_out_58_13;
wire x_out_58_14;
wire x_out_58_15;
wire x_out_58_18;
wire x_out_58_19;
wire x_out_58_2;
wire x_out_58_20;
wire x_out_58_21;
wire x_out_58_22;
wire x_out_58_23;
wire x_out_58_24;
wire x_out_58_25;
wire x_out_58_26;
wire x_out_58_27;
wire x_out_58_28;
wire x_out_58_29;
wire x_out_58_3;
wire x_out_58_30;
wire x_out_58_31;
wire x_out_58_32;
wire x_out_58_33;
wire x_out_58_4;
wire x_out_58_5;
wire x_out_58_6;
wire x_out_58_7;
wire x_out_58_8;
wire x_out_58_9;
wire x_out_59_0;
wire x_out_59_1;
wire x_out_59_10;
wire x_out_59_11;
wire x_out_59_12;
wire x_out_59_13;
wire x_out_59_14;
wire x_out_59_15;
wire x_out_59_18;
wire x_out_59_19;
wire x_out_59_2;
wire x_out_59_20;
wire x_out_59_21;
wire x_out_59_22;
wire x_out_59_23;
wire x_out_59_24;
wire x_out_59_25;
wire x_out_59_26;
wire x_out_59_27;
wire x_out_59_28;
wire x_out_59_29;
wire x_out_59_3;
wire x_out_59_30;
wire x_out_59_31;
wire x_out_59_32;
wire x_out_59_33;
wire x_out_59_4;
wire x_out_59_5;
wire x_out_59_6;
wire x_out_59_7;
wire x_out_59_8;
wire x_out_59_9;
wire x_out_5_0;
wire x_out_5_1;
wire x_out_5_10;
wire x_out_5_11;
wire x_out_5_12;
wire x_out_5_13;
wire x_out_5_14;
wire x_out_5_15;
wire x_out_5_18;
wire x_out_5_19;
wire x_out_5_2;
wire x_out_5_20;
wire x_out_5_21;
wire x_out_5_22;
wire x_out_5_23;
wire x_out_5_24;
wire x_out_5_25;
wire x_out_5_26;
wire x_out_5_27;
wire x_out_5_28;
wire x_out_5_29;
wire x_out_5_3;
wire x_out_5_30;
wire x_out_5_31;
wire x_out_5_32;
wire x_out_5_33;
wire x_out_5_4;
wire x_out_5_5;
wire x_out_5_6;
wire x_out_5_7;
wire x_out_5_8;
wire x_out_5_9;
wire x_out_60_0;
wire x_out_60_1;
wire x_out_60_10;
wire x_out_60_11;
wire x_out_60_12;
wire x_out_60_13;
wire x_out_60_14;
wire x_out_60_15;
wire x_out_60_18;
wire x_out_60_19;
wire x_out_60_2;
wire x_out_60_20;
wire x_out_60_21;
wire x_out_60_22;
wire x_out_60_23;
wire x_out_60_24;
wire x_out_60_25;
wire x_out_60_26;
wire x_out_60_27;
wire x_out_60_28;
wire x_out_60_29;
wire x_out_60_3;
wire x_out_60_30;
wire x_out_60_31;
wire x_out_60_32;
wire x_out_60_33;
wire x_out_60_4;
wire x_out_60_5;
wire x_out_60_6;
wire x_out_60_7;
wire x_out_60_8;
wire x_out_60_9;
wire x_out_61_0;
wire x_out_61_1;
wire x_out_61_10;
wire x_out_61_11;
wire x_out_61_12;
wire x_out_61_13;
wire x_out_61_14;
wire x_out_61_15;
wire x_out_61_18;
wire x_out_61_19;
wire x_out_61_2;
wire x_out_61_20;
wire x_out_61_21;
wire x_out_61_22;
wire x_out_61_23;
wire x_out_61_24;
wire x_out_61_25;
wire x_out_61_26;
wire x_out_61_27;
wire x_out_61_28;
wire x_out_61_29;
wire x_out_61_3;
wire x_out_61_30;
wire x_out_61_31;
wire x_out_61_32;
wire x_out_61_33;
wire x_out_61_4;
wire x_out_61_5;
wire x_out_61_6;
wire x_out_61_7;
wire x_out_61_8;
wire x_out_61_9;
wire x_out_62_0;
wire x_out_62_1;
wire x_out_62_10;
wire x_out_62_11;
wire x_out_62_12;
wire x_out_62_13;
wire x_out_62_14;
wire x_out_62_15;
wire x_out_62_18;
wire x_out_62_19;
wire x_out_62_2;
wire x_out_62_20;
wire x_out_62_21;
wire x_out_62_22;
wire x_out_62_23;
wire x_out_62_24;
wire x_out_62_25;
wire x_out_62_26;
wire x_out_62_27;
wire x_out_62_28;
wire x_out_62_29;
wire x_out_62_3;
wire x_out_62_30;
wire x_out_62_31;
wire x_out_62_32;
wire x_out_62_33;
wire x_out_62_4;
wire x_out_62_5;
wire x_out_62_6;
wire x_out_62_7;
wire x_out_62_8;
wire x_out_62_9;
wire x_out_63_0;
wire x_out_63_1;
wire x_out_63_10;
wire x_out_63_11;
wire x_out_63_12;
wire x_out_63_13;
wire x_out_63_14;
wire x_out_63_15;
wire x_out_63_18;
wire x_out_63_19;
wire x_out_63_2;
wire x_out_63_20;
wire x_out_63_21;
wire x_out_63_22;
wire x_out_63_23;
wire x_out_63_24;
wire x_out_63_25;
wire x_out_63_26;
wire x_out_63_27;
wire x_out_63_28;
wire x_out_63_29;
wire x_out_63_3;
wire x_out_63_30;
wire x_out_63_31;
wire x_out_63_32;
wire x_out_63_33;
wire x_out_63_4;
wire x_out_63_5;
wire x_out_63_6;
wire x_out_63_7;
wire x_out_63_8;
wire x_out_63_9;
wire x_out_6_0;
wire x_out_6_1;
wire x_out_6_10;
wire x_out_6_11;
wire x_out_6_12;
wire x_out_6_13;
wire x_out_6_14;
wire x_out_6_15;
wire x_out_6_18;
wire x_out_6_19;
wire x_out_6_2;
wire x_out_6_20;
wire x_out_6_21;
wire x_out_6_22;
wire x_out_6_23;
wire x_out_6_24;
wire x_out_6_25;
wire x_out_6_26;
wire x_out_6_27;
wire x_out_6_28;
wire x_out_6_29;
wire x_out_6_3;
wire x_out_6_30;
wire x_out_6_31;
wire x_out_6_32;
wire x_out_6_33;
wire x_out_6_4;
wire x_out_6_5;
wire x_out_6_6;
wire x_out_6_7;
wire x_out_6_8;
wire x_out_6_9;
wire x_out_7_0;
wire x_out_7_1;
wire x_out_7_10;
wire x_out_7_11;
wire x_out_7_12;
wire x_out_7_13;
wire x_out_7_14;
wire x_out_7_15;
wire x_out_7_18;
wire x_out_7_19;
wire x_out_7_2;
wire x_out_7_20;
wire x_out_7_21;
wire x_out_7_22;
wire x_out_7_23;
wire x_out_7_24;
wire x_out_7_25;
wire x_out_7_26;
wire x_out_7_27;
wire x_out_7_28;
wire x_out_7_29;
wire x_out_7_3;
wire x_out_7_30;
wire x_out_7_31;
wire x_out_7_32;
wire x_out_7_33;
wire x_out_7_4;
wire x_out_7_5;
wire x_out_7_6;
wire x_out_7_7;
wire x_out_7_8;
wire x_out_7_9;
wire x_out_8_0;
wire x_out_8_1;
wire x_out_8_10;
wire x_out_8_11;
wire x_out_8_12;
wire x_out_8_13;
wire x_out_8_14;
wire x_out_8_15;
wire x_out_8_18;
wire x_out_8_19;
wire x_out_8_2;
wire x_out_8_20;
wire x_out_8_21;
wire x_out_8_22;
wire x_out_8_23;
wire x_out_8_24;
wire x_out_8_25;
wire x_out_8_26;
wire x_out_8_27;
wire x_out_8_28;
wire x_out_8_29;
wire x_out_8_3;
wire x_out_8_30;
wire x_out_8_31;
wire x_out_8_32;
wire x_out_8_33;
wire x_out_8_4;
wire x_out_8_5;
wire x_out_8_6;
wire x_out_8_7;
wire x_out_8_8;
wire x_out_8_9;
wire x_out_9_0;
wire x_out_9_1;
wire x_out_9_10;
wire x_out_9_11;
wire x_out_9_12;
wire x_out_9_13;
wire x_out_9_14;
wire x_out_9_15;
wire x_out_9_18;
wire x_out_9_19;
wire x_out_9_2;
wire x_out_9_20;
wire x_out_9_21;
wire x_out_9_22;
wire x_out_9_23;
wire x_out_9_24;
wire x_out_9_25;
wire x_out_9_26;
wire x_out_9_27;
wire x_out_9_28;
wire x_out_9_29;
wire x_out_9_3;
wire x_out_9_30;
wire x_out_9_31;
wire x_out_9_32;
wire x_out_9_33;
wire x_out_9_4;
wire x_out_9_5;
wire x_out_9_6;
wire x_out_9_7;
wire x_out_9_8;
wire x_out_9_9;

// Start cells
in01f80 FE_OFC0_n_17395 ( .a(n_17395), .o(FE_OFN0_n_17395) );
in01f80 FE_OFC1000_n_17200 ( .a(n_17200), .o(FE_OFN1000_n_17200) );
in01f80 FE_OFC1001_n_17200 ( .a(FE_OFN1000_n_17200), .o(FE_OFN1001_n_17200) );
in01f80 FE_OFC1002_n_19855 ( .a(n_19855), .o(FE_OFN1002_n_19855) );
in01f80 FE_OFC1003_n_19855 ( .a(FE_OFN1002_n_19855), .o(FE_OFN1003_n_19855) );
in01f80 FE_OFC1004_n_23624 ( .a(n_23624), .o(FE_OFN1004_n_23624) );
in01f80 FE_OFC1005_n_23624 ( .a(FE_OFN1004_n_23624), .o(FE_OFN1005_n_23624) );
in01f80 FE_OFC1006_n_24950 ( .a(n_24950), .o(FE_OFN1006_n_24950) );
in01f80 FE_OFC1007_n_24950 ( .a(FE_OFN1006_n_24950), .o(FE_OFN1007_n_24950) );
in01f80 FE_OFC1008_n_27881 ( .a(n_27881), .o(FE_OFN1008_n_27881) );
in01f80 FE_OFC1009_n_27881 ( .a(FE_OFN1008_n_27881), .o(FE_OFN1009_n_27881) );
in01f80 FE_OFC100_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN100_n_27449) );
in01f80 FE_OFC1010_n_28328 ( .a(n_28328), .o(FE_OFN1010_n_28328) );
in01f80 FE_OFC1011_n_28328 ( .a(FE_OFN1010_n_28328), .o(FE_OFN1011_n_28328) );
in01f80 FE_OFC1012_n_28629 ( .a(n_28629), .o(FE_OFN1012_n_28629) );
in01f80 FE_OFC1014_n_16571 ( .a(n_16571), .o(FE_OFN1014_n_16571) );
in01f80 FE_OFC1015_n_16571 ( .a(FE_OFN1014_n_16571), .o(FE_OFN1015_n_16571) );
in01f80 FE_OFC1016_n_17433 ( .a(n_17433), .o(FE_OFN1016_n_17433) );
in01f80 FE_OFC1017_n_17433 ( .a(FE_OFN1016_n_17433), .o(FE_OFN1017_n_17433) );
in01f80 FE_OFC1018_n_22081 ( .a(n_22081), .o(FE_OFN1018_n_22081) );
in01f80 FE_OFC1019_n_22081 ( .a(FE_OFN1018_n_22081), .o(FE_OFN1019_n_22081) );
in01f80 FE_OFC101_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN101_n_27449) );
in01f80 FE_OFC1020_n_28703 ( .a(n_28703), .o(FE_OFN1020_n_28703) );
in01f80 FE_OFC1021_n_28703 ( .a(FE_OFN1020_n_28703), .o(FE_OFN1021_n_28703) );
in01f80 FE_OFC1028_n_14570 ( .a(n_14570), .o(FE_OFN1028_n_14570) );
in01f80 FE_OFC1029_n_14570 ( .a(FE_OFN1028_n_14570), .o(FE_OFN1029_n_14570) );
in01f80 FE_OFC102_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN102_n_27449) );
in01f80 FE_OFC1030_n_19666 ( .a(n_19666), .o(FE_OFN1030_n_19666) );
in01f80 FE_OFC1031_n_19666 ( .a(FE_OFN1030_n_19666), .o(FE_OFN1031_n_19666) );
in01f80 FE_OFC1034_n_21194 ( .a(n_21194), .o(FE_OFN1034_n_21194) );
in01f80 FE_OFC1035_n_21194 ( .a(FE_OFN1034_n_21194), .o(FE_OFN1035_n_21194) );
in01f80 FE_OFC1036_n_26168 ( .a(n_26168), .o(FE_OFN1036_n_26168) );
in01f80 FE_OFC1037_n_26168 ( .a(FE_OFN1036_n_26168), .o(FE_OFN1037_n_26168) );
in01f80 FE_OFC1038_n_27890 ( .a(n_27890), .o(FE_OFN1038_n_27890) );
in01f80 FE_OFC1039_n_27890 ( .a(FE_OFN1038_n_27890), .o(FE_OFN1039_n_27890) );
in01f80 FE_OFC103_n_27449 ( .a(FE_OFN90_n_27449), .o(FE_OFN103_n_27449) );
in01f80 FE_OFC1044_n_26162 ( .a(n_26162), .o(FE_OFN1044_n_26162) );
in01f80 FE_OFC1045_n_26162 ( .a(FE_OFN1044_n_26162), .o(FE_OFN1045_n_26162) );
in01f80 FE_OFC1046_n_27057 ( .a(n_27057), .o(FE_OFN1046_n_27057) );
in01f80 FE_OFC1047_n_27057 ( .a(FE_OFN1046_n_27057), .o(FE_OFN1047_n_27057) );
in01f80 FE_OFC104_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN104_n_27449) );
in01f80 FE_OFC1054_n_25805 ( .a(n_25805), .o(FE_OFN1054_n_25805) );
in01f80 FE_OFC1055_n_25805 ( .a(FE_OFN1054_n_25805), .o(FE_OFN1055_n_25805) );
in01f80 FE_OFC1056_n_18817 ( .a(n_18817), .o(FE_OFN1056_n_18817) );
in01f80 FE_OFC1057_n_18817 ( .a(FE_OFN1056_n_18817), .o(FE_OFN1057_n_18817) );
in01f80 FE_OFC1058_n_18610 ( .a(n_18610), .o(FE_OFN1058_n_18610) );
in01f80 FE_OFC1059_n_18610 ( .a(FE_OFN1058_n_18610), .o(FE_OFN1059_n_18610) );
in01f80 FE_OFC105_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN105_n_27449) );
in01f80 FE_OFC1060_n_19587 ( .a(n_19587), .o(FE_OFN1060_n_19587) );
in01f80 FE_OFC1061_n_19587 ( .a(FE_OFN1060_n_19587), .o(FE_OFN1061_n_19587) );
in01f80 FE_OFC106_n_27449 ( .a(FE_OFN91_n_27449), .o(FE_OFN106_n_27449) );
in01f80 FE_OFC1073_n_6399 ( .a(FE_OFN1129_n_6399), .o(FE_OFN1073_n_6399) );
in01f80 FE_OFC107_n_27449 ( .a(FE_OFN90_n_27449), .o(FE_OFN107_n_27449) );
in01f80 FE_OFC1080_n_14273 ( .a(n_14273), .o(FE_OFN1080_n_14273) );
in01f80 FE_OFC1081_n_14273 ( .a(FE_OFN1080_n_14273), .o(FE_OFN1081_n_14273) );
in01f80 FE_OFC1082_n_8877 ( .a(n_8877), .o(FE_OFN1082_n_8877) );
in01f80 FE_OFC1083_n_8877 ( .a(FE_OFN1082_n_8877), .o(FE_OFN1083_n_8877) );
in01f80 FE_OFC1084_n_14427 ( .a(n_14427), .o(FE_OFN1084_n_14427) );
in01f80 FE_OFC1085_n_14427 ( .a(FE_OFN1084_n_14427), .o(FE_OFN1085_n_14427) );
in01f80 FE_OFC1086_n_8974 ( .a(n_8974), .o(FE_OFN1086_n_8974) );
in01f80 FE_OFC1087_n_8974 ( .a(FE_OFN1086_n_8974), .o(FE_OFN1087_n_8974) );
in01f80 FE_OFC1088_n_8985 ( .a(n_8985), .o(FE_OFN1088_n_8985) );
in01f80 FE_OFC1089_n_8985 ( .a(FE_OFN1088_n_8985), .o(FE_OFN1089_n_8985) );
in01f80 FE_OFC108_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN108_n_27449) );
in01f80 FE_OFC1090_n_8621 ( .a(n_8621), .o(FE_OFN1090_n_8621) );
in01f80 FE_OFC1091_n_8621 ( .a(FE_OFN1090_n_8621), .o(FE_OFN1091_n_8621) );
in01f80 FE_OFC109_n_27449 ( .a(FE_OFN93_n_27449), .o(FE_OFN109_n_27449) );
in01f80 FE_OFC10_n_29204 ( .a(n_29204), .o(FE_OFN10_n_29204) );
in01f80 FE_OFC1100_n_12369 ( .a(n_12369), .o(FE_OFN1100_n_12369) );
in01f80 FE_OFC1101_n_12369 ( .a(FE_OFN1100_n_12369), .o(FE_OFN1101_n_12369) );
in01f80 FE_OFC1102_rst ( .a(rst), .o(FE_OFN1102_rst) );
in01f80 FE_OFC1103_rst ( .a(rst), .o(FE_OFN1103_rst) );
in01f80 FE_OFC1104_rst ( .a(rst), .o(FE_OFN1104_rst) );
in01f80 FE_OFC1105_rst ( .a(rst), .o(FE_OFN1105_rst) );
in01f80 FE_OFC1106_rst ( .a(FE_OFN1104_rst), .o(FE_OFN1106_rst) );
in01f80 FE_OFC1107_rst ( .a(FE_OFN1102_rst), .o(FE_OFN1107_rst) );
in01f80 FE_OFC1108_rst ( .a(FE_OFN1102_rst), .o(FE_OFN1108_rst) );
in01f80 FE_OFC1109_rst ( .a(FE_OFN1103_rst), .o(FE_OFN1109_rst) );
in01f80 FE_OFC1110_rst ( .a(FE_OFN1104_rst), .o(FE_OFN1110_rst) );
in01f80 FE_OFC1111_rst ( .a(FE_OFN1104_rst), .o(FE_OFN1111_rst) );
in01f80 FE_OFC1112_rst ( .a(FE_OFN1105_rst), .o(FE_OFN1112_rst) );
in01f80 FE_OFC1113_rst ( .a(FE_OFN1102_rst), .o(FE_OFN1113_rst) );
in01f80 FE_OFC1114_rst ( .a(FE_OFN1102_rst), .o(FE_OFN1114_rst) );
in01f80 FE_OFC1115_rst ( .a(FE_OFN1103_rst), .o(FE_OFN1115_rst) );
in01f80 FE_OFC1117_rst ( .a(FE_OFN1103_rst), .o(FE_OFN1117_rst) );
in01f80 FE_OFC1118_rst ( .a(FE_OFN1103_rst), .o(FE_OFN1118_rst) );
in01f80 FE_OFC1119_rst ( .a(FE_OFN1103_rst), .o(FE_OFN1119_rst) );
in01f80 FE_OFC111_n_27449 ( .a(FE_OFN94_n_27449), .o(FE_OFN111_n_27449) );
in01f80 FE_OFC1120_rst ( .a(FE_OFN1105_rst), .o(FE_OFN1120_rst) );
in01f80 FE_OFC1121_rst ( .a(FE_OFN1103_rst), .o(FE_OFN1121_rst) );
in01f80 FE_OFC1122_rst ( .a(FE_OFN1108_rst), .o(FE_OFN1122_rst) );
in01f80 FE_OFC1123_rst ( .a(FE_OFN1122_rst), .o(FE_OFN1123_rst) );
in01f80 FE_OFC1124_rst ( .a(FE_OFN1122_rst), .o(FE_OFN1124_rst) );
in01f80 FE_OFC1125_n_29632 ( .a(n_29632), .o(FE_OFN1125_n_29632) );
in01f80 FE_OFC1126_n_29632 ( .a(FE_OFN1125_n_29632), .o(FE_OFN1126_n_29632) );
in01f80 FE_OFC1127_n_29567 ( .a(n_29567), .o(FE_OFN1127_n_29567) );
in01f80 FE_OFC1128_n_29567 ( .a(FE_OFN1127_n_29567), .o(FE_OFN1128_n_29567) );
in01f80 FE_OFC1129_n_6399 ( .a(n_6399), .o(FE_OFN1129_n_6399) );
in01f80 FE_OFC1130_n_27986 ( .a(n_27986), .o(FE_OFN1130_n_27986) );
in01f80 FE_OFC1131_n_28629 ( .a(FE_OFN1012_n_28629), .o(FE_OFN1131_n_28629) );
in01f80 FE_OFC1132_n_28627 ( .a(FE_OFN1134_n_28627), .o(FE_OFN1132_n_28627) );
in01f80 FE_OFC1133_n_28782 ( .a(FE_OFN998_n_28782), .o(FE_OFN1133_n_28782) );
in01f80 FE_OFC1134_n_28627 ( .a(n_28627), .o(FE_OFN1134_n_28627) );
in01f80 FE_OFC1135_n_28794 ( .a(n_28794), .o(FE_OFN1135_n_28794) );
in01f80 FE_OFC1136_n_28794 ( .a(FE_OFN1135_n_28794), .o(FE_OFN1136_n_28794) );
in01f80 FE_OFC1137_n_28938 ( .a(n_28938), .o(FE_OFN1137_n_28938) );
in01f80 FE_OFC1138_n_28938 ( .a(FE_OFN1137_n_28938), .o(FE_OFN1138_n_28938) );
in01f80 FE_OFC1139_n_27012 ( .a(FE_OFN74_n_27012), .o(FE_OFN1139_n_27012) );
in01f80 FE_OFC113_n_27449 ( .a(FE_OFN106_n_27449), .o(FE_OFN113_n_27449) );
in01f80 FE_OFC1140_n_27012 ( .a(FE_OFN1139_n_27012), .o(FE_OFN1140_n_27012) );
in01f80 FE_OFC1141_n_27012 ( .a(FE_OFN1139_n_27012), .o(FE_OFN1141_n_27012) );
in01f80 FE_OFC1142_n_27012 ( .a(n_27012), .o(FE_OFN1142_n_27012) );
in01f80 FE_OFC1143_n_27012 ( .a(FE_OFN1142_n_27012), .o(FE_OFN1143_n_27012) );
in01f80 FE_OFC1144_n_27012 ( .a(FE_OFN1142_n_27012), .o(FE_OFN1144_n_27012) );
in01f80 FE_OFC1145_n_4860 ( .a(FE_OFN364_n_4860), .o(FE_OFN1145_n_4860) );
in01f80 FE_OFC1146_n_4860 ( .a(FE_OFN1145_n_4860), .o(FE_OFN1146_n_4860) );
in01f80 FE_OFC1147_n_4860 ( .a(FE_OFN1145_n_4860), .o(FE_OFN1147_n_4860) );
in01f80 FE_OFC1148_n_6525 ( .a(n_6525), .o(FE_OFN1148_n_6525) );
in01f80 FE_OFC1149_n_6525 ( .a(FE_OFN1148_n_6525), .o(FE_OFN1149_n_6525) );
in01f80 FE_OFC114_n_27449 ( .a(FE_OFN103_n_27449), .o(FE_OFN114_n_27449) );
in01f80 FE_OFC1150_n_3069 ( .a(FE_OFN309_n_3069), .o(FE_OFN1150_n_3069) );
in01f80 FE_OFC1151_n_3069 ( .a(FE_OFN1150_n_3069), .o(FE_OFN1151_n_3069) );
in01f80 FE_OFC1152_n_3069 ( .a(FE_OFN1150_n_3069), .o(FE_OFN1152_n_3069) );
in01f80 FE_OFC1153_n_14586 ( .a(FE_OFN86_n_14586), .o(FE_OFN1153_n_14586) );
in01f80 FE_OFC1154_n_14586 ( .a(FE_OFN1153_n_14586), .o(FE_OFN1154_n_14586) );
in01f80 FE_OFC1155_n_14586 ( .a(FE_OFN1153_n_14586), .o(FE_OFN1155_n_14586) );
in01f80 FE_OFC1156_n_26184 ( .a(FE_OFN175_n_26184), .o(FE_OFN1156_n_26184) );
in01f80 FE_OFC1157_n_26184 ( .a(FE_OFN1156_n_26184), .o(FE_OFN1157_n_26184) );
in01f80 FE_OFC1158_n_26184 ( .a(n_26184), .o(FE_OFN1158_n_26184) );
in01f80 FE_OFC1159_n_26184 ( .a(FE_OFN1158_n_26184), .o(FE_OFN1159_n_26184) );
in01f80 FE_OFC115_n_27449 ( .a(FE_OFN107_n_27449), .o(FE_OFN115_n_27449) );
in01f80 FE_OFC1160_n_26184 ( .a(FE_OFN1158_n_26184), .o(FE_OFN1160_n_26184) );
in01f80 FE_OFC1161_n_5003 ( .a(n_5003), .o(FE_OFN1161_n_5003) );
in01f80 FE_OFC1162_n_5003 ( .a(FE_OFN1161_n_5003), .o(FE_OFN1162_n_5003) );
in01f80 FE_OFC1163_n_4162 ( .a(n_4162), .o(FE_OFN1163_n_4162) );
in01f80 FE_OFC1164_n_4162 ( .a(n_4162), .o(FE_OFN1164_n_4162) );
in01f80 FE_OFC1165_n_4162 ( .a(FE_OFN1163_n_4162), .o(FE_OFN1165_n_4162) );
in01f80 FE_OFC1166_n_4162 ( .a(FE_OFN1163_n_4162), .o(FE_OFN1166_n_4162) );
in01f80 FE_OFC1167_n_4162 ( .a(FE_OFN1164_n_4162), .o(FE_OFN1167_n_4162) );
in01f80 FE_OFC1168_n_4162 ( .a(FE_OFN1164_n_4162), .o(FE_OFN1168_n_4162) );
in01f80 FE_OFC1169_n_4860 ( .a(n_4860), .o(FE_OFN1169_n_4860) );
in01f80 FE_OFC116_n_27449 ( .a(FE_OFN107_n_27449), .o(FE_OFN116_n_27449) );
in01f80 FE_OFC1170_n_4860 ( .a(n_4860), .o(FE_OFN1170_n_4860) );
in01f80 FE_OFC1171_n_4860 ( .a(FE_OFN1169_n_4860), .o(FE_OFN1171_n_4860) );
in01f80 FE_OFC1172_n_4860 ( .a(FE_OFN1170_n_4860), .o(FE_OFN1172_n_4860) );
in01f80 FE_OFC1173_n_4860 ( .a(FE_OFN1170_n_4860), .o(FE_OFN1173_n_4860) );
in01f80 FE_OFC1174_n_4860 ( .a(FE_OFN1169_n_4860), .o(FE_OFN1174_n_4860) );
in01f80 FE_OFC1175_n_28597 ( .a(n_28597), .o(FE_OFN1175_n_28597) );
in01f80 FE_OFC1176_n_28597 ( .a(FE_OFN1175_n_28597), .o(FE_OFN1176_n_28597) );
in01f80 FE_OFC1177_n_28597 ( .a(FE_OFN1175_n_28597), .o(FE_OFN1177_n_28597) );
in01f80 FE_OFC1178_n_17184 ( .a(n_17184), .o(FE_OFN1178_n_17184) );
in01f80 FE_OFC1179_n_17184 ( .a(FE_OFN1178_n_17184), .o(FE_OFN1179_n_17184) );
in01f80 FE_OFC117_n_27449 ( .a(FE_OFN104_n_27449), .o(FE_OFN117_n_27449) );
in01f80 FE_OFC1180_rst ( .a(FE_OFN1107_rst), .o(FE_OFN1180_rst) );
in01f80 FE_OFC1181_rst ( .a(FE_OFN1180_rst), .o(FE_OFN1181_rst) );
in01f80 FE_OFC1182_rst ( .a(FE_OFN1180_rst), .o(FE_OFN1182_rst) );
in01f80 FE_OFC1183_n_6701 ( .a(n_6701), .o(FE_OFN1183_n_6701) );
in01f80 FE_OFC1184_n_6701 ( .a(FE_OFN1183_n_6701), .o(FE_OFN1184_n_6701) );
in01f80 FE_OFC1185_n_12201 ( .a(n_12201), .o(FE_OFN1185_n_12201) );
in01f80 FE_OFC1186_n_12201 ( .a(FE_OFN1185_n_12201), .o(FE_OFN1186_n_12201) );
in01f80 FE_OFC1187_n_5249 ( .a(n_5249), .o(FE_OFN1187_n_5249) );
in01f80 FE_OFC1188_n_5249 ( .a(FE_OFN1187_n_5249), .o(FE_OFN1188_n_5249) );
in01f80 FE_OFC1189_n_13090 ( .a(n_13090), .o(FE_OFN1189_n_13090) );
in01f80 FE_OFC118_n_27449 ( .a(FE_OFN108_n_27449), .o(FE_OFN118_n_27449) );
in01f80 FE_OFC1190_n_13090 ( .a(FE_OFN1189_n_13090), .o(FE_OFN1190_n_13090) );
in01f80 FE_OFC1191_n_11896 ( .a(n_11896), .o(FE_OFN1191_n_11896) );
in01f80 FE_OFC1192_n_11896 ( .a(FE_OFN1191_n_11896), .o(FE_OFN1192_n_11896) );
in01f80 FE_OFC1193_n_12908 ( .a(n_12908), .o(FE_OFN1193_n_12908) );
in01f80 FE_OFC1194_n_12908 ( .a(FE_OFN1193_n_12908), .o(FE_OFN1194_n_12908) );
in01f80 FE_OFC1195_n_12016 ( .a(n_12016), .o(FE_OFN1195_n_12016) );
in01f80 FE_OFC1196_n_12016 ( .a(FE_OFN1195_n_12016), .o(FE_OFN1196_n_12016) );
in01f80 FE_OFC1197_n_13003 ( .a(n_13003), .o(FE_OFN1197_n_13003) );
in01f80 FE_OFC1198_n_13003 ( .a(FE_OFN1197_n_13003), .o(FE_OFN1198_n_13003) );
in01f80 FE_OFC1199_n_10340 ( .a(n_10340), .o(FE_OFN1199_n_10340) );
in01f80 FE_OFC119_n_27449 ( .a(FE_OFN109_n_27449), .o(FE_OFN119_n_27449) );
in01f80 FE_OFC11_n_29204 ( .a(FE_OFN10_n_29204), .o(FE_OFN11_n_29204) );
in01f80 FE_OFC1200_n_10340 ( .a(FE_OFN1199_n_10340), .o(FE_OFN1200_n_10340) );
in01f80 FE_OFC1201_n_5312 ( .a(n_5312), .o(FE_OFN1201_n_5312) );
in01f80 FE_OFC1202_n_5312 ( .a(FE_OFN1201_n_5312), .o(FE_OFN1202_n_5312) );
in01f80 FE_OFC1203_n_11679 ( .a(n_11679), .o(FE_OFN1203_n_11679) );
in01f80 FE_OFC1204_n_11679 ( .a(FE_OFN1203_n_11679), .o(FE_OFN1204_n_11679) );
in01f80 FE_OFC1205_n_9308 ( .a(n_9308), .o(FE_OFN1205_n_9308) );
in01f80 FE_OFC1206_n_9308 ( .a(FE_OFN1205_n_9308), .o(FE_OFN1206_n_9308) );
in01f80 FE_OFC1207_n_10456 ( .a(n_10456), .o(FE_OFN1207_n_10456) );
in01f80 FE_OFC1208_n_10456 ( .a(FE_OFN1207_n_10456), .o(FE_OFN1208_n_10456) );
in01f80 FE_OFC1209_n_10458 ( .a(n_10458), .o(FE_OFN1209_n_10458) );
in01f80 FE_OFC120_n_27449 ( .a(FE_OFN100_n_27449), .o(FE_OFN120_n_27449) );
in01f80 FE_OFC1210_n_10458 ( .a(FE_OFN1209_n_10458), .o(FE_OFN1210_n_10458) );
in01f80 FE_OFC1211_n_10465 ( .a(n_10465), .o(FE_OFN1211_n_10465) );
in01f80 FE_OFC1212_n_10465 ( .a(FE_OFN1211_n_10465), .o(FE_OFN1212_n_10465) );
in01f80 FE_OFC1213_n_10469 ( .a(n_10469), .o(FE_OFN1213_n_10469) );
in01f80 FE_OFC1214_n_10469 ( .a(FE_OFN1213_n_10469), .o(FE_OFN1214_n_10469) );
in01f80 FE_OFC1215_n_12761 ( .a(n_12761), .o(FE_OFN1215_n_12761) );
in01f80 FE_OFC1216_n_12761 ( .a(FE_OFN1215_n_12761), .o(FE_OFN1216_n_12761) );
in01f80 FE_OFC1217_n_13369 ( .a(n_13369), .o(FE_OFN1217_n_13369) );
in01f80 FE_OFC1218_n_13369 ( .a(FE_OFN1217_n_13369), .o(FE_OFN1218_n_13369) );
in01f80 FE_OFC1219_n_8798 ( .a(n_8798), .o(FE_OFN1219_n_8798) );
in01f80 FE_OFC121_n_27449 ( .a(FE_OFN122_n_27449), .o(FE_OFN121_n_27449) );
in01f80 FE_OFC1220_n_8798 ( .a(FE_OFN1219_n_8798), .o(FE_OFN1220_n_8798) );
in01f80 FE_OFC1221_n_6089 ( .a(n_6089), .o(FE_OFN1221_n_6089) );
in01f80 FE_OFC1222_n_6089 ( .a(FE_OFN1221_n_6089), .o(FE_OFN1222_n_6089) );
in01f80 FE_OFC1223_n_29433 ( .a(n_29433), .o(FE_OFN1223_n_29433) );
in01f80 FE_OFC1224_n_29433 ( .a(FE_OFN1223_n_29433), .o(FE_OFN1224_n_29433) );
in01f80 FE_OFC1225_n_10183 ( .a(n_10183), .o(FE_OFN1225_n_10183) );
in01f80 FE_OFC1226_n_10183 ( .a(FE_OFN1225_n_10183), .o(FE_OFN1226_n_10183) );
in01f80 FE_OFC1227_n_23261 ( .a(n_23261), .o(FE_OFN1227_n_23261) );
in01f80 FE_OFC1228_n_23261 ( .a(FE_OFN1227_n_23261), .o(FE_OFN1228_n_23261) );
in01f80 FE_OFC1229_n_24166 ( .a(n_24166), .o(FE_OFN1229_n_24166) );
in01f80 FE_OFC122_n_27449 ( .a(FE_OFN103_n_27449), .o(FE_OFN122_n_27449) );
in01f80 FE_OFC1230_n_24166 ( .a(FE_OFN1229_n_24166), .o(FE_OFN1230_n_24166) );
in01f80 FE_OFC1231_n_12068 ( .a(n_12068), .o(FE_OFN1231_n_12068) );
in01f80 FE_OFC1232_n_12068 ( .a(FE_OFN1231_n_12068), .o(FE_OFN1232_n_12068) );
in01f80 FE_OFC1233_n_4979 ( .a(n_4979), .o(FE_OFN1233_n_4979) );
in01f80 FE_OFC1234_n_4979 ( .a(FE_OFN1233_n_4979), .o(FE_OFN1234_n_4979) );
in01f80 FE_OFC1235_n_16615 ( .a(n_16615), .o(FE_OFN1235_n_16615) );
in01f80 FE_OFC1236_n_16615 ( .a(FE_OFN1235_n_16615), .o(FE_OFN1236_n_16615) );
in01f80 FE_OFC1237_n_10491 ( .a(n_10491), .o(FE_OFN1237_n_10491) );
in01f80 FE_OFC1238_n_10491 ( .a(FE_OFN1237_n_10491), .o(FE_OFN1238_n_10491) );
in01f80 FE_OFC1239_n_10499 ( .a(n_10499), .o(FE_OFN1239_n_10499) );
in01f80 FE_OFC123_n_27449 ( .a(FE_OFN104_n_27449), .o(FE_OFN123_n_27449) );
in01f80 FE_OFC1240_n_10499 ( .a(FE_OFN1239_n_10499), .o(FE_OFN1240_n_10499) );
in01f80 FE_OFC1241_n_29553 ( .a(n_29553), .o(FE_OFN1241_n_29553) );
in01f80 FE_OFC1242_n_29553 ( .a(FE_OFN1241_n_29553), .o(FE_OFN1242_n_29553) );
in01f80 FE_OFC1243_n_12940 ( .a(n_12940), .o(FE_OFN1243_n_12940) );
in01f80 FE_OFC1244_n_12940 ( .a(FE_OFN1243_n_12940), .o(FE_OFN1244_n_12940) );
in01f80 FE_OFC1245_n_4900 ( .a(n_4900), .o(FE_OFN1245_n_4900) );
in01f80 FE_OFC1246_n_4900 ( .a(FE_OFN1245_n_4900), .o(FE_OFN1246_n_4900) );
in01f80 FE_OFC1247_n_8470 ( .a(n_8470), .o(FE_OFN1247_n_8470) );
in01f80 FE_OFC1248_n_8470 ( .a(FE_OFN1247_n_8470), .o(FE_OFN1248_n_8470) );
in01f80 FE_OFC1249_n_5334 ( .a(n_5334), .o(FE_OFN1249_n_5334) );
in01f80 FE_OFC124_n_27449 ( .a(FE_OFN109_n_27449), .o(FE_OFN124_n_27449) );
in01f80 FE_OFC1250_n_5334 ( .a(FE_OFN1249_n_5334), .o(FE_OFN1250_n_5334) );
in01f80 FE_OFC1251_n_25296 ( .a(n_25296), .o(FE_OFN1251_n_25296) );
in01f80 FE_OFC1252_n_25296 ( .a(FE_OFN1251_n_25296), .o(FE_OFN1252_n_25296) );
in01f80 FE_OFC1253_n_12186 ( .a(n_12186), .o(FE_OFN1253_n_12186) );
in01f80 FE_OFC1254_n_12186 ( .a(FE_OFN1253_n_12186), .o(FE_OFN1254_n_12186) );
in01f80 FE_OFC1255_n_10520 ( .a(n_10520), .o(FE_OFN1255_n_10520) );
in01f80 FE_OFC1256_n_10520 ( .a(FE_OFN1255_n_10520), .o(FE_OFN1256_n_10520) );
in01f80 FE_OFC1257_n_4905 ( .a(n_4905), .o(FE_OFN1257_n_4905) );
in01f80 FE_OFC1258_n_4905 ( .a(FE_OFN1257_n_4905), .o(FE_OFN1258_n_4905) );
in01f80 FE_OFC1259_n_6178 ( .a(n_6178), .o(FE_OFN1259_n_6178) );
in01f80 FE_OFC125_n_27449 ( .a(FE_OFN109_n_27449), .o(FE_OFN125_n_27449) );
in01f80 FE_OFC1260_n_6178 ( .a(FE_OFN1259_n_6178), .o(FE_OFN1260_n_6178) );
in01f80 FE_OFC1261_n_6197 ( .a(n_6197), .o(FE_OFN1261_n_6197) );
in01f80 FE_OFC1262_n_6197 ( .a(FE_OFN1261_n_6197), .o(FE_OFN1262_n_6197) );
in01f80 FE_OFC1263_n_29354 ( .a(n_29354), .o(FE_OFN1263_n_29354) );
in01f80 FE_OFC1264_n_29354 ( .a(FE_OFN1263_n_29354), .o(FE_OFN1264_n_29354) );
in01f80 FE_OFC1265_n_16620 ( .a(n_16620), .o(FE_OFN1265_n_16620) );
in01f80 FE_OFC1266_n_16620 ( .a(FE_OFN1265_n_16620), .o(FE_OFN1266_n_16620) );
in01f80 FE_OFC1267_n_29314 ( .a(n_29314), .o(FE_OFN1267_n_29314) );
in01f80 FE_OFC1268_n_29314 ( .a(FE_OFN1267_n_29314), .o(FE_OFN1268_n_29314) );
in01f80 FE_OFC1269_n_29015 ( .a(n_29015), .o(FE_OFN1269_n_29015) );
in01f80 FE_OFC126_n_27449 ( .a(FE_OFN111_n_27449), .o(FE_OFN126_n_27449) );
in01f80 FE_OFC1270_n_29015 ( .a(FE_OFN1269_n_29015), .o(FE_OFN1270_n_29015) );
in01f80 FE_OFC1271_n_9600 ( .a(n_9600), .o(FE_OFN1271_n_9600) );
in01f80 FE_OFC1272_n_9600 ( .a(FE_OFN1271_n_9600), .o(FE_OFN1272_n_9600) );
in01f80 FE_OFC1273_n_8977 ( .a(n_8977), .o(FE_OFN1273_n_8977) );
in01f80 FE_OFC1274_n_8977 ( .a(FE_OFN1273_n_8977), .o(FE_OFN1274_n_8977) );
in01f80 FE_OFC1275_n_12754 ( .a(n_12754), .o(FE_OFN1275_n_12754) );
in01f80 FE_OFC1276_n_12754 ( .a(FE_OFN1275_n_12754), .o(FE_OFN1276_n_12754) );
in01f80 FE_OFC1277_n_6116 ( .a(n_6116), .o(FE_OFN1277_n_6116) );
in01f80 FE_OFC1278_n_6116 ( .a(FE_OFN1277_n_6116), .o(FE_OFN1278_n_6116) );
in01f80 FE_OFC1279_n_8068 ( .a(n_8068), .o(FE_OFN1279_n_8068) );
in01f80 FE_OFC127_n_27449 ( .a(FE_OFN111_n_27449), .o(FE_OFN127_n_27449) );
in01f80 FE_OFC1280_n_8068 ( .a(FE_OFN1279_n_8068), .o(FE_OFN1280_n_8068) );
in01f80 FE_OFC128_n_27449 ( .a(FE_OFN103_n_27449), .o(FE_OFN128_n_27449) );
in01f80 FE_OFC129_n_27449 ( .a(FE_OFN103_n_27449), .o(FE_OFN129_n_27449) );
in01f80 FE_OFC12_n_29204 ( .a(FE_OFN10_n_29204), .o(FE_OFN12_n_29204) );
in01f80 FE_OFC130_n_27449 ( .a(FE_OFN117_n_27449), .o(FE_OFN130_n_27449) );
in01f80 FE_OFC131_n_27449 ( .a(FE_OFN118_n_27449), .o(FE_OFN131_n_27449) );
in01f80 FE_OFC133_n_27449 ( .a(FE_OFN120_n_27449), .o(FE_OFN133_n_27449) );
in01f80 FE_OFC134_n_27449 ( .a(FE_OFN121_n_27449), .o(FE_OFN134_n_27449) );
in01f80 FE_OFC135_n_27449 ( .a(FE_OFN117_n_27449), .o(FE_OFN135_n_27449) );
in01f80 FE_OFC136_n_27449 ( .a(FE_OFN117_n_27449), .o(FE_OFN136_n_27449) );
in01f80 FE_OFC138_n_27449 ( .a(FE_OFN123_n_27449), .o(FE_OFN138_n_27449) );
in01f80 FE_OFC139_n_27449 ( .a(FE_OFN118_n_27449), .o(FE_OFN139_n_27449) );
in01f80 FE_OFC13_n_29068 ( .a(n_29068), .o(FE_OFN13_n_29068) );
in01f80 FE_OFC141_n_27449 ( .a(FE_OFN123_n_27449), .o(FE_OFN141_n_27449) );
in01f80 FE_OFC142_n_27449 ( .a(FE_OFN123_n_27449), .o(FE_OFN142_n_27449) );
in01f80 FE_OFC143_n_7361 ( .a(n_7361), .o(FE_OFN143_n_7361) );
in01f80 FE_OFC144_n_7361 ( .a(FE_OFN143_n_7361), .o(FE_OFN144_n_7361) );
in01f80 FE_OFC145_n_2667 ( .a(n_27012), .o(FE_OFN145_n_2667) );
in01f80 FE_OFC146_n_2667 ( .a(FE_OFN145_n_2667), .o(FE_OFN146_n_2667) );
in01f80 FE_OFC147_n_25677 ( .a(n_16028), .o(FE_OFN147_n_25677) );
in01f80 FE_OFC148_n_25677 ( .a(FE_OFN147_n_25677), .o(FE_OFN148_n_25677) );
in01f80 FE_OFC149_n_25677 ( .a(FE_OFN147_n_25677), .o(FE_OFN149_n_25677) );
in01f80 FE_OFC14_n_29068 ( .a(FE_OFN13_n_29068), .o(FE_OFN14_n_29068) );
in01f80 FE_OFC150_n_25677 ( .a(FE_OFN147_n_25677), .o(FE_OFN150_n_25677) );
in01f80 FE_OFC151_n_22615 ( .a(n_22615), .o(FE_OFN151_n_22615) );
in01f80 FE_OFC152_n_22615 ( .a(FE_OFN151_n_22615), .o(FE_OFN152_n_22615) );
in01f80 FE_OFC153_n_22615 ( .a(n_22615), .o(FE_OFN153_n_22615) );
in01f80 FE_OFC154_n_22615 ( .a(FE_OFN153_n_22615), .o(FE_OFN154_n_22615) );
in01f80 FE_OFC155_n_28014 ( .a(FE_OFN340_n_4860), .o(FE_OFN155_n_28014) );
in01f80 FE_OFC156_n_28014 ( .a(FE_OFN155_n_28014), .o(FE_OFN156_n_28014) );
in01f80 FE_OFC157_n_28014 ( .a(FE_OFN155_n_28014), .o(FE_OFN157_n_28014) );
in01f80 FE_OFC158_n_28014 ( .a(FE_OFN155_n_28014), .o(FE_OFN158_n_28014) );
in01f80 FE_OFC159_n_28014 ( .a(FE_OFN156_n_28014), .o(FE_OFN159_n_28014) );
in01f80 FE_OFC15_n_29068 ( .a(FE_OFN13_n_29068), .o(FE_OFN15_n_29068) );
in01f80 FE_OFC160_n_28014 ( .a(FE_OFN159_n_28014), .o(FE_OFN160_n_28014) );
in01f80 FE_OFC161_n_26454 ( .a(n_26454), .o(FE_OFN161_n_26454) );
in01f80 FE_OFC162_n_26454 ( .a(FE_OFN161_n_26454), .o(FE_OFN162_n_26454) );
in01f80 FE_OFC164_n_29269 ( .a(n_29269), .o(FE_OFN164_n_29269) );
in01f80 FE_OFC165_n_29269 ( .a(FE_OFN164_n_29269), .o(FE_OFN165_n_29269) );
in01f80 FE_OFC166_n_29269 ( .a(FE_OFN164_n_29269), .o(FE_OFN166_n_29269) );
in01f80 FE_OFC169_n_22948 ( .a(FE_OFN361_n_4860), .o(FE_OFN169_n_22948) );
in01f80 FE_OFC16_n_29617 ( .a(n_29617), .o(FE_OFN16_n_29617) );
in01f80 FE_OFC170_n_22948 ( .a(FE_OFN361_n_4860), .o(FE_OFN170_n_22948) );
in01f80 FE_OFC171_n_22948 ( .a(FE_OFN361_n_4860), .o(FE_OFN171_n_22948) );
in01f80 FE_OFC172_n_22948 ( .a(FE_OFN169_n_22948), .o(FE_OFN172_n_22948) );
in01f80 FE_OFC173_n_22948 ( .a(FE_OFN172_n_22948), .o(FE_OFN173_n_22948) );
in01f80 FE_OFC174_n_26184 ( .a(n_26184), .o(FE_OFN174_n_26184) );
in01f80 FE_OFC175_n_26184 ( .a(FE_OFN174_n_26184), .o(FE_OFN175_n_26184) );
in01f80 FE_OFC177_n_27681 ( .a(n_27681), .o(FE_OFN177_n_27681) );
in01f80 FE_OFC179_n_27681 ( .a(FE_OFN177_n_27681), .o(FE_OFN179_n_27681) );
in01f80 FE_OFC17_n_29617 ( .a(FE_OFN16_n_29617), .o(FE_OFN17_n_29617) );
in01f80 FE_OFC180_n_27681 ( .a(FE_OFN177_n_27681), .o(FE_OFN180_n_27681) );
in01f80 FE_OFC181_n_27681 ( .a(FE_OFN177_n_27681), .o(FE_OFN181_n_27681) );
in01f80 FE_OFC182_n_29402 ( .a(n_16028), .o(FE_OFN182_n_29402) );
in01f80 FE_OFC183_n_29402 ( .a(FE_OFN182_n_29402), .o(FE_OFN183_n_29402) );
in01f80 FE_OFC184_n_29402 ( .a(FE_OFN182_n_29402), .o(FE_OFN184_n_29402) );
in01f80 FE_OFC185_n_29496 ( .a(n_29496), .o(FE_OFN185_n_29496) );
in01f80 FE_OFC186_n_29496 ( .a(FE_OFN185_n_29496), .o(FE_OFN186_n_29496) );
in01f80 FE_OFC187_n_29496 ( .a(FE_OFN185_n_29496), .o(FE_OFN187_n_29496) );
in01f80 FE_OFC188_n_28362 ( .a(n_28362), .o(FE_OFN188_n_28362) );
in01f80 FE_OFC189_n_28362 ( .a(FE_OFN188_n_28362), .o(FE_OFN189_n_28362) );
in01f80 FE_OFC18_n_29617 ( .a(FE_OFN16_n_29617), .o(FE_OFN18_n_29617) );
in01f80 FE_OFC190_n_28362 ( .a(FE_OFN188_n_28362), .o(FE_OFN190_n_28362) );
in01f80 FE_OFC191_n_28928 ( .a(n_28928), .o(FE_OFN191_n_28928) );
in01f80 FE_OFC192_n_28928 ( .a(FE_OFN191_n_28928), .o(FE_OFN192_n_28928) );
in01f80 FE_OFC193_n_28928 ( .a(FE_OFN191_n_28928), .o(FE_OFN193_n_28928) );
in01f80 FE_OFC195_n_5003 ( .a(n_29104), .o(FE_OFN195_n_5003) );
in01f80 FE_OFC196_n_5003 ( .a(n_29104), .o(FE_OFN196_n_5003) );
in01f80 FE_OFC197_n_29637 ( .a(n_27681), .o(FE_OFN197_n_29637) );
in01f80 FE_OFC198_n_29637 ( .a(FE_OFN197_n_29637), .o(FE_OFN198_n_29637) );
in01f80 FE_OFC199_n_29637 ( .a(FE_OFN197_n_29637), .o(FE_OFN199_n_29637) );
in01f80 FE_OFC19_n_27452 ( .a(n_27452), .o(FE_OFN19_n_27452) );
in01f80 FE_OFC1_n_17395 ( .a(FE_OFN0_n_17395), .o(FE_OFN1_n_17395) );
in01f80 FE_OFC200_n_29637 ( .a(FE_OFN199_n_29637), .o(FE_OFN200_n_29637) );
in01f80 FE_OFC201_n_29637 ( .a(FE_OFN200_n_29637), .o(FE_OFN201_n_29637) );
in01f80 FE_OFC202_n_28771 ( .a(n_28771), .o(FE_OFN202_n_28771) );
in01f80 FE_OFC203_n_28771 ( .a(FE_OFN202_n_28771), .o(FE_OFN203_n_28771) );
in01f80 FE_OFC204_n_28771 ( .a(FE_OFN202_n_28771), .o(FE_OFN204_n_28771) );
in01f80 FE_OFC205_n_28771 ( .a(n_28771), .o(FE_OFN205_n_28771) );
in01f80 FE_OFC206_n_28771 ( .a(FE_OFN205_n_28771), .o(FE_OFN206_n_28771) );
in01f80 FE_OFC207_n_29661 ( .a(n_27681), .o(FE_OFN207_n_29661) );
in01f80 FE_OFC208_n_29661 ( .a(FE_OFN207_n_29661), .o(FE_OFN208_n_29661) );
in01f80 FE_OFC209_n_29661 ( .a(FE_OFN207_n_29661), .o(FE_OFN209_n_29661) );
in01f80 FE_OFC20_n_27452 ( .a(FE_OFN19_n_27452), .o(FE_OFN20_n_27452) );
in01f80 FE_OFC210_n_29661 ( .a(FE_OFN209_n_29661), .o(FE_OFN210_n_29661) );
in01f80 FE_OFC211_n_29661 ( .a(FE_OFN210_n_29661), .o(FE_OFN211_n_29661) );
in01f80 FE_OFC212_n_29661 ( .a(FE_OFN210_n_29661), .o(FE_OFN212_n_29661) );
in01f80 FE_OFC213_n_29687 ( .a(n_29687), .o(FE_OFN213_n_29687) );
in01f80 FE_OFC214_n_29687 ( .a(FE_OFN213_n_29687), .o(FE_OFN214_n_29687) );
in01f80 FE_OFC215_n_29687 ( .a(n_29687), .o(FE_OFN215_n_29687) );
in01f80 FE_OFC217_n_29687 ( .a(FE_OFN215_n_29687), .o(FE_OFN217_n_29687) );
in01f80 FE_OFC218_n_23315 ( .a(n_23315), .o(FE_OFN218_n_23315) );
in01f80 FE_OFC219_n_23315 ( .a(FE_OFN218_n_23315), .o(FE_OFN219_n_23315) );
in01f80 FE_OFC21_n_27452 ( .a(FE_OFN19_n_27452), .o(FE_OFN21_n_27452) );
in01f80 FE_OFC220_n_23315 ( .a(FE_OFN219_n_23315), .o(FE_OFN220_n_23315) );
in01f80 FE_OFC221_n_23315 ( .a(FE_OFN220_n_23315), .o(FE_OFN221_n_23315) );
in01f80 FE_OFC222_n_21642 ( .a(n_29269), .o(FE_OFN222_n_21642) );
in01f80 FE_OFC223_n_21642 ( .a(FE_OFN222_n_21642), .o(FE_OFN223_n_21642) );
in01f80 FE_OFC224_n_21642 ( .a(FE_OFN222_n_21642), .o(FE_OFN224_n_21642) );
in01f80 FE_OFC225_n_21642 ( .a(FE_OFN222_n_21642), .o(FE_OFN225_n_21642) );
in01f80 FE_OFC226_n_4162 ( .a(FE_OFN1165_n_4162), .o(FE_OFN226_n_4162) );
in01f80 FE_OFC227_n_4162 ( .a(FE_OFN1166_n_4162), .o(FE_OFN227_n_4162) );
in01f80 FE_OFC228_n_4162 ( .a(FE_OFN1168_n_4162), .o(FE_OFN228_n_4162) );
in01f80 FE_OFC230_n_4162 ( .a(FE_OFN226_n_4162), .o(FE_OFN230_n_4162) );
in01f80 FE_OFC231_n_4162 ( .a(FE_OFN1166_n_4162), .o(FE_OFN231_n_4162) );
in01f80 FE_OFC232_n_4162 ( .a(FE_OFN1165_n_4162), .o(FE_OFN232_n_4162) );
in01f80 FE_OFC234_n_4162 ( .a(FE_OFN227_n_4162), .o(FE_OFN234_n_4162) );
in01f80 FE_OFC235_n_4162 ( .a(FE_OFN228_n_4162), .o(FE_OFN235_n_4162) );
in01f80 FE_OFC236_n_4162 ( .a(FE_OFN232_n_4162), .o(FE_OFN236_n_4162) );
in01f80 FE_OFC237_n_4162 ( .a(FE_OFN226_n_4162), .o(FE_OFN237_n_4162) );
in01f80 FE_OFC238_n_4162 ( .a(FE_OFN1167_n_4162), .o(FE_OFN238_n_4162) );
in01f80 FE_OFC239_n_4162 ( .a(FE_OFN231_n_4162), .o(FE_OFN239_n_4162) );
in01f80 FE_OFC23_n_26609 ( .a(n_27452), .o(FE_OFN23_n_26609) );
in01f80 FE_OFC240_n_4162 ( .a(FE_OFN231_n_4162), .o(FE_OFN240_n_4162) );
in01f80 FE_OFC242_n_4162 ( .a(FE_OFN237_n_4162), .o(FE_OFN242_n_4162) );
in01f80 FE_OFC243_n_4162 ( .a(FE_OFN237_n_4162), .o(FE_OFN243_n_4162) );
in01f80 FE_OFC244_n_4162 ( .a(FE_OFN238_n_4162), .o(FE_OFN244_n_4162) );
in01f80 FE_OFC247_n_4162 ( .a(FE_OFN227_n_4162), .o(FE_OFN247_n_4162) );
in01f80 FE_OFC248_n_4162 ( .a(FE_OFN242_n_4162), .o(FE_OFN248_n_4162) );
in01f80 FE_OFC249_n_4162 ( .a(FE_OFN243_n_4162), .o(FE_OFN249_n_4162) );
in01f80 FE_OFC24_n_11489 ( .a(n_11489), .o(FE_OFN24_n_11489) );
in01f80 FE_OFC251_n_4162 ( .a(FE_OFN242_n_4162), .o(FE_OFN251_n_4162) );
in01f80 FE_OFC252_n_4280 ( .a(n_4280), .o(FE_OFN252_n_4280) );
in01f80 FE_OFC253_n_4280 ( .a(FE_OFN252_n_4280), .o(FE_OFN253_n_4280) );
in01f80 FE_OFC254_n_4280 ( .a(FE_OFN252_n_4280), .o(FE_OFN254_n_4280) );
in01f80 FE_OFC256_n_4280 ( .a(FE_OFN252_n_4280), .o(FE_OFN256_n_4280) );
in01f80 FE_OFC257_n_4280 ( .a(FE_OFN252_n_4280), .o(FE_OFN257_n_4280) );
in01f80 FE_OFC258_n_4280 ( .a(FE_OFN252_n_4280), .o(FE_OFN258_n_4280) );
in01f80 FE_OFC259_n_4280 ( .a(FE_OFN252_n_4280), .o(FE_OFN259_n_4280) );
in01f80 FE_OFC25_n_11489 ( .a(FE_OFN24_n_11489), .o(FE_OFN25_n_11489) );
in01f80 FE_OFC260_n_4280 ( .a(FE_OFN252_n_4280), .o(FE_OFN260_n_4280) );
in01f80 FE_OFC261_n_4280 ( .a(FE_OFN258_n_4280), .o(FE_OFN261_n_4280) );
in01f80 FE_OFC262_n_4280 ( .a(FE_OFN258_n_4280), .o(FE_OFN262_n_4280) );
in01f80 FE_OFC264_n_4280 ( .a(FE_OFN261_n_4280), .o(FE_OFN264_n_4280) );
in01f80 FE_OFC265_n_4280 ( .a(FE_OFN262_n_4280), .o(FE_OFN265_n_4280) );
in01f80 FE_OFC266_n_4280 ( .a(FE_OFN261_n_4280), .o(FE_OFN266_n_4280) );
in01f80 FE_OFC267_n_4280 ( .a(FE_OFN261_n_4280), .o(FE_OFN267_n_4280) );
in01f80 FE_OFC268_n_4280 ( .a(FE_OFN261_n_4280), .o(FE_OFN268_n_4280) );
in01f80 FE_OFC269_n_4280 ( .a(FE_OFN261_n_4280), .o(FE_OFN269_n_4280) );
in01f80 FE_OFC26_n_13676 ( .a(n_13676), .o(FE_OFN26_n_13676) );
in01f80 FE_OFC270_n_16028 ( .a(n_16028), .o(FE_OFN270_n_16028) );
in01f80 FE_OFC271_n_16028 ( .a(FE_OFN270_n_16028), .o(FE_OFN271_n_16028) );
in01f80 FE_OFC272_n_16893 ( .a(n_16893), .o(FE_OFN272_n_16893) );
in01f80 FE_OFC273_n_16893 ( .a(FE_OFN272_n_16893), .o(FE_OFN273_n_16893) );
in01f80 FE_OFC274_n_16893 ( .a(FE_OFN272_n_16893), .o(FE_OFN274_n_16893) );
in01f80 FE_OFC275_n_16893 ( .a(n_16893), .o(FE_OFN275_n_16893) );
in01f80 FE_OFC276_n_16893 ( .a(FE_OFN275_n_16893), .o(FE_OFN276_n_16893) );
in01f80 FE_OFC277_n_16893 ( .a(FE_OFN275_n_16893), .o(FE_OFN277_n_16893) );
in01f80 FE_OFC278_n_16656 ( .a(n_16656), .o(FE_OFN278_n_16656) );
in01f80 FE_OFC279_n_16656 ( .a(FE_OFN278_n_16656), .o(FE_OFN279_n_16656) );
in01f80 FE_OFC27_n_13676 ( .a(FE_OFN26_n_13676), .o(FE_OFN27_n_13676) );
in01f80 FE_OFC280_n_16656 ( .a(FE_OFN278_n_16656), .o(FE_OFN280_n_16656) );
in01f80 FE_OFC281_n_7349 ( .a(n_7349), .o(FE_OFN281_n_7349) );
in01f80 FE_OFC282_n_7349 ( .a(FE_OFN281_n_7349), .o(FE_OFN282_n_7349) );
in01f80 FE_OFC283_n_29266 ( .a(n_29266), .o(FE_OFN283_n_29266) );
in01f80 FE_OFC284_n_29266 ( .a(n_29266), .o(FE_OFN284_n_29266) );
in01f80 FE_OFC285_n_29266 ( .a(FE_OFN283_n_29266), .o(FE_OFN285_n_29266) );
in01f80 FE_OFC286_n_29266 ( .a(FE_OFN283_n_29266), .o(FE_OFN286_n_29266) );
in01f80 FE_OFC287_n_29266 ( .a(FE_OFN284_n_29266), .o(FE_OFN287_n_29266) );
in01f80 FE_OFC288_n_29266 ( .a(FE_OFN284_n_29266), .o(FE_OFN288_n_29266) );
in01f80 FE_OFC289_n_27194 ( .a(n_27194), .o(FE_OFN289_n_27194) );
in01f80 FE_OFC28_n_13676 ( .a(FE_OFN26_n_13676), .o(FE_OFN28_n_13676) );
in01f80 FE_OFC290_n_27194 ( .a(FE_OFN289_n_27194), .o(FE_OFN290_n_27194) );
in01f80 FE_OFC291_n_3069 ( .a(n_4280), .o(FE_OFN291_n_3069) );
in01f80 FE_OFC292_n_3069 ( .a(FE_OFN291_n_3069), .o(FE_OFN292_n_3069) );
in01f80 FE_OFC293_n_3069 ( .a(FE_OFN291_n_3069), .o(FE_OFN293_n_3069) );
in01f80 FE_OFC294_n_3069 ( .a(FE_OFN291_n_3069), .o(FE_OFN294_n_3069) );
in01f80 FE_OFC295_n_3069 ( .a(FE_OFN291_n_3069), .o(FE_OFN295_n_3069) );
in01f80 FE_OFC296_n_3069 ( .a(FE_OFN291_n_3069), .o(FE_OFN296_n_3069) );
in01f80 FE_OFC297_n_3069 ( .a(FE_OFN291_n_3069), .o(FE_OFN297_n_3069) );
in01f80 FE_OFC298_n_3069 ( .a(FE_OFN293_n_3069), .o(FE_OFN298_n_3069) );
in01f80 FE_OFC299_n_3069 ( .a(FE_OFN291_n_3069), .o(FE_OFN299_n_3069) );
in01f80 FE_OFC29_n_13676 ( .a(FE_OFN26_n_13676), .o(FE_OFN29_n_13676) );
in01f80 FE_OFC2_n_28682 ( .a(n_28682), .o(FE_OFN2_n_28682) );
in01f80 FE_OFC300_n_3069 ( .a(FE_OFN291_n_3069), .o(FE_OFN300_n_3069) );
in01f80 FE_OFC301_n_3069 ( .a(FE_OFN296_n_3069), .o(FE_OFN301_n_3069) );
in01f80 FE_OFC302_n_3069 ( .a(FE_OFN295_n_3069), .o(FE_OFN302_n_3069) );
in01f80 FE_OFC303_n_3069 ( .a(FE_OFN298_n_3069), .o(FE_OFN303_n_3069) );
in01f80 FE_OFC304_n_3069 ( .a(FE_OFN296_n_3069), .o(FE_OFN304_n_3069) );
in01f80 FE_OFC305_n_3069 ( .a(FE_OFN300_n_3069), .o(FE_OFN305_n_3069) );
in01f80 FE_OFC306_n_3069 ( .a(FE_OFN302_n_3069), .o(FE_OFN306_n_3069) );
in01f80 FE_OFC307_n_3069 ( .a(FE_OFN302_n_3069), .o(FE_OFN307_n_3069) );
in01f80 FE_OFC308_n_3069 ( .a(FE_OFN301_n_3069), .o(FE_OFN308_n_3069) );
in01f80 FE_OFC309_n_3069 ( .a(FE_OFN301_n_3069), .o(FE_OFN309_n_3069) );
in01f80 FE_OFC30_n_13676 ( .a(FE_OFN26_n_13676), .o(FE_OFN30_n_13676) );
in01f80 FE_OFC310_n_3069 ( .a(FE_OFN301_n_3069), .o(FE_OFN310_n_3069) );
in01f80 FE_OFC311_n_3069 ( .a(FE_OFN304_n_3069), .o(FE_OFN311_n_3069) );
in01f80 FE_OFC312_n_3069 ( .a(FE_OFN305_n_3069), .o(FE_OFN312_n_3069) );
in01f80 FE_OFC313_n_3069 ( .a(FE_OFN304_n_3069), .o(FE_OFN313_n_3069) );
in01f80 FE_OFC314_n_3069 ( .a(FE_OFN305_n_3069), .o(FE_OFN314_n_3069) );
in01f80 FE_OFC315_n_26999 ( .a(n_26999), .o(FE_OFN315_n_26999) );
in01f80 FE_OFC316_n_26999 ( .a(FE_OFN315_n_26999), .o(FE_OFN316_n_26999) );
in01f80 FE_OFC317_n_27400 ( .a(n_27400), .o(FE_OFN317_n_27400) );
in01f80 FE_OFC318_n_27400 ( .a(FE_OFN317_n_27400), .o(FE_OFN318_n_27400) );
in01f80 FE_OFC320_n_4860 ( .a(FE_OFN1172_n_4860), .o(FE_OFN320_n_4860) );
in01f80 FE_OFC321_n_4860 ( .a(n_4860), .o(FE_OFN321_n_4860) );
in01f80 FE_OFC322_n_4860 ( .a(n_4860), .o(FE_OFN322_n_4860) );
in01f80 FE_OFC324_n_4860 ( .a(FE_OFN320_n_4860), .o(FE_OFN324_n_4860) );
in01f80 FE_OFC325_n_4860 ( .a(FE_OFN1173_n_4860), .o(FE_OFN325_n_4860) );
in01f80 FE_OFC326_n_4860 ( .a(FE_OFN321_n_4860), .o(FE_OFN326_n_4860) );
in01f80 FE_OFC327_n_4860 ( .a(FE_OFN1171_n_4860), .o(FE_OFN327_n_4860) );
in01f80 FE_OFC329_n_4860 ( .a(FE_OFN321_n_4860), .o(FE_OFN329_n_4860) );
in01f80 FE_OFC32_n_27986 ( .a(FE_OFN1130_n_27986), .o(FE_OFN32_n_27986) );
in01f80 FE_OFC330_n_4860 ( .a(FE_OFN321_n_4860), .o(FE_OFN330_n_4860) );
in01f80 FE_OFC331_n_4860 ( .a(FE_OFN322_n_4860), .o(FE_OFN331_n_4860) );
in01f80 FE_OFC332_n_4860 ( .a(FE_OFN322_n_4860), .o(FE_OFN332_n_4860) );
in01f80 FE_OFC334_n_4860 ( .a(FE_OFN325_n_4860), .o(FE_OFN334_n_4860) );
in01f80 FE_OFC335_n_4860 ( .a(FE_OFN327_n_4860), .o(FE_OFN335_n_4860) );
in01f80 FE_OFC336_n_4860 ( .a(FE_OFN327_n_4860), .o(FE_OFN336_n_4860) );
in01f80 FE_OFC337_n_4860 ( .a(FE_OFN1171_n_4860), .o(FE_OFN337_n_4860) );
in01f80 FE_OFC338_n_4860 ( .a(FE_OFN1171_n_4860), .o(FE_OFN338_n_4860) );
in01f80 FE_OFC339_n_4860 ( .a(FE_OFN331_n_4860), .o(FE_OFN339_n_4860) );
in01f80 FE_OFC33_n_15183 ( .a(n_15183), .o(FE_OFN33_n_15183) );
in01f80 FE_OFC340_n_4860 ( .a(FE_OFN332_n_4860), .o(FE_OFN340_n_4860) );
in01f80 FE_OFC341_n_4860 ( .a(FE_OFN335_n_4860), .o(FE_OFN341_n_4860) );
in01f80 FE_OFC342_n_4860 ( .a(FE_OFN334_n_4860), .o(FE_OFN342_n_4860) );
in01f80 FE_OFC343_n_4860 ( .a(FE_OFN334_n_4860), .o(FE_OFN343_n_4860) );
in01f80 FE_OFC344_n_4860 ( .a(FE_OFN334_n_4860), .o(FE_OFN344_n_4860) );
in01f80 FE_OFC345_n_4860 ( .a(FE_OFN337_n_4860), .o(FE_OFN345_n_4860) );
in01f80 FE_OFC347_n_4860 ( .a(FE_OFN338_n_4860), .o(FE_OFN347_n_4860) );
in01f80 FE_OFC349_n_4860 ( .a(FE_OFN340_n_4860), .o(FE_OFN349_n_4860) );
in01f80 FE_OFC34_n_15183 ( .a(FE_OFN33_n_15183), .o(FE_OFN34_n_15183) );
in01f80 FE_OFC350_n_4860 ( .a(FE_OFN339_n_4860), .o(FE_OFN350_n_4860) );
in01f80 FE_OFC352_n_4860 ( .a(FE_OFN339_n_4860), .o(FE_OFN352_n_4860) );
in01f80 FE_OFC353_n_4860 ( .a(FE_OFN341_n_4860), .o(FE_OFN353_n_4860) );
in01f80 FE_OFC355_n_4860 ( .a(FE_OFN342_n_4860), .o(FE_OFN355_n_4860) );
in01f80 FE_OFC357_n_4860 ( .a(FE_OFN343_n_4860), .o(FE_OFN357_n_4860) );
in01f80 FE_OFC358_n_4860 ( .a(FE_OFN344_n_4860), .o(FE_OFN358_n_4860) );
in01f80 FE_OFC359_n_4860 ( .a(FE_OFN345_n_4860), .o(FE_OFN359_n_4860) );
in01f80 FE_OFC35_n_15183 ( .a(FE_OFN33_n_15183), .o(FE_OFN35_n_15183) );
in01f80 FE_OFC360_n_4860 ( .a(FE_OFN342_n_4860), .o(FE_OFN360_n_4860) );
in01f80 FE_OFC361_n_4860 ( .a(FE_OFN344_n_4860), .o(FE_OFN361_n_4860) );
in01f80 FE_OFC363_n_4860 ( .a(FE_OFN339_n_4860), .o(FE_OFN363_n_4860) );
in01f80 FE_OFC364_n_4860 ( .a(FE_OFN359_n_4860), .o(FE_OFN364_n_4860) );
in01f80 FE_OFC368_n_26312 ( .a(n_27449), .o(FE_OFN368_n_26312) );
in01f80 FE_OFC369_n_26312 ( .a(n_27449), .o(FE_OFN369_n_26312) );
in01f80 FE_OFC370_n_15817 ( .a(n_15817), .o(FE_OFN370_n_15817) );
in01f80 FE_OFC371_n_15817 ( .a(FE_OFN370_n_15817), .o(FE_OFN371_n_15817) );
in01f80 FE_OFC372_n_15853 ( .a(n_15853), .o(FE_OFN372_n_15853) );
in01f80 FE_OFC373_n_15853 ( .a(FE_OFN372_n_15853), .o(FE_OFN373_n_15853) );
in01f80 FE_OFC374_n_14224 ( .a(n_14224), .o(FE_OFN374_n_14224) );
in01f80 FE_OFC375_n_14224 ( .a(FE_OFN374_n_14224), .o(FE_OFN375_n_14224) );
in01f80 FE_OFC376_n_14285 ( .a(n_14285), .o(FE_OFN376_n_14285) );
in01f80 FE_OFC377_n_14285 ( .a(FE_OFN376_n_14285), .o(FE_OFN377_n_14285) );
in01f80 FE_OFC378_n_13985 ( .a(n_13985), .o(FE_OFN378_n_13985) );
in01f80 FE_OFC379_n_13985 ( .a(FE_OFN378_n_13985), .o(FE_OFN379_n_13985) );
in01f80 FE_OFC37_n_17184 ( .a(n_13676), .o(FE_OFN37_n_17184) );
in01f80 FE_OFC380_n_16289 ( .a(n_16289), .o(FE_OFN380_n_16289) );
in01f80 FE_OFC381_n_16289 ( .a(n_16289), .o(FE_OFN381_n_16289) );
in01f80 FE_OFC382_n_16289 ( .a(FE_OFN380_n_16289), .o(FE_OFN382_n_16289) );
in01f80 FE_OFC383_n_16289 ( .a(FE_OFN380_n_16289), .o(FE_OFN383_n_16289) );
in01f80 FE_OFC384_n_16289 ( .a(FE_OFN381_n_16289), .o(FE_OFN384_n_16289) );
in01f80 FE_OFC385_n_16289 ( .a(FE_OFN381_n_16289), .o(FE_OFN385_n_16289) );
in01f80 FE_OFC386_n_17236 ( .a(n_17236), .o(FE_OFN386_n_17236) );
in01f80 FE_OFC387_n_17236 ( .a(FE_OFN386_n_17236), .o(FE_OFN387_n_17236) );
in01f80 FE_OFC388_n_16991 ( .a(n_16991), .o(FE_OFN388_n_16991) );
in01f80 FE_OFC389_n_16991 ( .a(FE_OFN388_n_16991), .o(FE_OFN389_n_16991) );
in01f80 FE_OFC38_n_17184 ( .a(n_13676), .o(FE_OFN38_n_17184) );
in01f80 FE_OFC390_n_15554 ( .a(n_15554), .o(FE_OFN390_n_15554) );
in01f80 FE_OFC391_n_15554 ( .a(FE_OFN390_n_15554), .o(FE_OFN391_n_15554) );
in01f80 FE_OFC392_n_14663 ( .a(n_14663), .o(FE_OFN392_n_14663) );
in01f80 FE_OFC393_n_14663 ( .a(FE_OFN392_n_14663), .o(FE_OFN393_n_14663) );
in01f80 FE_OFC394_n_14720 ( .a(n_14720), .o(FE_OFN394_n_14720) );
in01f80 FE_OFC396_n_14720 ( .a(FE_OFN394_n_14720), .o(FE_OFN396_n_14720) );
in01f80 FE_OFC397_n_8616 ( .a(n_8616), .o(FE_OFN397_n_8616) );
in01f80 FE_OFC398_n_8616 ( .a(FE_OFN397_n_8616), .o(FE_OFN398_n_8616) );
in01f80 FE_OFC399_n_28303 ( .a(n_28303), .o(FE_OFN399_n_28303) );
in01f80 FE_OFC39_n_25450 ( .a(n_25450), .o(FE_OFN39_n_25450) );
in01f80 FE_OFC3_n_28682 ( .a(FE_OFN2_n_28682), .o(FE_OFN3_n_28682) );
in01f80 FE_OFC400_n_28303 ( .a(FE_OFN399_n_28303), .o(FE_OFN400_n_28303) );
in01f80 FE_OFC402_n_28303 ( .a(FE_OFN399_n_28303), .o(FE_OFN402_n_28303) );
in01f80 FE_OFC404_n_28303 ( .a(FE_OFN399_n_28303), .o(FE_OFN404_n_28303) );
in01f80 FE_OFC405_n_28303 ( .a(FE_OFN399_n_28303), .o(FE_OFN405_n_28303) );
in01f80 FE_OFC406_n_28303 ( .a(FE_OFN399_n_28303), .o(FE_OFN406_n_28303) );
in01f80 FE_OFC407_n_28303 ( .a(FE_OFN406_n_28303), .o(FE_OFN407_n_28303) );
in01f80 FE_OFC408_n_28303 ( .a(FE_OFN406_n_28303), .o(FE_OFN408_n_28303) );
in01f80 FE_OFC409_n_28303 ( .a(FE_OFN399_n_28303), .o(FE_OFN409_n_28303) );
in01f80 FE_OFC40_n_25450 ( .a(FE_OFN39_n_25450), .o(FE_OFN40_n_25450) );
in01f80 FE_OFC410_n_28303 ( .a(FE_OFN399_n_28303), .o(FE_OFN410_n_28303) );
in01f80 FE_OFC411_n_28303 ( .a(FE_OFN408_n_28303), .o(FE_OFN411_n_28303) );
in01f80 FE_OFC412_n_28303 ( .a(FE_OFN408_n_28303), .o(FE_OFN412_n_28303) );
in01f80 FE_OFC413_n_28303 ( .a(FE_OFN407_n_28303), .o(FE_OFN413_n_28303) );
in01f80 FE_OFC414_n_28303 ( .a(FE_OFN408_n_28303), .o(FE_OFN414_n_28303) );
in01f80 FE_OFC416_n_28303 ( .a(FE_OFN407_n_28303), .o(FE_OFN416_n_28303) );
in01f80 FE_OFC417_n_28303 ( .a(FE_OFN407_n_28303), .o(FE_OFN417_n_28303) );
in01f80 FE_OFC419_n_16909 ( .a(n_28303), .o(FE_OFN419_n_16909) );
in01f80 FE_OFC41_n_26563 ( .a(n_26563), .o(FE_OFN41_n_26563) );
in01f80 FE_OFC420_n_16909 ( .a(n_16909), .o(FE_OFN420_n_16909) );
in01f80 FE_OFC421_n_16909 ( .a(FE_OFN420_n_16909), .o(FE_OFN421_n_16909) );
in01f80 FE_OFC422_n_16909 ( .a(FE_OFN420_n_16909), .o(FE_OFN422_n_16909) );
in01f80 FE_OFC423_n_16296 ( .a(n_16296), .o(FE_OFN423_n_16296) );
in01f80 FE_OFC424_n_16296 ( .a(FE_OFN423_n_16296), .o(FE_OFN424_n_16296) );
in01f80 FE_OFC425_n_23661 ( .a(n_23661), .o(FE_OFN425_n_23661) );
in01f80 FE_OFC426_n_23661 ( .a(FE_OFN425_n_23661), .o(FE_OFN426_n_23661) );
in01f80 FE_OFC427_n_17707 ( .a(n_17707), .o(FE_OFN427_n_17707) );
in01f80 FE_OFC428_n_17707 ( .a(FE_OFN427_n_17707), .o(FE_OFN428_n_17707) );
in01f80 FE_OFC429_n_26458 ( .a(n_26458), .o(FE_OFN429_n_26458) );
in01f80 FE_OFC42_n_26563 ( .a(FE_OFN41_n_26563), .o(FE_OFN42_n_26563) );
in01f80 FE_OFC430_n_26458 ( .a(FE_OFN429_n_26458), .o(FE_OFN430_n_26458) );
in01f80 FE_OFC431_n_20518 ( .a(n_20518), .o(FE_OFN431_n_20518) );
in01f80 FE_OFC432_n_20518 ( .a(FE_OFN431_n_20518), .o(FE_OFN432_n_20518) );
in01f80 FE_OFC433_n_23637 ( .a(n_23637), .o(FE_OFN433_n_23637) );
in01f80 FE_OFC434_n_23637 ( .a(FE_OFN433_n_23637), .o(FE_OFN434_n_23637) );
in01f80 FE_OFC435_n_26167 ( .a(n_26167), .o(FE_OFN435_n_26167) );
in01f80 FE_OFC436_n_26167 ( .a(FE_OFN435_n_26167), .o(FE_OFN436_n_26167) );
in01f80 FE_OFC437_n_27889 ( .a(n_27889), .o(FE_OFN437_n_27889) );
in01f80 FE_OFC438_n_27889 ( .a(FE_OFN437_n_27889), .o(FE_OFN438_n_27889) );
in01f80 FE_OFC43_n_25810 ( .a(n_25810), .o(FE_OFN43_n_25810) );
in01f80 FE_OFC443_n_19118 ( .a(n_19118), .o(FE_OFN443_n_19118) );
in01f80 FE_OFC444_n_19118 ( .a(FE_OFN443_n_19118), .o(FE_OFN444_n_19118) );
in01f80 FE_OFC445_n_24948 ( .a(n_24948), .o(FE_OFN445_n_24948) );
in01f80 FE_OFC446_n_24948 ( .a(FE_OFN445_n_24948), .o(FE_OFN446_n_24948) );
in01f80 FE_OFC449_n_17680 ( .a(n_17680), .o(FE_OFN449_n_17680) );
in01f80 FE_OFC44_n_25810 ( .a(FE_OFN43_n_25810), .o(FE_OFN44_n_25810) );
in01f80 FE_OFC450_n_17680 ( .a(FE_OFN449_n_17680), .o(FE_OFN450_n_17680) );
in01f80 FE_OFC451_n_23152 ( .a(n_23152), .o(FE_OFN451_n_23152) );
in01f80 FE_OFC452_n_23152 ( .a(FE_OFN451_n_23152), .o(FE_OFN452_n_23152) );
in01f80 FE_OFC453_n_24837 ( .a(n_24837), .o(FE_OFN453_n_24837) );
in01f80 FE_OFC454_n_24837 ( .a(FE_OFN453_n_24837), .o(FE_OFN454_n_24837) );
in01f80 FE_OFC455_n_8508 ( .a(n_8508), .o(FE_OFN455_n_8508) );
in01f80 FE_OFC456_n_8508 ( .a(FE_OFN455_n_8508), .o(FE_OFN456_n_8508) );
in01f80 FE_OFC457_n_5621 ( .a(n_5621), .o(FE_OFN457_n_5621) );
in01f80 FE_OFC458_n_5621 ( .a(FE_OFN457_n_5621), .o(FE_OFN458_n_5621) );
in01f80 FE_OFC459_n_13371 ( .a(n_13371), .o(FE_OFN459_n_13371) );
in01f80 FE_OFC45_n_17233 ( .a(n_17233), .o(FE_OFN45_n_17233) );
in01f80 FE_OFC460_n_13371 ( .a(FE_OFN459_n_13371), .o(FE_OFN460_n_13371) );
in01f80 FE_OFC461_n_21334 ( .a(n_21334), .o(FE_OFN461_n_21334) );
in01f80 FE_OFC462_n_21334 ( .a(FE_OFN461_n_21334), .o(FE_OFN462_n_21334) );
in01f80 FE_OFC46_n_17233 ( .a(FE_OFN45_n_17233), .o(FE_OFN46_n_17233) );
in01f80 FE_OFC473_n_5257 ( .a(n_5257), .o(FE_OFN473_n_5257) );
in01f80 FE_OFC474_n_5257 ( .a(FE_OFN473_n_5257), .o(FE_OFN474_n_5257) );
in01f80 FE_OFC477_n_11170 ( .a(n_11170), .o(FE_OFN477_n_11170) );
in01f80 FE_OFC478_n_11170 ( .a(FE_OFN477_n_11170), .o(FE_OFN478_n_11170) );
in01f80 FE_OFC479_n_12184 ( .a(n_12184), .o(FE_OFN479_n_12184) );
in01f80 FE_OFC47_n_17099 ( .a(n_17099), .o(FE_OFN47_n_17099) );
in01f80 FE_OFC480_n_12184 ( .a(FE_OFN479_n_12184), .o(FE_OFN480_n_12184) );
in01f80 FE_OFC481_n_13520 ( .a(n_13520), .o(FE_OFN481_n_13520) );
in01f80 FE_OFC482_n_13520 ( .a(FE_OFN481_n_13520), .o(FE_OFN482_n_13520) );
in01f80 FE_OFC483_n_12038 ( .a(n_12038), .o(FE_OFN483_n_12038) );
in01f80 FE_OFC484_n_12038 ( .a(FE_OFN483_n_12038), .o(FE_OFN484_n_12038) );
in01f80 FE_OFC485_n_17500 ( .a(n_17500), .o(FE_OFN485_n_17500) );
in01f80 FE_OFC486_n_17500 ( .a(FE_OFN485_n_17500), .o(FE_OFN486_n_17500) );
in01f80 FE_OFC487_n_27256 ( .a(n_27256), .o(FE_OFN487_n_27256) );
in01f80 FE_OFC488_n_27256 ( .a(FE_OFN487_n_27256), .o(FE_OFN488_n_27256) );
in01f80 FE_OFC489_n_20516 ( .a(n_20516), .o(FE_OFN489_n_20516) );
in01f80 FE_OFC48_n_17099 ( .a(FE_OFN47_n_17099), .o(FE_OFN48_n_17099) );
in01f80 FE_OFC490_n_20516 ( .a(FE_OFN489_n_20516), .o(FE_OFN490_n_20516) );
in01f80 FE_OFC491_n_28765 ( .a(n_28765), .o(FE_OFN491_n_28765) );
in01f80 FE_OFC492_n_28765 ( .a(FE_OFN491_n_28765), .o(FE_OFN492_n_28765) );
in01f80 FE_OFC493_n_18414 ( .a(n_18414), .o(FE_OFN493_n_18414) );
in01f80 FE_OFC494_n_18414 ( .a(FE_OFN493_n_18414), .o(FE_OFN494_n_18414) );
in01f80 FE_OFC495_n_21648 ( .a(n_21648), .o(FE_OFN495_n_21648) );
in01f80 FE_OFC496_n_21648 ( .a(FE_OFN495_n_21648), .o(FE_OFN496_n_21648) );
in01f80 FE_OFC497_n_20677 ( .a(n_20677), .o(FE_OFN497_n_20677) );
in01f80 FE_OFC498_n_20677 ( .a(FE_OFN497_n_20677), .o(FE_OFN498_n_20677) );
in01f80 FE_OFC4_n_28682 ( .a(FE_OFN2_n_28682), .o(FE_OFN4_n_28682) );
in01f80 FE_OFC507_n_22083 ( .a(n_22083), .o(FE_OFN507_n_22083) );
in01f80 FE_OFC508_n_22083 ( .a(FE_OFN507_n_22083), .o(FE_OFN508_n_22083) );
in01f80 FE_OFC511_n_19847 ( .a(n_19847), .o(FE_OFN511_n_19847) );
in01f80 FE_OFC512_n_19847 ( .a(FE_OFN511_n_19847), .o(FE_OFN512_n_19847) );
in01f80 FE_OFC513_n_23620 ( .a(n_23620), .o(FE_OFN513_n_23620) );
in01f80 FE_OFC514_n_23620 ( .a(FE_OFN513_n_23620), .o(FE_OFN514_n_23620) );
in01f80 FE_OFC515_n_28406 ( .a(n_28406), .o(FE_OFN515_n_28406) );
in01f80 FE_OFC516_n_28406 ( .a(FE_OFN515_n_28406), .o(FE_OFN516_n_28406) );
in01f80 FE_OFC517_n_20894 ( .a(n_20894), .o(FE_OFN517_n_20894) );
in01f80 FE_OFC518_n_20894 ( .a(FE_OFN517_n_20894), .o(FE_OFN518_n_20894) );
in01f80 FE_OFC519_n_22315 ( .a(n_22315), .o(FE_OFN519_n_22315) );
in01f80 FE_OFC51_n_27012 ( .a(n_27012), .o(FE_OFN51_n_27012) );
in01f80 FE_OFC520_n_22315 ( .a(FE_OFN519_n_22315), .o(FE_OFN520_n_22315) );
in01f80 FE_OFC521_n_25685 ( .a(n_25685), .o(FE_OFN521_n_25685) );
in01f80 FE_OFC522_n_25685 ( .a(FE_OFN521_n_25685), .o(FE_OFN522_n_25685) );
in01f80 FE_OFC523_n_21282 ( .a(n_21282), .o(FE_OFN523_n_21282) );
in01f80 FE_OFC524_n_21282 ( .a(FE_OFN523_n_21282), .o(FE_OFN524_n_21282) );
in01f80 FE_OFC529_n_16938 ( .a(n_16938), .o(FE_OFN529_n_16938) );
in01f80 FE_OFC530_n_16938 ( .a(FE_OFN529_n_16938), .o(FE_OFN530_n_16938) );
in01f80 FE_OFC531_n_12317 ( .a(n_12317), .o(FE_OFN531_n_12317) );
in01f80 FE_OFC532_n_12317 ( .a(FE_OFN531_n_12317), .o(FE_OFN532_n_12317) );
in01f80 FE_OFC533_n_13775 ( .a(n_13775), .o(FE_OFN533_n_13775) );
in01f80 FE_OFC534_n_13775 ( .a(FE_OFN533_n_13775), .o(FE_OFN534_n_13775) );
in01f80 FE_OFC535_n_17798 ( .a(n_17798), .o(FE_OFN535_n_17798) );
in01f80 FE_OFC536_n_17798 ( .a(FE_OFN535_n_17798), .o(FE_OFN536_n_17798) );
in01f80 FE_OFC537_n_10328 ( .a(n_10328), .o(FE_OFN537_n_10328) );
in01f80 FE_OFC538_n_10328 ( .a(FE_OFN537_n_10328), .o(FE_OFN538_n_10328) );
in01f80 FE_OFC539_n_17809 ( .a(n_17809), .o(FE_OFN539_n_17809) );
in01f80 FE_OFC540_n_17809 ( .a(FE_OFN539_n_17809), .o(FE_OFN540_n_17809) );
in01f80 FE_OFC541_n_23570 ( .a(n_23570), .o(FE_OFN541_n_23570) );
in01f80 FE_OFC542_n_23570 ( .a(FE_OFN541_n_23570), .o(FE_OFN542_n_23570) );
in01f80 FE_OFC543_n_9030 ( .a(n_9030), .o(FE_OFN543_n_9030) );
in01f80 FE_OFC544_n_9030 ( .a(FE_OFN543_n_9030), .o(FE_OFN544_n_9030) );
in01f80 FE_OFC545_n_9036 ( .a(n_9036), .o(FE_OFN545_n_9036) );
in01f80 FE_OFC546_n_9036 ( .a(FE_OFN545_n_9036), .o(FE_OFN546_n_9036) );
in01f80 FE_OFC547_n_10452 ( .a(n_10452), .o(FE_OFN547_n_10452) );
in01f80 FE_OFC548_n_10452 ( .a(FE_OFN547_n_10452), .o(FE_OFN548_n_10452) );
in01f80 FE_OFC549_n_6072 ( .a(n_6072), .o(FE_OFN549_n_6072) );
in01f80 FE_OFC54_n_27012 ( .a(n_27012), .o(FE_OFN54_n_27012) );
in01f80 FE_OFC550_n_6072 ( .a(FE_OFN549_n_6072), .o(FE_OFN550_n_6072) );
in01f80 FE_OFC551_n_9482 ( .a(n_9482), .o(FE_OFN551_n_9482) );
in01f80 FE_OFC552_n_9482 ( .a(FE_OFN551_n_9482), .o(FE_OFN552_n_9482) );
in01f80 FE_OFC553_n_9468 ( .a(n_9468), .o(FE_OFN553_n_9468) );
in01f80 FE_OFC554_n_9468 ( .a(FE_OFN553_n_9468), .o(FE_OFN554_n_9468) );
in01f80 FE_OFC555_n_23580 ( .a(n_23580), .o(FE_OFN555_n_23580) );
in01f80 FE_OFC556_n_23580 ( .a(FE_OFN555_n_23580), .o(FE_OFN556_n_23580) );
in01f80 FE_OFC557_n_26546 ( .a(n_26546), .o(FE_OFN557_n_26546) );
in01f80 FE_OFC558_n_26546 ( .a(FE_OFN557_n_26546), .o(FE_OFN558_n_26546) );
in01f80 FE_OFC56_n_27012 ( .a(FE_OFN61_n_27012), .o(FE_OFN56_n_27012) );
in01f80 FE_OFC571_n_12800 ( .a(n_12800), .o(FE_OFN571_n_12800) );
in01f80 FE_OFC572_n_12800 ( .a(FE_OFN571_n_12800), .o(FE_OFN572_n_12800) );
in01f80 FE_OFC573_n_10137 ( .a(n_10137), .o(FE_OFN573_n_10137) );
in01f80 FE_OFC574_n_10137 ( .a(FE_OFN573_n_10137), .o(FE_OFN574_n_10137) );
in01f80 FE_OFC575_n_10136 ( .a(n_10136), .o(FE_OFN575_n_10136) );
in01f80 FE_OFC576_n_10136 ( .a(FE_OFN575_n_10136), .o(FE_OFN576_n_10136) );
in01f80 FE_OFC577_n_6424 ( .a(n_6424), .o(FE_OFN577_n_6424) );
in01f80 FE_OFC578_n_6424 ( .a(FE_OFN577_n_6424), .o(FE_OFN578_n_6424) );
in01f80 FE_OFC579_n_19119 ( .a(n_19119), .o(FE_OFN579_n_19119) );
in01f80 FE_OFC57_n_27012 ( .a(n_27012), .o(FE_OFN57_n_27012) );
in01f80 FE_OFC580_n_19119 ( .a(FE_OFN579_n_19119), .o(FE_OFN580_n_19119) );
in01f80 FE_OFC583_n_18103 ( .a(n_18103), .o(FE_OFN583_n_18103) );
in01f80 FE_OFC584_n_18103 ( .a(FE_OFN583_n_18103), .o(FE_OFN584_n_18103) );
in01f80 FE_OFC585_n_19447 ( .a(n_19447), .o(FE_OFN585_n_19447) );
in01f80 FE_OFC586_n_19447 ( .a(FE_OFN585_n_19447), .o(FE_OFN586_n_19447) );
in01f80 FE_OFC589_n_20904 ( .a(n_20904), .o(FE_OFN589_n_20904) );
in01f80 FE_OFC58_n_27012 ( .a(n_27012), .o(FE_OFN58_n_27012) );
in01f80 FE_OFC590_n_20904 ( .a(FE_OFN589_n_20904), .o(FE_OFN590_n_20904) );
in01f80 FE_OFC595_n_16896 ( .a(n_16896), .o(FE_OFN595_n_16896) );
in01f80 FE_OFC596_n_16896 ( .a(FE_OFN595_n_16896), .o(FE_OFN596_n_16896) );
in01f80 FE_OFC597_n_17615 ( .a(n_17615), .o(FE_OFN597_n_17615) );
in01f80 FE_OFC598_n_17615 ( .a(FE_OFN597_n_17615), .o(FE_OFN598_n_17615) );
in01f80 FE_OFC599_n_16000 ( .a(n_16000), .o(FE_OFN599_n_16000) );
in01f80 FE_OFC5_n_28597 ( .a(n_28597), .o(FE_OFN5_n_28597) );
in01f80 FE_OFC600_n_16000 ( .a(FE_OFN599_n_16000), .o(FE_OFN600_n_16000) );
in01f80 FE_OFC601_n_17761 ( .a(n_17761), .o(FE_OFN601_n_17761) );
in01f80 FE_OFC602_n_17761 ( .a(FE_OFN601_n_17761), .o(FE_OFN602_n_17761) );
in01f80 FE_OFC603_n_21535 ( .a(n_21535), .o(FE_OFN603_n_21535) );
in01f80 FE_OFC604_n_21535 ( .a(FE_OFN603_n_21535), .o(FE_OFN604_n_21535) );
in01f80 FE_OFC605_n_25225 ( .a(n_25225), .o(FE_OFN605_n_25225) );
in01f80 FE_OFC606_n_25225 ( .a(FE_OFN605_n_25225), .o(FE_OFN606_n_25225) );
in01f80 FE_OFC60_n_27012 ( .a(FE_OFN51_n_27012), .o(FE_OFN60_n_27012) );
in01f80 FE_OFC611_n_5698 ( .a(n_5698), .o(FE_OFN611_n_5698) );
in01f80 FE_OFC612_n_5698 ( .a(FE_OFN611_n_5698), .o(FE_OFN612_n_5698) );
in01f80 FE_OFC613_n_20110 ( .a(n_20110), .o(FE_OFN613_n_20110) );
in01f80 FE_OFC614_n_20110 ( .a(FE_OFN613_n_20110), .o(FE_OFN614_n_20110) );
in01f80 FE_OFC61_n_27012 ( .a(n_27012), .o(FE_OFN61_n_27012) );
in01f80 FE_OFC623_n_17378 ( .a(n_17378), .o(FE_OFN623_n_17378) );
in01f80 FE_OFC624_n_17378 ( .a(FE_OFN623_n_17378), .o(FE_OFN624_n_17378) );
in01f80 FE_OFC625_n_26697 ( .a(n_26697), .o(FE_OFN625_n_26697) );
in01f80 FE_OFC626_n_26697 ( .a(FE_OFN625_n_26697), .o(FE_OFN626_n_26697) );
in01f80 FE_OFC627_n_15605 ( .a(n_15605), .o(FE_OFN627_n_15605) );
in01f80 FE_OFC628_n_15605 ( .a(FE_OFN627_n_15605), .o(FE_OFN628_n_15605) );
in01f80 FE_OFC629_n_19358 ( .a(n_19358), .o(FE_OFN629_n_19358) );
in01f80 FE_OFC62_n_27012 ( .a(FE_OFN54_n_27012), .o(FE_OFN62_n_27012) );
in01f80 FE_OFC630_n_19358 ( .a(FE_OFN629_n_19358), .o(FE_OFN630_n_19358) );
in01f80 FE_OFC631_n_21154 ( .a(n_21154), .o(FE_OFN631_n_21154) );
in01f80 FE_OFC632_n_21154 ( .a(FE_OFN631_n_21154), .o(FE_OFN632_n_21154) );
in01f80 FE_OFC633_n_27731 ( .a(n_27731), .o(FE_OFN633_n_27731) );
in01f80 FE_OFC634_n_27731 ( .a(FE_OFN633_n_27731), .o(FE_OFN634_n_27731) );
in01f80 FE_OFC635_n_26260 ( .a(n_26260), .o(FE_OFN635_n_26260) );
in01f80 FE_OFC636_n_26260 ( .a(FE_OFN635_n_26260), .o(FE_OFN636_n_26260) );
in01f80 FE_OFC63_n_27012 ( .a(FE_OFN54_n_27012), .o(FE_OFN63_n_27012) );
in01f80 FE_OFC641_n_12432 ( .a(n_12432), .o(FE_OFN641_n_12432) );
in01f80 FE_OFC642_n_12432 ( .a(FE_OFN641_n_12432), .o(FE_OFN642_n_12432) );
in01f80 FE_OFC645_n_6732 ( .a(n_6732), .o(FE_OFN645_n_6732) );
in01f80 FE_OFC646_n_6732 ( .a(FE_OFN645_n_6732), .o(FE_OFN646_n_6732) );
in01f80 FE_OFC647_n_22008 ( .a(n_22008), .o(FE_OFN647_n_22008) );
in01f80 FE_OFC648_n_22008 ( .a(FE_OFN647_n_22008), .o(FE_OFN648_n_22008) );
in01f80 FE_OFC649_n_23576 ( .a(n_23576), .o(FE_OFN649_n_23576) );
in01f80 FE_OFC64_n_27012 ( .a(FE_OFN57_n_27012), .o(FE_OFN64_n_27012) );
in01f80 FE_OFC650_n_23576 ( .a(FE_OFN649_n_23576), .o(FE_OFN650_n_23576) );
in01f80 FE_OFC655_n_10503 ( .a(n_10503), .o(FE_OFN655_n_10503) );
in01f80 FE_OFC656_n_10503 ( .a(FE_OFN655_n_10503), .o(FE_OFN656_n_10503) );
in01f80 FE_OFC657_n_10424 ( .a(n_10424), .o(FE_OFN657_n_10424) );
in01f80 FE_OFC658_n_10424 ( .a(FE_OFN657_n_10424), .o(FE_OFN658_n_10424) );
in01f80 FE_OFC659_n_19445 ( .a(n_19445), .o(FE_OFN659_n_19445) );
in01f80 FE_OFC65_n_27012 ( .a(FE_OFN57_n_27012), .o(FE_OFN65_n_27012) );
in01f80 FE_OFC660_n_19445 ( .a(FE_OFN659_n_19445), .o(FE_OFN660_n_19445) );
in01f80 FE_OFC661_n_27899 ( .a(n_27899), .o(FE_OFN661_n_27899) );
in01f80 FE_OFC662_n_27899 ( .a(FE_OFN661_n_27899), .o(FE_OFN662_n_27899) );
in01f80 FE_OFC663_n_22027 ( .a(n_22027), .o(FE_OFN663_n_22027) );
in01f80 FE_OFC664_n_22027 ( .a(FE_OFN663_n_22027), .o(FE_OFN664_n_22027) );
in01f80 FE_OFC665_n_26759 ( .a(n_26759), .o(FE_OFN665_n_26759) );
in01f80 FE_OFC666_n_26759 ( .a(FE_OFN665_n_26759), .o(FE_OFN666_n_26759) );
in01f80 FE_OFC671_n_17494 ( .a(n_17494), .o(FE_OFN671_n_17494) );
in01f80 FE_OFC672_n_17494 ( .a(FE_OFN671_n_17494), .o(FE_OFN672_n_17494) );
in01f80 FE_OFC673_n_6720 ( .a(n_6720), .o(FE_OFN673_n_6720) );
in01f80 FE_OFC674_n_6720 ( .a(FE_OFN673_n_6720), .o(FE_OFN674_n_6720) );
in01f80 FE_OFC675_n_6824 ( .a(n_6824), .o(FE_OFN675_n_6824) );
in01f80 FE_OFC676_n_6824 ( .a(FE_OFN675_n_6824), .o(FE_OFN676_n_6824) );
in01f80 FE_OFC679_n_9691 ( .a(n_9691), .o(FE_OFN679_n_9691) );
in01f80 FE_OFC680_n_9691 ( .a(FE_OFN679_n_9691), .o(FE_OFN680_n_9691) );
in01f80 FE_OFC681_n_18155 ( .a(n_18155), .o(FE_OFN681_n_18155) );
in01f80 FE_OFC682_n_18155 ( .a(FE_OFN681_n_18155), .o(FE_OFN682_n_18155) );
in01f80 FE_OFC683_n_22025 ( .a(n_22025), .o(FE_OFN683_n_22025) );
in01f80 FE_OFC684_n_22025 ( .a(FE_OFN683_n_22025), .o(FE_OFN684_n_22025) );
in01f80 FE_OFC685_n_22968 ( .a(n_22968), .o(FE_OFN685_n_22968) );
in01f80 FE_OFC686_n_22968 ( .a(FE_OFN685_n_22968), .o(FE_OFN686_n_22968) );
in01f80 FE_OFC687_n_20109 ( .a(n_20109), .o(FE_OFN687_n_20109) );
in01f80 FE_OFC688_n_20109 ( .a(FE_OFN687_n_20109), .o(FE_OFN688_n_20109) );
in01f80 FE_OFC689_n_16216 ( .a(n_16216), .o(FE_OFN689_n_16216) );
in01f80 FE_OFC68_n_27012 ( .a(FE_OFN58_n_27012), .o(FE_OFN68_n_27012) );
in01f80 FE_OFC690_n_16216 ( .a(FE_OFN689_n_16216), .o(FE_OFN690_n_16216) );
in01f80 FE_OFC691_n_6708 ( .a(n_6708), .o(FE_OFN691_n_6708) );
in01f80 FE_OFC692_n_6708 ( .a(FE_OFN691_n_6708), .o(FE_OFN692_n_6708) );
in01f80 FE_OFC695_n_19853 ( .a(n_19853), .o(FE_OFN695_n_19853) );
in01f80 FE_OFC696_n_19853 ( .a(FE_OFN695_n_19853), .o(FE_OFN696_n_19853) );
in01f80 FE_OFC697_n_22333 ( .a(n_22333), .o(FE_OFN697_n_22333) );
in01f80 FE_OFC698_n_22333 ( .a(FE_OFN697_n_22333), .o(FE_OFN698_n_22333) );
in01f80 FE_OFC69_n_27012 ( .a(FE_OFN51_n_27012), .o(FE_OFN69_n_27012) );
in01f80 FE_OFC6_n_28597 ( .a(FE_OFN5_n_28597), .o(FE_OFN6_n_28597) );
in01f80 FE_OFC703_n_10462 ( .a(n_10462), .o(FE_OFN703_n_10462) );
in01f80 FE_OFC704_n_10462 ( .a(FE_OFN703_n_10462), .o(FE_OFN704_n_10462) );
in01f80 FE_OFC705_n_6444 ( .a(n_6444), .o(FE_OFN705_n_6444) );
in01f80 FE_OFC706_n_6444 ( .a(FE_OFN705_n_6444), .o(FE_OFN706_n_6444) );
in01f80 FE_OFC707_n_8059 ( .a(n_8059), .o(FE_OFN707_n_8059) );
in01f80 FE_OFC708_n_8059 ( .a(FE_OFN707_n_8059), .o(FE_OFN708_n_8059) );
in01f80 FE_OFC709_n_20192 ( .a(n_20192), .o(FE_OFN709_n_20192) );
in01f80 FE_OFC710_n_20192 ( .a(FE_OFN709_n_20192), .o(FE_OFN710_n_20192) );
in01f80 FE_OFC715_n_29187 ( .a(n_29187), .o(FE_OFN715_n_29187) );
in01f80 FE_OFC716_n_29187 ( .a(FE_OFN715_n_29187), .o(FE_OFN716_n_29187) );
in01f80 FE_OFC717_n_18993 ( .a(n_18993), .o(FE_OFN717_n_18993) );
in01f80 FE_OFC718_n_18993 ( .a(FE_OFN717_n_18993), .o(FE_OFN718_n_18993) );
in01f80 FE_OFC719_n_20807 ( .a(n_20807), .o(FE_OFN719_n_20807) );
in01f80 FE_OFC71_n_27012 ( .a(FE_OFN62_n_27012), .o(FE_OFN71_n_27012) );
in01f80 FE_OFC720_n_20807 ( .a(FE_OFN719_n_20807), .o(FE_OFN720_n_20807) );
in01f80 FE_OFC721_n_17438 ( .a(n_17438), .o(FE_OFN721_n_17438) );
in01f80 FE_OFC722_n_17438 ( .a(FE_OFN721_n_17438), .o(FE_OFN722_n_17438) );
in01f80 FE_OFC723_n_19019 ( .a(n_19019), .o(FE_OFN723_n_19019) );
in01f80 FE_OFC724_n_19019 ( .a(FE_OFN723_n_19019), .o(FE_OFN724_n_19019) );
in01f80 FE_OFC725_n_5240 ( .a(n_5240), .o(FE_OFN725_n_5240) );
in01f80 FE_OFC726_n_5240 ( .a(FE_OFN725_n_5240), .o(FE_OFN726_n_5240) );
in01f80 FE_OFC727_n_23636 ( .a(n_23636), .o(FE_OFN727_n_23636) );
in01f80 FE_OFC728_n_23636 ( .a(FE_OFN727_n_23636), .o(FE_OFN728_n_23636) );
in01f80 FE_OFC729_n_27888 ( .a(n_27888), .o(FE_OFN729_n_27888) );
in01f80 FE_OFC72_n_27012 ( .a(FE_OFN61_n_27012), .o(FE_OFN72_n_27012) );
in01f80 FE_OFC730_n_27888 ( .a(FE_OFN729_n_27888), .o(FE_OFN730_n_27888) );
in01f80 FE_OFC733_n_22952 ( .a(n_22952), .o(FE_OFN733_n_22952) );
in01f80 FE_OFC734_n_22952 ( .a(FE_OFN733_n_22952), .o(FE_OFN734_n_22952) );
in01f80 FE_OFC739_n_20195 ( .a(n_20195), .o(FE_OFN739_n_20195) );
in01f80 FE_OFC740_n_20195 ( .a(FE_OFN739_n_20195), .o(FE_OFN740_n_20195) );
in01f80 FE_OFC741_n_24025 ( .a(n_24025), .o(FE_OFN741_n_24025) );
in01f80 FE_OFC742_n_24025 ( .a(FE_OFN741_n_24025), .o(FE_OFN742_n_24025) );
in01f80 FE_OFC743_n_25732 ( .a(n_25732), .o(FE_OFN743_n_25732) );
in01f80 FE_OFC744_n_25732 ( .a(FE_OFN743_n_25732), .o(FE_OFN744_n_25732) );
in01f80 FE_OFC745_n_26604 ( .a(n_26604), .o(FE_OFN745_n_26604) );
in01f80 FE_OFC746_n_26604 ( .a(FE_OFN745_n_26604), .o(FE_OFN746_n_26604) );
in01f80 FE_OFC747_n_16529 ( .a(n_16529), .o(FE_OFN747_n_16529) );
in01f80 FE_OFC748_n_16529 ( .a(FE_OFN747_n_16529), .o(FE_OFN748_n_16529) );
in01f80 FE_OFC749_n_20252 ( .a(n_20252), .o(FE_OFN749_n_20252) );
in01f80 FE_OFC74_n_27012 ( .a(FE_OFN61_n_27012), .o(FE_OFN74_n_27012) );
in01f80 FE_OFC750_n_20252 ( .a(FE_OFN749_n_20252), .o(FE_OFN750_n_20252) );
in01f80 FE_OFC751_n_20252 ( .a(FE_OFN749_n_20252), .o(FE_OFN751_n_20252) );
in01f80 FE_OFC752_n_22913 ( .a(n_22913), .o(FE_OFN752_n_22913) );
in01f80 FE_OFC753_n_22913 ( .a(FE_OFN752_n_22913), .o(FE_OFN753_n_22913) );
in01f80 FE_OFC75_n_27012 ( .a(FE_OFN61_n_27012), .o(FE_OFN75_n_27012) );
in01f80 FE_OFC760_n_9661 ( .a(n_9661), .o(FE_OFN760_n_9661) );
in01f80 FE_OFC761_n_9661 ( .a(FE_OFN760_n_9661), .o(FE_OFN761_n_9661) );
in01f80 FE_OFC762_n_8501 ( .a(n_8501), .o(FE_OFN762_n_8501) );
in01f80 FE_OFC763_n_8501 ( .a(FE_OFN762_n_8501), .o(FE_OFN763_n_8501) );
in01f80 FE_OFC764_n_5707 ( .a(n_5707), .o(FE_OFN764_n_5707) );
in01f80 FE_OFC765_n_5707 ( .a(FE_OFN764_n_5707), .o(FE_OFN765_n_5707) );
in01f80 FE_OFC766_n_20476 ( .a(n_20476), .o(FE_OFN766_n_20476) );
in01f80 FE_OFC767_n_20476 ( .a(FE_OFN766_n_20476), .o(FE_OFN767_n_20476) );
in01f80 FE_OFC768_n_17379 ( .a(n_17379), .o(FE_OFN768_n_17379) );
in01f80 FE_OFC769_n_17379 ( .a(FE_OFN768_n_17379), .o(FE_OFN769_n_17379) );
in01f80 FE_OFC76_n_27012 ( .a(FE_OFN61_n_27012), .o(FE_OFN76_n_27012) );
in01f80 FE_OFC770_n_20323 ( .a(n_20323), .o(FE_OFN770_n_20323) );
in01f80 FE_OFC771_n_20323 ( .a(FE_OFN770_n_20323), .o(FE_OFN771_n_20323) );
in01f80 FE_OFC772_n_26698 ( .a(n_26698), .o(FE_OFN772_n_26698) );
in01f80 FE_OFC773_n_26698 ( .a(FE_OFN772_n_26698), .o(FE_OFN773_n_26698) );
in01f80 FE_OFC778_n_12158 ( .a(n_12158), .o(FE_OFN778_n_12158) );
in01f80 FE_OFC779_n_12158 ( .a(FE_OFN778_n_12158), .o(FE_OFN779_n_12158) );
in01f80 FE_OFC77_n_27012 ( .a(FE_OFN71_n_27012), .o(FE_OFN77_n_27012) );
in01f80 FE_OFC782_n_10771 ( .a(n_10771), .o(FE_OFN782_n_10771) );
in01f80 FE_OFC783_n_10771 ( .a(FE_OFN782_n_10771), .o(FE_OFN783_n_10771) );
in01f80 FE_OFC784_n_10198 ( .a(n_10198), .o(FE_OFN784_n_10198) );
in01f80 FE_OFC785_n_10198 ( .a(FE_OFN784_n_10198), .o(FE_OFN785_n_10198) );
in01f80 FE_OFC786_n_8855 ( .a(n_8855), .o(FE_OFN786_n_8855) );
in01f80 FE_OFC787_n_8855 ( .a(FE_OFN786_n_8855), .o(FE_OFN787_n_8855) );
in01f80 FE_OFC788_n_20913 ( .a(n_20913), .o(FE_OFN788_n_20913) );
in01f80 FE_OFC789_n_20913 ( .a(FE_OFN788_n_20913), .o(FE_OFN789_n_20913) );
in01f80 FE_OFC78_n_27012 ( .a(FE_OFN71_n_27012), .o(FE_OFN78_n_27012) );
in01f80 FE_OFC790_n_28272 ( .a(n_28272), .o(FE_OFN790_n_28272) );
in01f80 FE_OFC791_n_28272 ( .a(FE_OFN790_n_28272), .o(FE_OFN791_n_28272) );
in01f80 FE_OFC7_n_28597 ( .a(FE_OFN5_n_28597), .o(FE_OFN7_n_28597) );
in01f80 FE_OFC800_n_6782 ( .a(n_6782), .o(FE_OFN800_n_6782) );
in01f80 FE_OFC801_n_6782 ( .a(FE_OFN800_n_6782), .o(FE_OFN801_n_6782) );
in01f80 FE_OFC802_n_6771 ( .a(n_6771), .o(FE_OFN802_n_6771) );
in01f80 FE_OFC803_n_6771 ( .a(FE_OFN802_n_6771), .o(FE_OFN803_n_6771) );
in01f80 FE_OFC806_n_23617 ( .a(n_23617), .o(FE_OFN806_n_23617) );
in01f80 FE_OFC807_n_23617 ( .a(FE_OFN806_n_23617), .o(FE_OFN807_n_23617) );
in01f80 FE_OFC808_n_24927 ( .a(n_24927), .o(FE_OFN808_n_24927) );
in01f80 FE_OFC809_n_24927 ( .a(FE_OFN808_n_24927), .o(FE_OFN809_n_24927) );
in01f80 FE_OFC80_n_27012 ( .a(FE_OFN71_n_27012), .o(FE_OFN80_n_27012) );
in01f80 FE_OFC810_n_12878 ( .a(n_12878), .o(FE_OFN810_n_12878) );
in01f80 FE_OFC811_n_12878 ( .a(FE_OFN810_n_12878), .o(FE_OFN811_n_12878) );
in01f80 FE_OFC812_n_15982 ( .a(n_15982), .o(FE_OFN812_n_15982) );
in01f80 FE_OFC813_n_15982 ( .a(FE_OFN812_n_15982), .o(FE_OFN813_n_15982) );
in01f80 FE_OFC814_n_12310 ( .a(n_12310), .o(FE_OFN814_n_12310) );
in01f80 FE_OFC815_n_12310 ( .a(FE_OFN814_n_12310), .o(FE_OFN815_n_12310) );
in01f80 FE_OFC816_n_13135 ( .a(n_13135), .o(FE_OFN816_n_13135) );
in01f80 FE_OFC817_n_13135 ( .a(FE_OFN816_n_13135), .o(FE_OFN817_n_13135) );
in01f80 FE_OFC818_n_20821 ( .a(n_20821), .o(FE_OFN818_n_20821) );
in01f80 FE_OFC819_n_20821 ( .a(FE_OFN818_n_20821), .o(FE_OFN819_n_20821) );
in01f80 FE_OFC81_n_6529 ( .a(n_6529), .o(FE_OFN81_n_6529) );
in01f80 FE_OFC820_n_24644 ( .a(n_24644), .o(FE_OFN820_n_24644) );
in01f80 FE_OFC821_n_24644 ( .a(FE_OFN820_n_24644), .o(FE_OFN821_n_24644) );
in01f80 FE_OFC826_n_3772 ( .a(n_3772), .o(FE_OFN826_n_3772) );
in01f80 FE_OFC827_n_3772 ( .a(FE_OFN826_n_3772), .o(FE_OFN827_n_3772) );
in01f80 FE_OFC828_n_8424 ( .a(n_8424), .o(FE_OFN828_n_8424) );
in01f80 FE_OFC829_n_8424 ( .a(FE_OFN828_n_8424), .o(FE_OFN829_n_8424) );
in01f80 FE_OFC82_n_6529 ( .a(FE_OFN81_n_6529), .o(FE_OFN82_n_6529) );
in01f80 FE_OFC830_n_14863 ( .a(n_14863), .o(FE_OFN830_n_14863) );
in01f80 FE_OFC831_n_14863 ( .a(FE_OFN830_n_14863), .o(FE_OFN831_n_14863) );
in01f80 FE_OFC834_n_16760 ( .a(n_16760), .o(FE_OFN834_n_16760) );
in01f80 FE_OFC835_n_16760 ( .a(FE_OFN834_n_16760), .o(FE_OFN835_n_16760) );
in01f80 FE_OFC83_n_11673 ( .a(n_11673), .o(FE_OFN83_n_11673) );
in01f80 FE_OFC842_n_10412 ( .a(n_10412), .o(FE_OFN842_n_10412) );
in01f80 FE_OFC843_n_10412 ( .a(FE_OFN842_n_10412), .o(FE_OFN843_n_10412) );
in01f80 FE_OFC844_n_7616 ( .a(n_7616), .o(FE_OFN844_n_7616) );
in01f80 FE_OFC845_n_7616 ( .a(FE_OFN844_n_7616), .o(FE_OFN845_n_7616) );
in01f80 FE_OFC846_n_22340 ( .a(n_22340), .o(FE_OFN846_n_22340) );
in01f80 FE_OFC847_n_22340 ( .a(FE_OFN846_n_22340), .o(FE_OFN847_n_22340) );
in01f80 FE_OFC848_n_23567 ( .a(n_23567), .o(FE_OFN848_n_23567) );
in01f80 FE_OFC849_n_23567 ( .a(FE_OFN848_n_23567), .o(FE_OFN849_n_23567) );
in01f80 FE_OFC84_n_11673 ( .a(FE_OFN83_n_11673), .o(FE_OFN84_n_11673) );
in01f80 FE_OFC850_n_27728 ( .a(n_27728), .o(FE_OFN850_n_27728) );
in01f80 FE_OFC851_n_27728 ( .a(FE_OFN850_n_27728), .o(FE_OFN851_n_27728) );
in01f80 FE_OFC852_n_27880 ( .a(n_27880), .o(FE_OFN852_n_27880) );
in01f80 FE_OFC853_n_27880 ( .a(FE_OFN852_n_27880), .o(FE_OFN853_n_27880) );
in01f80 FE_OFC856_n_12565 ( .a(n_12565), .o(FE_OFN856_n_12565) );
in01f80 FE_OFC857_n_12565 ( .a(FE_OFN856_n_12565), .o(FE_OFN857_n_12565) );
in01f80 FE_OFC858_n_14125 ( .a(n_14125), .o(FE_OFN858_n_14125) );
in01f80 FE_OFC859_n_14125 ( .a(FE_OFN858_n_14125), .o(FE_OFN859_n_14125) );
in01f80 FE_OFC85_n_14586 ( .a(n_4860), .o(FE_OFN85_n_14586) );
in01f80 FE_OFC860_n_10492 ( .a(n_10492), .o(FE_OFN860_n_10492) );
in01f80 FE_OFC861_n_10492 ( .a(FE_OFN860_n_10492), .o(FE_OFN861_n_10492) );
in01f80 FE_OFC862_n_10495 ( .a(n_10495), .o(FE_OFN862_n_10495) );
in01f80 FE_OFC863_n_10495 ( .a(FE_OFN862_n_10495), .o(FE_OFN863_n_10495) );
in01f80 FE_OFC864_n_10501 ( .a(n_10501), .o(FE_OFN864_n_10501) );
in01f80 FE_OFC865_n_10501 ( .a(FE_OFN864_n_10501), .o(FE_OFN865_n_10501) );
in01f80 FE_OFC866_n_6151 ( .a(n_6151), .o(FE_OFN866_n_6151) );
in01f80 FE_OFC867_n_6151 ( .a(FE_OFN866_n_6151), .o(FE_OFN867_n_6151) );
in01f80 FE_OFC868_n_10506 ( .a(n_10506), .o(FE_OFN868_n_10506) );
in01f80 FE_OFC869_n_10506 ( .a(FE_OFN868_n_10506), .o(FE_OFN869_n_10506) );
in01f80 FE_OFC86_n_14586 ( .a(FE_OFN85_n_14586), .o(FE_OFN86_n_14586) );
in01f80 FE_OFC870_n_6154 ( .a(n_6154), .o(FE_OFN870_n_6154) );
in01f80 FE_OFC871_n_6154 ( .a(FE_OFN870_n_6154), .o(FE_OFN871_n_6154) );
in01f80 FE_OFC872_n_8070 ( .a(n_8070), .o(FE_OFN872_n_8070) );
in01f80 FE_OFC873_n_8070 ( .a(FE_OFN872_n_8070), .o(FE_OFN873_n_8070) );
in01f80 FE_OFC874_n_6157 ( .a(n_6157), .o(FE_OFN874_n_6157) );
in01f80 FE_OFC875_n_6157 ( .a(FE_OFN874_n_6157), .o(FE_OFN875_n_6157) );
in01f80 FE_OFC876_n_22329 ( .a(n_22329), .o(FE_OFN876_n_22329) );
in01f80 FE_OFC877_n_22329 ( .a(FE_OFN876_n_22329), .o(FE_OFN877_n_22329) );
in01f80 FE_OFC878_n_28229 ( .a(n_28229), .o(FE_OFN878_n_28229) );
in01f80 FE_OFC879_n_28229 ( .a(FE_OFN878_n_28229), .o(FE_OFN879_n_28229) );
in01f80 FE_OFC87_n_27449 ( .a(n_27449), .o(FE_OFN87_n_27449) );
in01f80 FE_OFC884_n_28405 ( .a(n_28405), .o(FE_OFN884_n_28405) );
in01f80 FE_OFC885_n_28405 ( .a(FE_OFN884_n_28405), .o(FE_OFN885_n_28405) );
in01f80 FE_OFC888_n_18291 ( .a(n_18291), .o(FE_OFN888_n_18291) );
in01f80 FE_OFC889_n_18291 ( .a(FE_OFN888_n_18291), .o(FE_OFN889_n_18291) );
in01f80 FE_OFC88_n_27449 ( .a(n_27449), .o(FE_OFN88_n_27449) );
in01f80 FE_OFC890_n_22165 ( .a(n_22165), .o(FE_OFN890_n_22165) );
in01f80 FE_OFC891_n_22165 ( .a(FE_OFN890_n_22165), .o(FE_OFN891_n_22165) );
in01f80 FE_OFC892_n_20806 ( .a(n_20806), .o(FE_OFN892_n_20806) );
in01f80 FE_OFC893_n_20806 ( .a(FE_OFN892_n_20806), .o(FE_OFN893_n_20806) );
in01f80 FE_OFC894_n_15923 ( .a(n_15923), .o(FE_OFN894_n_15923) );
in01f80 FE_OFC895_n_15923 ( .a(FE_OFN894_n_15923), .o(FE_OFN895_n_15923) );
in01f80 FE_OFC896_n_15930 ( .a(n_15930), .o(FE_OFN896_n_15930) );
in01f80 FE_OFC897_n_15930 ( .a(FE_OFN896_n_15930), .o(FE_OFN897_n_15930) );
in01f80 FE_OFC898_n_19332 ( .a(n_19332), .o(FE_OFN898_n_19332) );
in01f80 FE_OFC899_n_19332 ( .a(FE_OFN898_n_19332), .o(FE_OFN899_n_19332) );
in01f80 FE_OFC89_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN89_n_27449) );
in01f80 FE_OFC8_n_11667 ( .a(n_11667), .o(FE_OFN8_n_11667) );
in01f80 FE_OFC900_n_26098 ( .a(n_26098), .o(FE_OFN900_n_26098) );
in01f80 FE_OFC901_n_26098 ( .a(FE_OFN900_n_26098), .o(FE_OFN901_n_26098) );
in01f80 FE_OFC902_n_20903 ( .a(n_20903), .o(FE_OFN902_n_20903) );
in01f80 FE_OFC903_n_20903 ( .a(FE_OFN902_n_20903), .o(FE_OFN903_n_20903) );
in01f80 FE_OFC904_n_24967 ( .a(n_24967), .o(FE_OFN904_n_24967) );
in01f80 FE_OFC905_n_24967 ( .a(FE_OFN904_n_24967), .o(FE_OFN905_n_24967) );
in01f80 FE_OFC90_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN90_n_27449) );
in01f80 FE_OFC910_n_19850 ( .a(n_19850), .o(FE_OFN910_n_19850) );
in01f80 FE_OFC911_n_19850 ( .a(FE_OFN910_n_19850), .o(FE_OFN911_n_19850) );
in01f80 FE_OFC912_n_28409 ( .a(n_28409), .o(FE_OFN912_n_28409) );
in01f80 FE_OFC913_n_28409 ( .a(FE_OFN912_n_28409), .o(FE_OFN913_n_28409) );
in01f80 FE_OFC916_n_19297 ( .a(n_19297), .o(FE_OFN916_n_19297) );
in01f80 FE_OFC917_n_19297 ( .a(FE_OFN916_n_19297), .o(FE_OFN917_n_19297) );
in01f80 FE_OFC918_n_19575 ( .a(n_19575), .o(FE_OFN918_n_19575) );
in01f80 FE_OFC919_n_19575 ( .a(FE_OFN918_n_19575), .o(FE_OFN919_n_19575) );
in01f80 FE_OFC91_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN91_n_27449) );
in01f80 FE_OFC920_n_22498 ( .a(n_22498), .o(FE_OFN920_n_22498) );
in01f80 FE_OFC921_n_22498 ( .a(FE_OFN920_n_22498), .o(FE_OFN921_n_22498) );
in01f80 FE_OFC922_n_24430 ( .a(n_24430), .o(FE_OFN922_n_24430) );
in01f80 FE_OFC923_n_24430 ( .a(FE_OFN922_n_24430), .o(FE_OFN923_n_24430) );
in01f80 FE_OFC92_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN92_n_27449) );
in01f80 FE_OFC930_n_4898 ( .a(n_4898), .o(FE_OFN930_n_4898) );
in01f80 FE_OFC931_n_4898 ( .a(FE_OFN930_n_4898), .o(FE_OFN931_n_4898) );
in01f80 FE_OFC932_n_4950 ( .a(n_4950), .o(FE_OFN932_n_4950) );
in01f80 FE_OFC933_n_4950 ( .a(FE_OFN932_n_4950), .o(FE_OFN933_n_4950) );
in01f80 FE_OFC934_n_22317 ( .a(n_22317), .o(FE_OFN934_n_22317) );
in01f80 FE_OFC935_n_22317 ( .a(FE_OFN934_n_22317), .o(FE_OFN935_n_22317) );
in01f80 FE_OFC936_n_27359 ( .a(n_27359), .o(FE_OFN936_n_27359) );
in01f80 FE_OFC937_n_27359 ( .a(FE_OFN936_n_27359), .o(FE_OFN937_n_27359) );
in01f80 FE_OFC938_n_21084 ( .a(n_21084), .o(FE_OFN938_n_21084) );
in01f80 FE_OFC939_n_21084 ( .a(FE_OFN938_n_21084), .o(FE_OFN939_n_21084) );
in01f80 FE_OFC93_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN93_n_27449) );
in01f80 FE_OFC940_n_23815 ( .a(n_23815), .o(FE_OFN940_n_23815) );
in01f80 FE_OFC941_n_23815 ( .a(FE_OFN940_n_23815), .o(FE_OFN941_n_23815) );
in01f80 FE_OFC942_n_24127 ( .a(n_24127), .o(FE_OFN942_n_24127) );
in01f80 FE_OFC943_n_24127 ( .a(FE_OFN942_n_24127), .o(FE_OFN943_n_24127) );
in01f80 FE_OFC944_n_27398 ( .a(n_27398), .o(FE_OFN944_n_27398) );
in01f80 FE_OFC945_n_27398 ( .a(FE_OFN944_n_27398), .o(FE_OFN945_n_27398) );
in01f80 FE_OFC94_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN94_n_27449) );
in01f80 FE_OFC952_n_13421 ( .a(n_13421), .o(FE_OFN952_n_13421) );
in01f80 FE_OFC953_n_13421 ( .a(FE_OFN952_n_13421), .o(FE_OFN953_n_13421) );
in01f80 FE_OFC956_n_13438 ( .a(n_13438), .o(FE_OFN956_n_13438) );
in01f80 FE_OFC957_n_13438 ( .a(FE_OFN956_n_13438), .o(FE_OFN957_n_13438) );
in01f80 FE_OFC95_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN95_n_27449) );
in01f80 FE_OFC962_n_9280 ( .a(n_9280), .o(FE_OFN962_n_9280) );
in01f80 FE_OFC963_n_9280 ( .a(FE_OFN962_n_9280), .o(FE_OFN963_n_9280) );
in01f80 FE_OFC964_n_9283 ( .a(n_9283), .o(FE_OFN964_n_9283) );
in01f80 FE_OFC965_n_9283 ( .a(FE_OFN964_n_9283), .o(FE_OFN965_n_9283) );
in01f80 FE_OFC966_n_9286 ( .a(n_9286), .o(FE_OFN966_n_9286) );
in01f80 FE_OFC967_n_9286 ( .a(FE_OFN966_n_9286), .o(FE_OFN967_n_9286) );
in01f80 FE_OFC96_n_27449 ( .a(FE_OFN88_n_27449), .o(FE_OFN96_n_27449) );
in01f80 FE_OFC970_n_6854 ( .a(n_6854), .o(FE_OFN970_n_6854) );
in01f80 FE_OFC971_n_6854 ( .a(FE_OFN970_n_6854), .o(FE_OFN971_n_6854) );
in01f80 FE_OFC972_n_6822 ( .a(n_6822), .o(FE_OFN972_n_6822) );
in01f80 FE_OFC973_n_6822 ( .a(FE_OFN972_n_6822), .o(FE_OFN973_n_6822) );
in01f80 FE_OFC978_n_12566 ( .a(n_12566), .o(FE_OFN978_n_12566) );
in01f80 FE_OFC979_n_12566 ( .a(FE_OFN978_n_12566), .o(FE_OFN979_n_12566) );
in01f80 FE_OFC980_n_16353 ( .a(n_16353), .o(FE_OFN980_n_16353) );
in01f80 FE_OFC981_n_16353 ( .a(FE_OFN980_n_16353), .o(FE_OFN981_n_16353) );
in01f80 FE_OFC986_n_12804 ( .a(n_12804), .o(FE_OFN986_n_12804) );
in01f80 FE_OFC987_n_12804 ( .a(FE_OFN986_n_12804), .o(FE_OFN987_n_12804) );
in01f80 FE_OFC988_n_13374 ( .a(n_13374), .o(FE_OFN988_n_13374) );
in01f80 FE_OFC989_n_13374 ( .a(FE_OFN988_n_13374), .o(FE_OFN989_n_13374) );
in01f80 FE_OFC98_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN98_n_27449) );
in01f80 FE_OFC990_n_5720 ( .a(n_5720), .o(FE_OFN990_n_5720) );
in01f80 FE_OFC991_n_5720 ( .a(FE_OFN990_n_5720), .o(FE_OFN991_n_5720) );
in01f80 FE_OFC992_n_16934 ( .a(n_16934), .o(FE_OFN992_n_16934) );
in01f80 FE_OFC993_n_16934 ( .a(FE_OFN992_n_16934), .o(FE_OFN993_n_16934) );
in01f80 FE_OFC994_n_22325 ( .a(n_22325), .o(FE_OFN994_n_22325) );
in01f80 FE_OFC995_n_22325 ( .a(FE_OFN994_n_22325), .o(FE_OFN995_n_22325) );
in01f80 FE_OFC996_n_23622 ( .a(n_23622), .o(FE_OFN996_n_23622) );
in01f80 FE_OFC997_n_23622 ( .a(FE_OFN996_n_23622), .o(FE_OFN997_n_23622) );
in01f80 FE_OFC998_n_28782 ( .a(n_28782), .o(FE_OFN998_n_28782) );
in01f80 FE_OFC99_n_27449 ( .a(FE_OFN87_n_27449), .o(FE_OFN99_n_27449) );
in01f80 FE_OFC9_n_11667 ( .a(FE_OFN8_n_11667), .o(FE_OFN9_n_11667) );
in01f80 drc573191 ( .a(n_32744), .o(n_27231) );
oa12f80 g2 ( .a(n_8894), .b(n_32731), .c(n_13262), .o(n_32732) );
oa22f80 g539494 ( .a(n_29360), .b(FE_OFN295_n_3069), .c(n_638), .d(FE_OFN360_n_4860), .o(n_29580) );
oa22f80 g539495 ( .a(n_29271), .b(FE_OFN187_n_29496), .c(n_1950), .d(FE_OFN17_n_29617), .o(n_29497) );
oa22f80 g539496 ( .a(n_29593), .b(FE_OFN410_n_28303), .c(n_74), .d(FE_OFN130_n_27449), .o(n_29685) );
oa22f80 g539502 ( .a(n_29185), .b(FE_OFN295_n_3069), .c(n_47), .d(FE_OFN74_n_27012), .o(n_29415) );
oa22f80 g539503 ( .a(n_29594), .b(n_29683), .c(n_1138), .d(FE_OFN68_n_27012), .o(n_29669) );
oa22f80 g539504 ( .a(FE_OFN1126_n_29632), .b(n_29683), .c(n_1785), .d(FE_OFN349_n_4860), .o(n_29695) );
oa22f80 g539505 ( .a(n_29707), .b(FE_OFN402_n_28303), .c(n_1922), .d(FE_OFN1146_n_4860), .o(n_29710) );
ao12f80 g539519 ( .a(n_29193), .b(n_29192), .c(n_29191), .o(n_29360) );
ao12f80 g539520 ( .a(n_29128), .b(n_29127), .c(n_29135), .o(n_29271) );
ao12f80 g539521 ( .a(n_29469), .b(n_29468), .c(n_29467), .o(n_29593) );
oa22f80 g539522 ( .a(n_29673), .b(n_29698), .c(n_1103), .d(FE_OFN357_n_4860), .o(n_29706) );
oa22f80 g539523 ( .a(n_29633), .b(n_29698), .c(n_1817), .d(FE_OFN336_n_4860), .o(n_29699) );
oa22f80 g539524 ( .a(n_29526), .b(FE_OFN208_n_29661), .c(n_1945), .d(FE_OFN358_n_4860), .o(n_29662) );
oa22f80 g539525 ( .a(n_29653), .b(n_29664), .c(n_429), .d(FE_OFN347_n_4860), .o(n_29705) );
oa22f80 g539526 ( .a(n_29700), .b(FE_OFN211_n_29661), .c(n_1420), .d(FE_OFN100_n_27449), .o(n_29709) );
no02f80 g539547 ( .a(n_29192), .b(n_29191), .o(n_29193) );
no02f80 g539548 ( .a(n_29127), .b(n_29135), .o(n_29128) );
no02f80 g539549 ( .a(n_29468), .b(n_29467), .o(n_29469) );
ao12f80 g539550 ( .a(n_29064), .b(n_29063), .c(n_29062), .o(n_29185) );
ao12f80 g539551 ( .a(n_29536), .b(n_29535), .c(n_29534), .o(n_29632) );
ao12f80 g539552 ( .a(n_29703), .b(n_29702), .c(n_29701), .o(n_29707) );
ao12f80 g539553 ( .a(n_29473), .b(n_29472), .c(n_29471), .o(n_29594) );
oa22f80 g539554 ( .a(n_29609), .b(FE_OFN412_n_28303), .c(n_1132), .d(FE_OFN124_n_27449), .o(n_29672) );
oa22f80 g539555 ( .a(n_29607), .b(FE_OFN410_n_28303), .c(n_932), .d(FE_OFN350_n_4860), .o(n_29670) );
oa22f80 g539556 ( .a(n_29557), .b(n_29496), .c(n_855), .d(FE_OFN358_n_4860), .o(n_29651) );
oa22f80 g539557 ( .a(n_29605), .b(FE_OFN412_n_28303), .c(n_1815), .d(FE_OFN326_n_4860), .o(n_29667) );
oa22f80 g539558 ( .a(n_29604), .b(n_29683), .c(n_14), .d(FE_OFN68_n_27012), .o(n_29684) );
oa22f80 g539559 ( .a(n_29602), .b(n_29683), .c(n_838), .d(FE_OFN324_n_4860), .o(n_29681) );
oa22f80 g539560 ( .a(n_29494), .b(FE_OFN416_n_28303), .c(n_1901), .d(FE_OFN104_n_27449), .o(n_29649) );
oa22f80 g539561 ( .a(n_29367), .b(n_29698), .c(n_1935), .d(FE_OFN95_n_27449), .o(n_29584) );
oa22f80 g539562 ( .a(n_29491), .b(n_29698), .c(n_793), .d(FE_OFN95_n_27449), .o(n_29644) );
oa22f80 g539563 ( .a(FE_OFN1242_n_29553), .b(n_29691), .c(n_1776), .d(FE_OFN68_n_27012), .o(n_29656) );
oa22f80 g539564 ( .a(n_29694), .b(FE_OFN201_n_29637), .c(n_1030), .d(FE_OFN69_n_27012), .o(n_29708) );
oa22f80 g539565 ( .a(n_29490), .b(FE_OFN201_n_29637), .c(n_1788), .d(FE_OFN128_n_27449), .o(n_29638) );
oa22f80 g539566 ( .a(n_29432), .b(FE_OFN208_n_29661), .c(n_65), .d(FE_OFN122_n_27449), .o(n_29622) );
no02f80 g539597 ( .a(n_29535), .b(n_29534), .o(n_29536) );
no02f80 g539598 ( .a(n_29702), .b(n_29701), .o(n_29703) );
no02f80 g539599 ( .a(n_29472), .b(n_29471), .o(n_29473) );
no02f80 g539600 ( .a(n_29063), .b(n_29062), .o(n_29064) );
oa12f80 g539601 ( .a(n_28718), .b(n_28858), .c(n_29062), .o(n_29192) );
ao22s80 g539602 ( .a(n_29136), .b(n_28927), .c(n_29070), .d(x_in_52_14), .o(n_29468) );
ao12f80 g539603 ( .a(n_29636), .b(n_29635), .c(n_29634), .o(n_29673) );
ao12f80 g539604 ( .a(n_29564), .b(n_29563), .c(n_29562), .o(n_29633) );
oa22f80 g539605 ( .a(n_28487), .b(FE_OFN211_n_29661), .c(n_1292), .d(FE_OFN125_n_27449), .o(n_28763) );
ao12f80 g539606 ( .a(n_29450), .b(n_29449), .c(n_29448), .o(n_29526) );
ao12f80 g539607 ( .a(n_29614), .b(n_29613), .c(n_29612), .o(n_29653) );
ao12f80 g539608 ( .a(n_29677), .b(n_29676), .c(n_29675), .o(n_29700) );
ao12f80 g539609 ( .a(n_28796), .b(n_28927), .c(x_in_52_14), .o(n_29127) );
ao12f80 g539610 ( .a(n_28797), .b(n_28927), .c(x_in_52_15), .o(n_29467) );
oa22f80 g539611 ( .a(n_29579), .b(FE_OFN251_n_4162), .c(n_242), .d(FE_OFN119_n_27449), .o(n_29652) );
oa22f80 g539612 ( .a(n_29643), .b(n_29691), .c(n_1844), .d(FE_OFN1146_n_4860), .o(n_29693) );
oa22f80 g539613 ( .a(n_29642), .b(n_29691), .c(n_588), .d(FE_OFN336_n_4860), .o(n_29692) );
oa22f80 g539614 ( .a(n_29641), .b(n_29691), .c(n_741), .d(FE_OFN1123_rst), .o(n_29689) );
oa22f80 g539615 ( .a(n_29640), .b(n_29691), .c(n_808), .d(FE_OFN122_n_27449), .o(n_29686) );
oa22f80 g539616 ( .a(n_29627), .b(n_29691), .c(n_1925), .d(FE_OFN68_n_27012), .o(n_29668) );
oa22f80 g539617 ( .a(n_29626), .b(n_29664), .c(n_1368), .d(FE_OFN63_n_27012), .o(n_29665) );
oa22f80 g539618 ( .a(n_29639), .b(FE_OFN217_n_29687), .c(n_1053), .d(FE_OFN92_n_27449), .o(n_29696) );
oa22f80 g539619 ( .a(n_29505), .b(FE_OFN409_n_28303), .c(n_1923), .d(FE_OFN99_n_27449), .o(n_29650) );
oa22f80 g539620 ( .a(n_29625), .b(n_29687), .c(n_238), .d(FE_OFN99_n_27449), .o(n_29682) );
oa22f80 g539621 ( .a(n_29624), .b(n_29691), .c(n_17), .d(FE_OFN96_n_27449), .o(n_29680) );
oa22f80 g539622 ( .a(n_29623), .b(n_29691), .c(n_835), .d(n_27449), .o(n_29678) );
oa22f80 g539623 ( .a(n_29575), .b(n_29691), .c(n_697), .d(FE_OFN349_n_4860), .o(n_29660) );
oa22f80 g539624 ( .a(n_29503), .b(n_29664), .c(n_1018), .d(FE_OFN56_n_27012), .o(n_29647) );
oa22f80 g539625 ( .a(n_29384), .b(n_29664), .c(n_164), .d(FE_OFN63_n_27012), .o(n_29583) );
oa22f80 g539626 ( .a(n_29501), .b(FE_OFN269_n_4280), .c(n_502), .d(FE_OFN1143_n_27012), .o(n_29646) );
oa22f80 g539627 ( .a(n_29216), .b(n_22019), .c(n_426), .d(FE_OFN63_n_27012), .o(n_29454) );
oa22f80 g539628 ( .a(n_29574), .b(FE_OFN268_n_4280), .c(n_664), .d(FE_OFN329_n_4860), .o(n_29657) );
oa22f80 g539629 ( .a(n_28392), .b(n_28486), .c(n_306), .d(FE_OFN72_n_27012), .o(n_28716) );
no02f80 g539658 ( .a(n_29635), .b(n_29634), .o(n_29636) );
no02f80 g539659 ( .a(n_29563), .b(n_29562), .o(n_29564) );
no02f80 g539660 ( .a(n_29449), .b(n_29448), .o(n_29450) );
no02f80 g539661 ( .a(n_28927), .b(x_in_52_15), .o(n_28797) );
na03f80 g539662 ( .a(n_28477), .b(n_28355), .c(n_4340), .o(n_28708) );
no02f80 g539663 ( .a(n_29613), .b(n_29612), .o(n_29614) );
no02f80 g539664 ( .a(n_28719), .b(n_28858), .o(n_29063) );
no02f80 g539665 ( .a(n_28927), .b(x_in_52_14), .o(n_28796) );
no02f80 g539666 ( .a(n_29676), .b(n_29675), .o(n_29677) );
oa12f80 g539667 ( .a(n_28389), .b(n_29438), .c(n_28599), .o(n_29535) );
oa12f80 g539668 ( .a(n_28181), .b(n_29674), .c(n_28360), .o(n_29702) );
oa12f80 g539669 ( .a(n_27867), .b(n_29369), .c(n_28177), .o(n_29472) );
ao12f80 g539670 ( .a(n_29508), .b(n_29507), .c(n_29581), .o(n_29609) );
ao12f80 g539671 ( .a(n_29521), .b(n_29520), .c(n_29519), .o(n_29607) );
ao12f80 g539672 ( .a(n_29460), .b(n_29562), .c(n_29459), .o(n_29557) );
ao12f80 g539673 ( .a(n_29518), .b(n_29517), .c(n_29516), .o(n_29605) );
ao12f80 g539674 ( .a(n_29514), .b(n_29513), .c(n_29512), .o(n_29604) );
ao12f80 g539675 ( .a(n_29511), .b(n_29510), .c(n_29509), .o(n_29602) );
ao12f80 g539676 ( .a(n_29393), .b(n_29392), .c(n_29455), .o(n_29494) );
oa12f80 g539677 ( .a(n_28636), .b(n_28644), .c(x_in_52_15), .o(n_29191) );
ao12f80 g539678 ( .a(n_29243), .b(n_29242), .c(n_29333), .o(n_29367) );
ao12f80 g539679 ( .a(n_29389), .b(n_29388), .c(n_29438), .o(n_29491) );
ao12f80 g539680 ( .a(n_29458), .b(n_29457), .c(n_29456), .o(n_29553) );
ao12f80 g539681 ( .a(n_29391), .b(n_29489), .c(n_29390), .o(n_29490) );
ao12f80 g539682 ( .a(n_29659), .b(n_29674), .c(n_29658), .o(n_29694) );
ao12f80 g539683 ( .a(n_29335), .b(n_29369), .c(n_29334), .o(n_29432) );
oa22f80 g539684 ( .a(n_29359), .b(FE_OFN300_n_3069), .c(n_1470), .d(FE_OFN91_n_27449), .o(n_29540) );
oa22f80 g539685 ( .a(n_29420), .b(FE_OFN309_n_3069), .c(n_1451), .d(FE_OFN134_n_27449), .o(n_29601) );
oa22f80 g539686 ( .a(n_29419), .b(FE_OFN313_n_3069), .c(n_1625), .d(FE_OFN361_n_4860), .o(n_29600) );
oa22f80 g539687 ( .a(n_29418), .b(FE_OFN313_n_3069), .c(n_568), .d(FE_OFN1174_n_4860), .o(n_29598) );
oa22f80 g539688 ( .a(n_29358), .b(n_22019), .c(n_828), .d(FE_OFN1115_rst), .o(n_29533) );
oa22f80 g539689 ( .a(n_29417), .b(n_22019), .c(n_909), .d(FE_OFN1117_rst), .o(n_29596) );
oa22f80 g539690 ( .a(n_29357), .b(FE_OFN299_n_3069), .c(n_880), .d(FE_OFN350_n_4860), .o(n_29532) );
oa22f80 g539691 ( .a(n_29356), .b(FE_OFN267_n_4280), .c(n_1019), .d(FE_OFN326_n_4860), .o(n_29530) );
oa22f80 g539692 ( .a(n_29274), .b(FE_OFN258_n_4280), .c(n_1325), .d(FE_OFN77_n_27012), .o(n_29470) );
oa22f80 g539693 ( .a(n_29355), .b(n_4280), .c(n_1041), .d(FE_OFN78_n_27012), .o(n_29528) );
oa22f80 g539694 ( .a(FE_OFN1264_n_29354), .b(n_22019), .c(n_335), .d(FE_OFN1171_n_4860), .o(n_29525) );
oa22f80 g539695 ( .a(n_29182), .b(FE_OFN296_n_3069), .c(n_1444), .d(FE_OFN352_n_4860), .o(n_29416) );
oa22f80 g539696 ( .a(n_29466), .b(FE_OFN294_n_3069), .c(n_1506), .d(FE_OFN1109_rst), .o(n_29631) );
oa22f80 g539697 ( .a(n_28434), .b(FE_OFN259_n_4280), .c(n_1517), .d(FE_OFN130_n_27449), .o(n_28759) );
oa22f80 g539698 ( .a(n_29111), .b(n_23291), .c(n_1637), .d(FE_OFN1117_rst), .o(n_29353) );
oa22f80 g539699 ( .a(n_29273), .b(FE_OFN253_n_4280), .c(n_480), .d(FE_OFN1121_rst), .o(n_29465) );
oa22f80 g539700 ( .a(n_29272), .b(FE_OFN297_n_3069), .c(n_340), .d(FE_OFN352_n_4860), .o(n_29464) );
oa22f80 g539701 ( .a(n_29181), .b(FE_OFN300_n_3069), .c(n_296), .d(FE_OFN60_n_27012), .o(n_29410) );
oa22f80 g539702 ( .a(n_29110), .b(FE_OFN259_n_4280), .c(n_1165), .d(FE_OFN108_n_27449), .o(n_29350) );
oa22f80 g539703 ( .a(n_29413), .b(FE_OFN310_n_3069), .c(n_1326), .d(FE_OFN134_n_27449), .o(n_29592) );
oa22f80 g539704 ( .a(n_29412), .b(FE_OFN299_n_3069), .c(n_24), .d(FE_OFN74_n_27012), .o(n_29589) );
oa22f80 g539705 ( .a(n_29351), .b(FE_OFN297_n_3069), .c(n_277), .d(FE_OFN78_n_27012), .o(n_29524) );
oa22f80 g539706 ( .a(n_29411), .b(FE_OFN300_n_3069), .c(n_486), .d(FE_OFN91_n_27449), .o(n_29588) );
oa22f80 g539707 ( .a(n_29515), .b(FE_OFN214_n_29687), .c(n_1348), .d(FE_OFN363_n_4860), .o(n_29629) );
oa22f80 g539708 ( .a(n_29630), .b(FE_OFN214_n_29687), .c(n_1256), .d(FE_OFN1109_rst), .o(n_29688) );
oa22f80 g539709 ( .a(n_29409), .b(n_4280), .c(n_1563), .d(FE_OFN1109_rst), .o(n_29587) );
oa22f80 g539710 ( .a(n_29040), .b(FE_OFN259_n_4280), .c(n_1755), .d(FE_OFN130_n_27449), .o(n_29256) );
oa22f80 g539711 ( .a(n_29421), .b(FE_OFN314_n_3069), .c(n_1867), .d(FE_OFN12_n_29204), .o(n_29585) );
oa22f80 g539712 ( .a(n_28105), .b(n_28644), .c(n_1612), .d(FE_OFN100_n_27449), .o(n_28645) );
no02f80 g539762 ( .a(n_29520), .b(n_29519), .o(n_29521) );
no02f80 g539763 ( .a(n_29517), .b(n_29516), .o(n_29518) );
no02f80 g539764 ( .a(n_29562), .b(n_29459), .o(n_29460) );
no02f80 g539765 ( .a(n_29513), .b(n_29512), .o(n_29514) );
no02f80 g539766 ( .a(n_29510), .b(n_29509), .o(n_29511) );
no02f80 g539767 ( .a(n_29392), .b(n_29455), .o(n_29393) );
na02f80 g539768 ( .a(n_28644), .b(x_in_52_15), .o(n_28636) );
no02f80 g539769 ( .a(n_29457), .b(n_29456), .o(n_29458) );
no02f80 g539770 ( .a(n_29489), .b(n_29390), .o(n_29391) );
no02f80 g539771 ( .a(n_29369), .b(n_29334), .o(n_29335) );
in01f80 g539772 ( .a(n_28718), .o(n_28719) );
na02f80 g539773 ( .a(n_28644), .b(x_in_52_14), .o(n_28718) );
no02f80 g539774 ( .a(n_28644), .b(x_in_52_14), .o(n_28858) );
no02f80 g539775 ( .a(n_29507), .b(n_29581), .o(n_29508) );
no02f80 g539776 ( .a(n_29242), .b(n_29333), .o(n_29243) );
no02f80 g539777 ( .a(n_29388), .b(n_29438), .o(n_29389) );
oa12f80 g539778 ( .a(n_28393), .b(n_29581), .c(n_28603), .o(n_29635) );
oa12f80 g539779 ( .a(n_28198), .b(n_29333), .c(n_28361), .o(n_29449) );
no02f80 g539780 ( .a(n_29674), .b(n_29658), .o(n_29659) );
ao12f80 g539781 ( .a(n_28357), .b(n_28482), .c(n_29455), .o(n_29563) );
oa12f80 g539782 ( .a(n_28401), .b(n_27994), .c(n_28400), .o(n_28635) );
oa12f80 g539783 ( .a(n_28258), .b(n_28260), .c(n_28104), .o(n_28511) );
ao22s80 g539784 ( .a(n_29072), .b(x_in_36_14), .c(n_29506), .d(n_27456), .o(n_29676) );
oa12f80 g539785 ( .a(n_27996), .b(n_29502), .c(n_27800), .o(n_29613) );
oa12f80 g539786 ( .a(rst), .b(n_28354), .c(n_28391), .o(n_28392) );
ao12f80 g539787 ( .a(n_29552), .b(n_29551), .c(n_29550), .o(n_29643) );
ao12f80 g539788 ( .a(n_29549), .b(n_29548), .c(n_29547), .o(n_29642) );
ao12f80 g539789 ( .a(n_29546), .b(n_29545), .c(n_29544), .o(n_29641) );
ao12f80 g539790 ( .a(n_29543), .b(n_29542), .c(n_29541), .o(n_29640) );
ao12f80 g539791 ( .a(n_29431), .b(n_29430), .c(n_29429), .o(n_29579) );
ao12f80 g539792 ( .a(n_29488), .b(n_29487), .c(n_29486), .o(n_29627) );
ao12f80 g539793 ( .a(n_29485), .b(n_29484), .c(n_29483), .o(n_29626) );
ao12f80 g539794 ( .a(n_29539), .b(n_29538), .c(n_29537), .o(n_29639) );
ao12f80 g539795 ( .a(n_29366), .b(n_29365), .c(n_29364), .o(n_29505) );
ao12f80 g539796 ( .a(n_29482), .b(n_29481), .c(n_29480), .o(n_29625) );
ao12f80 g539797 ( .a(n_29479), .b(n_29478), .c(n_29477), .o(n_29624) );
ao12f80 g539798 ( .a(n_29476), .b(n_29475), .c(n_29474), .o(n_29623) );
ao12f80 g539799 ( .a(n_29428), .b(n_29427), .c(n_29426), .o(n_29575) );
ao22s80 g539800 ( .a(n_29502), .b(n_28111), .c(n_29313), .d(n_28110), .o(n_29503) );
ao12f80 g539801 ( .a(n_29189), .b(n_29188), .c(FE_OFN716_n_29187), .o(n_29384) );
ao12f80 g539802 ( .a(n_28644), .b(n_26577), .c(n_26926), .o(n_28927) );
ao12f80 g539803 ( .a(n_29363), .b(n_29362), .c(n_29361), .o(n_29501) );
ao12f80 g539804 ( .a(n_29066), .b(n_29129), .c(n_29065), .o(n_29216) );
ao12f80 g539805 ( .a(n_29424), .b(n_29423), .c(n_29422), .o(n_29574) );
oa22f80 g539806 ( .a(n_29312), .b(n_29664), .c(n_704), .d(FE_OFN347_n_4860), .o(n_29500) );
oa22f80 g539807 ( .a(n_29382), .b(n_29664), .c(n_1463), .d(n_27709), .o(n_29573) );
oa22f80 g539808 ( .a(n_29380), .b(FE_OFN416_n_28303), .c(n_1134), .d(FE_OFN1117_rst), .o(n_29572) );
oa22f80 g539809 ( .a(n_29452), .b(n_29687), .c(n_1648), .d(n_29068), .o(n_29620) );
oa22f80 g539810 ( .a(n_29444), .b(FE_OFN217_n_29687), .c(n_1831), .d(n_29617), .o(n_29619) );
oa22f80 g539811 ( .a(n_29447), .b(FE_OFN294_n_3069), .c(n_672), .d(FE_OFN17_n_29617), .o(n_29618) );
oa22f80 g539812 ( .a(n_29215), .b(n_27681), .c(n_1889), .d(FE_OFN1112_rst), .o(n_29446) );
oa22f80 g539813 ( .a(n_29378), .b(FE_OFN307_n_3069), .c(n_1469), .d(FE_OFN1106_rst), .o(n_29570) );
oa22f80 g539814 ( .a(n_29376), .b(n_22019), .c(n_1230), .d(FE_OFN1117_rst), .o(n_29569) );
oa22f80 g539815 ( .a(n_29374), .b(FE_OFN293_n_3069), .c(n_8), .d(FE_OFN1109_rst), .o(n_29566) );
oa22f80 g539816 ( .a(n_29443), .b(FE_OFN297_n_3069), .c(n_1775), .d(FE_OFN104_n_27449), .o(n_29616) );
oa22f80 g539817 ( .a(n_28476), .b(FE_OFN306_n_3069), .c(n_536), .d(FE_OFN125_n_27449), .o(n_28494) );
oa22f80 g539818 ( .a(n_29311), .b(n_22019), .c(n_1133), .d(FE_OFN347_n_4860), .o(n_29498) );
oa22f80 g539819 ( .a(FE_OFN1128_n_29567), .b(n_29664), .c(n_1571), .d(FE_OFN1108_rst), .o(n_29654) );
oa22f80 g539820 ( .a(n_29442), .b(FE_OFN307_n_3069), .c(n_55), .d(FE_OFN1106_rst), .o(n_29611) );
oa22f80 g539821 ( .a(n_29372), .b(FE_OFN294_n_3069), .c(n_1746), .d(FE_OFN138_n_27449), .o(n_29561) );
oa22f80 g539822 ( .a(n_29441), .b(FE_OFN217_n_29687), .c(n_675), .d(FE_OFN96_n_27449), .o(n_29608) );
oa22f80 g539823 ( .a(n_29371), .b(FE_OFN214_n_29687), .c(n_749), .d(FE_OFN131_n_27449), .o(n_29559) );
oa22f80 g539824 ( .a(n_29440), .b(FE_OFN236_n_4162), .c(n_273), .d(FE_OFN64_n_27012), .o(n_29606) );
oa22f80 g539825 ( .a(n_29310), .b(FE_OFN414_n_28303), .c(n_1898), .d(FE_OFN116_n_27449), .o(n_29495) );
oa22f80 g539826 ( .a(n_29439), .b(FE_OFN414_n_28303), .c(n_1546), .d(FE_OFN116_n_27449), .o(n_29603) );
oa22f80 g539827 ( .a(n_29370), .b(FE_OFN412_n_28303), .c(n_341), .d(FE_OFN124_n_27449), .o(n_29556) );
oa22f80 g539828 ( .a(n_29071), .b(FE_OFN186_n_29496), .c(n_1161), .d(FE_OFN125_n_27449), .o(n_29300) );
oa22f80 g539829 ( .a(n_29213), .b(FE_OFN414_n_28303), .c(n_1350), .d(FE_OFN116_n_27449), .o(n_29437) );
oa22f80 g539830 ( .a(n_29309), .b(FE_OFN312_n_3069), .c(n_449), .d(FE_OFN124_n_27449), .o(n_29493) );
oa22f80 g539831 ( .a(n_29307), .b(FE_OFN166_n_29269), .c(n_1693), .d(FE_OFN108_n_27449), .o(n_29492) );
in01f80 g539832 ( .a(n_28486), .o(n_28487) );
oa22f80 g539833 ( .a(n_28021), .b(n_21777), .c(n_3364), .d(x_in_25_15), .o(n_28486) );
no02f80 g539850 ( .a(n_28394), .b(n_28603), .o(n_29507) );
no02f80 g539851 ( .a(n_29551), .b(n_29550), .o(n_29552) );
no02f80 g539852 ( .a(n_29548), .b(n_29547), .o(n_29549) );
no02f80 g539853 ( .a(n_29545), .b(n_29544), .o(n_29546) );
no02f80 g539854 ( .a(n_29542), .b(n_29541), .o(n_29543) );
no02f80 g539855 ( .a(n_29430), .b(n_29429), .o(n_29431) );
na02f80 g539856 ( .a(n_28356), .b(n_28482), .o(n_29392) );
no02f80 g539857 ( .a(n_29487), .b(n_29486), .o(n_29488) );
no02f80 g539858 ( .a(n_29484), .b(n_29483), .o(n_29485) );
no02f80 g539859 ( .a(n_29538), .b(n_29537), .o(n_29539) );
no02f80 g539860 ( .a(n_29365), .b(n_29364), .o(n_29366) );
no02f80 g539861 ( .a(n_29481), .b(n_29480), .o(n_29482) );
no02f80 g539862 ( .a(n_29478), .b(n_29477), .o(n_29479) );
no02f80 g539863 ( .a(n_29475), .b(n_29474), .o(n_29476) );
no02f80 g539864 ( .a(n_28199), .b(n_28361), .o(n_29242) );
no02f80 g539865 ( .a(n_29427), .b(n_29426), .o(n_29428) );
no02f80 g539866 ( .a(n_28390), .b(n_28599), .o(n_29388) );
no02f80 g539867 ( .a(n_29188), .b(FE_OFN716_n_29187), .o(n_29189) );
na02f80 g539868 ( .a(n_29135), .b(n_616), .o(n_29136) );
no02f80 g539869 ( .a(n_29129), .b(n_29065), .o(n_29066) );
no02f80 g539870 ( .a(n_29423), .b(n_29422), .o(n_29424) );
no02f80 g539871 ( .a(n_28360), .b(n_28182), .o(n_29658) );
no02f80 g539872 ( .a(n_29362), .b(n_29361), .o(n_29363) );
oa12f80 g539873 ( .a(n_28092), .b(n_29276), .c(n_28266), .o(n_29457) );
oa12f80 g539874 ( .a(n_28356), .b(n_27821), .c(n_27857), .o(n_28357) );
oa12f80 g539875 ( .a(n_28260), .b(n_80), .c(FE_OFN100_n_27449), .o(n_28261) );
ao22s80 g539876 ( .a(n_27861), .b(n_27675), .c(x_out_43_32), .d(n_27400), .o(n_28258) );
ao12f80 g539877 ( .a(n_27705), .b(n_29129), .c(n_28047), .o(n_29369) );
ao12f80 g539878 ( .a(n_29504), .b(n_29489), .c(x_in_20_13), .o(n_29674) );
ao12f80 g539879 ( .a(n_28225), .b(n_28264), .c(n_29186), .o(n_29438) );
na03f80 g539880 ( .a(n_27993), .b(n_28354), .c(n_28400), .o(n_28355) );
na03f80 g539881 ( .a(n_28391), .b(n_28476), .c(rst), .o(n_28477) );
oa12f80 g539882 ( .a(FE_OFN1109_rst), .b(n_28039), .c(n_28104), .o(n_28105) );
ao12f80 g539883 ( .a(n_29331), .b(n_29330), .c(n_29383), .o(n_29421) );
ao12f80 g539884 ( .a(n_28169), .b(n_28168), .c(n_29429), .o(n_29634) );
ao12f80 g539885 ( .a(n_29235), .b(n_29234), .c(n_29233), .o(n_29359) );
ao12f80 g539886 ( .a(n_29329), .b(n_29328), .c(n_29327), .o(n_29420) );
ao12f80 g539887 ( .a(n_29326), .b(n_29325), .c(n_29324), .o(n_29419) );
ao12f80 g539888 ( .a(n_29232), .b(n_29231), .c(FE_OFN1268_n_29314), .o(n_29358) );
ao12f80 g539889 ( .a(n_29323), .b(n_29322), .c(n_29321), .o(n_29418) );
ao12f80 g539890 ( .a(n_29320), .b(n_29319), .c(n_29318), .o(n_29417) );
ao12f80 g539891 ( .a(n_29230), .b(n_29229), .c(n_29228), .o(n_29357) );
ao12f80 g539892 ( .a(n_28037), .b(n_28254), .c(n_28036), .o(n_29520) );
ao12f80 g539893 ( .a(n_29157), .b(n_29156), .c(n_29155), .o(n_29274) );
ao12f80 g539894 ( .a(n_29227), .b(n_29226), .c(n_29225), .o(n_29356) );
ao12f80 g539895 ( .a(n_28035), .b(n_28247), .c(n_28034), .o(n_29517) );
oa12f80 g539896 ( .a(n_28290), .b(n_28289), .c(x_in_6_15), .o(n_29562) );
ao12f80 g539897 ( .a(n_28033), .b(n_28246), .c(n_28032), .o(n_29513) );
ao12f80 g539898 ( .a(n_29224), .b(n_29223), .c(n_29222), .o(n_29355) );
ao12f80 g539899 ( .a(n_29221), .b(n_29220), .c(n_29219), .o(n_29354) );
ao12f80 g539900 ( .a(n_28031), .b(n_29234), .c(n_28030), .o(n_29510) );
ao12f80 g539901 ( .a(n_29087), .b(n_29086), .c(n_29085), .o(n_29182) );
in01f80 g539902 ( .a(n_28644), .o(n_28434) );
na02f80 g539903 ( .a(n_28046), .b(n_28173), .o(n_28644) );
ao12f80 g539904 ( .a(n_29387), .b(n_29386), .c(n_29385), .o(n_29466) );
ao12f80 g539905 ( .a(n_28960), .b(n_28959), .c(n_29074), .o(n_29111) );
ao12f80 g539906 ( .a(n_29154), .b(n_29153), .c(n_29152), .o(n_29273) );
ao12f80 g539907 ( .a(n_29151), .b(n_29150), .c(n_29186), .o(n_29272) );
ao12f80 g539908 ( .a(n_29083), .b(n_29082), .c(n_29081), .o(n_29181) );
ao12f80 g539909 ( .a(n_28955), .b(n_28954), .c(n_29075), .o(n_29110) );
ao12f80 g539910 ( .a(n_29317), .b(n_29316), .c(n_29315), .o(n_29413) );
ao22s80 g539911 ( .a(n_28254), .b(n_29241), .c(n_27851), .d(n_29240), .o(n_29412) );
ao12f80 g539912 ( .a(n_29218), .b(n_29217), .c(n_29276), .o(n_29351) );
ao22s80 g539913 ( .a(n_28247), .b(n_29239), .c(n_27842), .d(n_29238), .o(n_29411) );
ao12f80 g539914 ( .a(n_29578), .b(n_29577), .c(n_29576), .o(n_29630) );
oa12f80 g539915 ( .a(n_28060), .b(n_28221), .c(x_in_20_15), .o(n_29701) );
ao12f80 g539916 ( .a(n_28873), .b(n_28939), .c(n_28872), .o(n_29040) );
ao22s80 g539917 ( .a(n_28246), .b(n_29237), .c(n_27835), .d(n_29236), .o(n_29409) );
oa22f80 g539918 ( .a(n_29067), .b(FE_OFN166_n_29269), .c(n_757), .d(FE_OFN91_n_27449), .o(n_29270) );
oa22f80 g539919 ( .a(n_29134), .b(FE_OFN265_n_4280), .c(n_22), .d(FE_OFN1181_rst), .o(n_29349) );
oa22f80 g539920 ( .a(n_29133), .b(FE_OFN264_n_4280), .c(n_739), .d(n_29104), .o(n_29347) );
oa22f80 g539921 ( .a(n_29132), .b(FE_OFN254_n_4280), .c(n_1137), .d(FE_OFN361_n_4860), .o(n_29346) );
oa22f80 g539922 ( .a(n_29131), .b(FE_OFN313_n_3069), .c(n_203), .d(FE_OFN1174_n_4860), .o(n_29344) );
oa22f80 g539923 ( .a(n_29130), .b(FE_OFN308_n_3069), .c(n_1560), .d(FE_OFN287_n_29266), .o(n_29343) );
oa22f80 g539924 ( .a(n_29061), .b(FE_OFN299_n_3069), .c(n_1093), .d(FE_OFN286_n_29266), .o(n_29268) );
oa22f80 g539925 ( .a(n_28937), .b(FE_OFN257_n_4280), .c(n_1951), .d(n_29261), .o(n_29178) );
oa22f80 g539926 ( .a(n_29060), .b(FE_OFN308_n_3069), .c(n_460), .d(n_29264), .o(n_29265) );
oa22f80 g539927 ( .a(n_29059), .b(FE_OFN230_n_4162), .c(n_1178), .d(n_29261), .o(n_29263) );
oa22f80 g539928 ( .a(n_29058), .b(FE_OFN248_n_4162), .c(n_1944), .d(FE_OFN91_n_27449), .o(n_29260) );
oa22f80 g539929 ( .a(n_28847), .b(n_29683), .c(n_62), .d(FE_OFN95_n_27449), .o(n_29108) );
oa22f80 g539930 ( .a(n_29057), .b(FE_OFN234_n_4162), .c(n_1320), .d(FE_OFN133_n_27449), .o(n_29258) );
oa22f80 g539931 ( .a(n_29056), .b(n_16028), .c(n_488), .d(n_25680), .o(n_29257) );
oa22f80 g539932 ( .a(n_29126), .b(FE_OFN184_n_29402), .c(n_1078), .d(n_29261), .o(n_29342) );
oa22f80 g539933 ( .a(n_29125), .b(FE_OFN234_n_4162), .c(n_942), .d(FE_OFN363_n_4860), .o(n_29341) );
oa22f80 g539934 ( .a(n_28846), .b(FE_OFN236_n_4162), .c(n_1496), .d(FE_OFN357_n_4860), .o(n_29103) );
oa22f80 g539935 ( .a(n_29124), .b(n_4162), .c(n_489), .d(FE_OFN1181_rst), .o(n_29340) );
oa22f80 g539936 ( .a(n_29055), .b(FE_OFN236_n_4162), .c(n_1265), .d(FE_OFN1106_rst), .o(n_29254) );
oa22f80 g539937 ( .a(n_29054), .b(FE_OFN184_n_29402), .c(n_1279), .d(n_27449), .o(n_29253) );
oa22f80 g539938 ( .a(n_28845), .b(FE_OFN410_n_28303), .c(n_1071), .d(FE_OFN76_n_27012), .o(n_29101) );
oa22f80 g539939 ( .a(n_29053), .b(n_28303), .c(n_686), .d(n_27449), .o(n_29252) );
oa22f80 g539940 ( .a(n_29123), .b(FE_OFN297_n_3069), .c(n_1081), .d(FE_OFN1117_rst), .o(n_29338) );
oa22f80 g539941 ( .a(n_28936), .b(n_4162), .c(n_265), .d(FE_OFN134_n_27449), .o(n_29176) );
oa22f80 g539942 ( .a(n_28935), .b(FE_OFN307_n_3069), .c(n_129), .d(FE_OFN99_n_27449), .o(n_29175) );
oa22f80 g539943 ( .a(n_29275), .b(FE_OFN313_n_3069), .c(n_911), .d(FE_OFN77_n_27012), .o(n_29522) );
oa22f80 g539944 ( .a(n_29122), .b(FE_OFN307_n_3069), .c(n_701), .d(FE_OFN64_n_27012), .o(n_29408) );
oa22f80 g539945 ( .a(n_29052), .b(n_28771), .c(n_1772), .d(FE_OFN138_n_27449), .o(n_29337) );
oa22f80 g539946 ( .a(n_29121), .b(FE_OFN303_n_3069), .c(n_1364), .d(FE_OFN335_n_4860), .o(n_29406) );
oa22f80 g539947 ( .a(n_29051), .b(FE_OFN313_n_3069), .c(n_1114), .d(FE_OFN1174_n_4860), .o(n_29336) );
oa22f80 g539948 ( .a(n_29120), .b(FE_OFN307_n_3069), .c(n_716), .d(FE_OFN357_n_4860), .o(n_29404) );
oa22f80 g539949 ( .a(n_28764), .b(FE_OFN296_n_3069), .c(n_1333), .d(FE_OFN80_n_27012), .o(n_29100) );
oa22f80 g539950 ( .a(n_28934), .b(n_29269), .c(n_404), .d(FE_OFN138_n_27449), .o(n_29251) );
oa22f80 g539951 ( .a(n_28933), .b(n_29269), .c(n_478), .d(FE_OFN1121_rst), .o(n_29250) );
oa22f80 g539952 ( .a(n_29119), .b(FE_OFN184_n_29402), .c(n_1174), .d(FE_OFN1114_rst), .o(n_29403) );
oa22f80 g539953 ( .a(n_29184), .b(FE_OFN183_n_29402), .c(n_1391), .d(FE_OFN1120_rst), .o(n_29463) );
oa22f80 g539954 ( .a(n_28844), .b(FE_OFN300_n_3069), .c(n_361), .d(FE_OFN1106_rst), .o(n_29174) );
oa22f80 g539955 ( .a(n_28843), .b(FE_OFN254_n_4280), .c(n_1183), .d(FE_OFN358_n_4860), .o(n_29171) );
oa22f80 g539956 ( .a(n_29118), .b(FE_OFN265_n_4280), .c(n_474), .d(FE_OFN353_n_4860), .o(n_29401) );
oa22f80 g539957 ( .a(n_29116), .b(FE_OFN239_n_4162), .c(n_130), .d(FE_OFN135_n_27449), .o(n_29400) );
oa22f80 g539958 ( .a(n_29115), .b(FE_OFN413_n_28303), .c(n_914), .d(FE_OFN78_n_27012), .o(n_29399) );
oa22f80 g539959 ( .a(n_29114), .b(FE_OFN412_n_28303), .c(n_1037), .d(FE_OFN91_n_27449), .o(n_29398) );
oa22f80 g539960 ( .a(n_29183), .b(FE_OFN265_n_4280), .c(n_1312), .d(FE_OFN128_n_27449), .o(n_29462) );
oa22f80 g539961 ( .a(n_28666), .b(FE_OFN410_n_28303), .c(n_804), .d(FE_OFN360_n_4860), .o(n_28981) );
oa22f80 g539962 ( .a(n_27834), .b(n_4280), .c(n_1702), .d(FE_OFN360_n_4860), .o(n_28324) );
oa22f80 g539963 ( .a(n_29113), .b(n_4280), .c(n_1618), .d(FE_OFN101_n_27449), .o(n_29396) );
oa22f80 g539964 ( .a(n_28842), .b(FE_OFN269_n_4280), .c(n_790), .d(FE_OFN115_n_27449), .o(n_29167) );
oa22f80 g539965 ( .a(n_29112), .b(FE_OFN264_n_4280), .c(n_933), .d(n_29264), .o(n_29394) );
ao22s80 g539966 ( .a(n_27992), .b(n_28400), .c(x_out_38_31), .d(n_5003), .o(n_28401) );
oa22f80 g539967 ( .a(n_28223), .b(n_28222), .c(n_28221), .d(x_in_20_13), .o(n_29390) );
ao22s80 g539968 ( .a(n_29277), .b(n_27652), .c(n_29278), .d(n_27651), .o(n_29515) );
no02f80 g540031 ( .a(n_29330), .b(n_29383), .o(n_29331) );
in01f80 g540032 ( .a(n_28393), .o(n_28394) );
na02f80 g540033 ( .a(n_28291), .b(x_in_60_14), .o(n_28393) );
no02f80 g540034 ( .a(n_28291), .b(x_in_60_14), .o(n_28603) );
no02f80 g540035 ( .a(n_29234), .b(n_29233), .o(n_29235) );
no02f80 g540036 ( .a(n_29328), .b(n_29327), .o(n_29329) );
no02f80 g540037 ( .a(n_29231), .b(FE_OFN1268_n_29314), .o(n_29232) );
no02f80 g540038 ( .a(n_29325), .b(n_29324), .o(n_29326) );
no02f80 g540039 ( .a(n_29322), .b(n_29321), .o(n_29323) );
no02f80 g540040 ( .a(n_29319), .b(n_29318), .o(n_29320) );
no02f80 g540041 ( .a(n_29229), .b(n_29228), .o(n_29230) );
no02f80 g540042 ( .a(n_29226), .b(n_29225), .o(n_29227) );
no02f80 g540043 ( .a(n_29156), .b(n_29155), .o(n_29157) );
na02f80 g540044 ( .a(n_28289), .b(x_in_6_15), .o(n_28290) );
no02f80 g540045 ( .a(n_29223), .b(n_29222), .o(n_29224) );
no02f80 g540046 ( .a(n_29220), .b(n_29219), .o(n_29221) );
no02f80 g540047 ( .a(n_29086), .b(n_29085), .o(n_29087) );
na02f80 g540048 ( .a(n_27984), .b(x_in_6_14), .o(n_28356) );
na02f80 g540049 ( .a(n_27985), .b(n_1489), .o(n_28482) );
no02f80 g540050 ( .a(n_28959), .b(n_29074), .o(n_28960) );
in01f80 g540051 ( .a(n_28198), .o(n_28199) );
na02f80 g540052 ( .a(n_28079), .b(x_in_32_14), .o(n_28198) );
no02f80 g540053 ( .a(n_28079), .b(x_in_32_14), .o(n_28361) );
no02f80 g540054 ( .a(n_29153), .b(n_29152), .o(n_29154) );
no02f80 g540055 ( .a(n_29150), .b(n_29186), .o(n_29151) );
in01f80 g540056 ( .a(n_28389), .o(n_28390) );
na02f80 g540057 ( .a(n_28288), .b(x_in_48_14), .o(n_28389) );
no02f80 g540058 ( .a(n_28288), .b(x_in_48_14), .o(n_28599) );
no02f80 g540059 ( .a(n_29082), .b(n_29081), .o(n_29083) );
no02f80 g540060 ( .a(n_28954), .b(n_29075), .o(n_28955) );
no02f80 g540061 ( .a(n_29316), .b(n_29315), .o(n_29317) );
no02f80 g540062 ( .a(n_29217), .b(n_29276), .o(n_29218) );
no02f80 g540063 ( .a(n_28221), .b(x_in_20_14), .o(n_28360) );
in01f80 g540064 ( .a(n_28181), .o(n_28182) );
na02f80 g540065 ( .a(n_28221), .b(x_in_20_14), .o(n_28181) );
na02f80 g540066 ( .a(n_28221), .b(x_in_20_15), .o(n_28060) );
no02f80 g540067 ( .a(n_28939), .b(n_28872), .o(n_28873) );
no02f80 g540068 ( .a(n_29386), .b(n_29385), .o(n_29387) );
no02f80 g540069 ( .a(n_27868), .b(n_28177), .o(n_29334) );
na02f80 g540070 ( .a(n_29425), .b(n_29194), .o(n_29506) );
no02f80 g540071 ( .a(n_29577), .b(n_29576), .o(n_29578) );
na02f80 g540072 ( .a(n_27706), .b(n_28047), .o(n_29065) );
na02f80 g540073 ( .a(n_27852), .b(n_6644), .o(n_28046) );
na02f80 g540074 ( .a(n_27853), .b(n_6645), .o(n_28173) );
no02f80 g540075 ( .a(n_28168), .b(n_29429), .o(n_28169) );
na02f80 g540076 ( .a(n_28039), .b(FE_OFN1109_rst), .o(n_28260) );
no02f80 g540077 ( .a(n_28254), .b(n_28036), .o(n_28037) );
oa12f80 g540078 ( .a(n_27962), .b(FE_OFN1268_n_29314), .c(n_28120), .o(n_29430) );
no02f80 g540079 ( .a(n_28247), .b(n_28034), .o(n_28035) );
no02f80 g540080 ( .a(n_28246), .b(n_28032), .o(n_28033) );
no02f80 g540081 ( .a(n_29234), .b(n_28030), .o(n_28031) );
oa12f80 g540082 ( .a(n_27627), .b(n_29075), .c(n_27865), .o(n_29188) );
ao12f80 g540083 ( .a(n_28223), .b(n_29332), .c(n_28222), .o(n_29504) );
oa12f80 g540084 ( .a(n_28006), .b(n_29248), .c(n_27827), .o(n_29551) );
oa12f80 g540085 ( .a(n_28119), .b(n_29247), .c(n_27960), .o(n_29548) );
oa12f80 g540086 ( .a(n_28118), .b(n_29246), .c(n_27958), .o(n_29545) );
oa12f80 g540087 ( .a(n_28117), .b(n_29245), .c(n_27956), .o(n_29542) );
oa12f80 g540088 ( .a(n_28005), .b(n_29166), .c(n_27822), .o(n_29519) );
oa12f80 g540089 ( .a(n_28002), .b(n_29165), .c(n_27819), .o(n_29516) );
oa12f80 g540090 ( .a(n_28116), .b(n_27954), .c(n_29092), .o(n_29459) );
oa12f80 g540091 ( .a(n_28001), .b(n_29164), .c(n_27817), .o(n_29512) );
oa12f80 g540092 ( .a(n_28115), .b(n_29163), .c(n_27952), .o(n_29509) );
oa12f80 g540093 ( .a(n_28114), .b(n_27950), .c(n_28966), .o(n_29455) );
oa12f80 g540094 ( .a(n_27814), .b(n_29381), .c(n_27383), .o(n_29487) );
oa12f80 g540095 ( .a(n_27635), .b(n_29379), .c(n_27191), .o(n_29484) );
oa12f80 g540096 ( .a(n_2709), .b(n_29451), .c(n_2152), .o(n_29538) );
oa12f80 g540097 ( .a(n_27634), .b(n_29214), .c(n_27189), .o(n_29365) );
oa12f80 g540098 ( .a(n_27633), .b(n_29377), .c(n_27187), .o(n_29481) );
oa12f80 g540099 ( .a(n_27632), .b(n_29375), .c(n_27185), .o(n_29478) );
oa12f80 g540100 ( .a(n_27631), .b(n_29373), .c(n_27183), .o(n_29475) );
oa12f80 g540101 ( .a(n_28113), .b(n_29091), .c(n_27946), .o(n_29427) );
in01f80 g540102 ( .a(n_29313), .o(n_29502) );
oa12f80 g540103 ( .a(n_28112), .b(n_28964), .c(n_27943), .o(n_29313) );
oa12f80 g540104 ( .a(n_27643), .b(n_29308), .c(n_27387), .o(n_29423) );
oa12f80 g540105 ( .a(n_27991), .b(n_611), .c(FE_OFN94_n_27449), .o(n_28144) );
oa12f80 g540106 ( .a(n_27757), .b(n_29212), .c(n_27271), .o(n_29362) );
ao12f80 g540107 ( .a(n_9560), .b(n_28009), .c(n_11547), .o(n_28021) );
ao12f80 g540108 ( .a(n_28227), .b(n_28265), .c(n_29383), .o(n_29581) );
ao12f80 g540109 ( .a(n_27941), .b(n_27995), .c(n_29074), .o(n_29333) );
oa12f80 g540110 ( .a(n_27715), .b(n_1825), .c(FE_OFN1146_n_4860), .o(n_28019) );
ao12f80 g540111 ( .a(n_29148), .b(n_29147), .c(n_29146), .o(n_29312) );
ao22s80 g540112 ( .a(n_29381), .b(n_27949), .c(n_29162), .d(n_27948), .o(n_29382) );
ao22s80 g540113 ( .a(n_29379), .b(n_27813), .c(n_29161), .d(n_27812), .o(n_29380) );
ao22s80 g540114 ( .a(n_29451), .b(n_3713), .c(n_29244), .d(n_3712), .o(n_29452) );
ao12f80 g540115 ( .a(n_29299), .b(n_29298), .c(n_29297), .o(n_29447) );
ao22s80 g540116 ( .a(n_29214), .b(n_27811), .c(n_28965), .d(n_27810), .o(n_29215) );
ao12f80 g540117 ( .a(n_29296), .b(n_29295), .c(n_29294), .o(n_29444) );
ao22s80 g540118 ( .a(n_29377), .b(n_27809), .c(n_29160), .d(n_27808), .o(n_29378) );
ao22s80 g540119 ( .a(n_29375), .b(n_27807), .c(n_29159), .d(n_27806), .o(n_29376) );
ao22s80 g540120 ( .a(n_29373), .b(n_27805), .c(n_29158), .d(n_27804), .o(n_29374) );
ao12f80 g540121 ( .a(n_29293), .b(n_29292), .c(n_29291), .o(n_29443) );
ao12f80 g540122 ( .a(n_29145), .b(n_29144), .c(n_29143), .o(n_29311) );
ao12f80 g540123 ( .a(n_29435), .b(n_29434), .c(FE_OFN1224_n_29433), .o(n_29567) );
ao12f80 g540124 ( .a(n_29290), .b(n_29289), .c(n_29288), .o(n_29442) );
ao12f80 g540125 ( .a(n_29203), .b(n_29202), .c(n_29201), .o(n_29372) );
ao12f80 g540126 ( .a(n_29287), .b(n_29286), .c(n_29285), .o(n_29441) );
ao12f80 g540127 ( .a(n_29200), .b(n_29199), .c(n_29198), .o(n_29371) );
ao12f80 g540128 ( .a(n_29284), .b(n_29283), .c(n_29282), .o(n_29440) );
ao12f80 g540129 ( .a(n_27864), .b(n_27863), .c(FE_OFN716_n_29187), .o(n_29448) );
ao12f80 g540130 ( .a(n_29142), .b(n_29141), .c(n_29140), .o(n_29310) );
ao12f80 g540131 ( .a(n_29281), .b(n_29280), .c(n_29279), .o(n_29439) );
ao12f80 g540132 ( .a(n_28109), .b(n_28108), .c(n_29456), .o(n_29534) );
ao12f80 g540133 ( .a(n_29197), .b(n_29196), .c(n_29195), .o(n_29370) );
ao12f80 g540134 ( .a(n_28851), .b(n_28850), .c(n_28849), .o(n_29071) );
in01f80 g540135 ( .a(n_28354), .o(n_28476) );
oa22f80 g540136 ( .a(n_27612), .b(n_12284), .c(n_28009), .d(n_12285), .o(n_28354) );
in01f80 g540137 ( .a(n_29135), .o(n_29070) );
ao22s80 g540138 ( .a(n_28715), .b(n_27667), .c(n_28939), .d(x_in_52_13), .o(n_29135) );
ao22s80 g540139 ( .a(n_29212), .b(n_27909), .c(n_28963), .d(n_27908), .o(n_29213) );
ao22s80 g540140 ( .a(n_29308), .b(n_27831), .c(n_29090), .d(n_27830), .o(n_29309) );
ao12f80 g540141 ( .a(n_29139), .b(n_29138), .c(n_29137), .o(n_29307) );
oa22f80 g540142 ( .a(n_29088), .b(FE_OFN184_n_29402), .c(n_1487), .d(FE_OFN347_n_4860), .o(n_29306) );
oa22f80 g540143 ( .a(n_28962), .b(FE_OFN184_n_29402), .c(n_735), .d(FE_OFN347_n_4860), .o(n_29211) );
oa22f80 g540144 ( .a(n_28958), .b(FE_OFN409_n_28303), .c(n_566), .d(FE_OFN125_n_27449), .o(n_29210) );
oa22f80 g540145 ( .a(n_29084), .b(n_29683), .c(n_105), .d(FE_OFN105_n_27449), .o(n_29305) );
oa22f80 g540146 ( .a(n_29149), .b(n_29683), .c(n_711), .d(FE_OFN105_n_27449), .o(n_29368) );
oa22f80 g540147 ( .a(n_28957), .b(FE_OFN411_n_28303), .c(n_1875), .d(FE_OFN192_n_28928), .o(n_29208) );
oa22f80 g540148 ( .a(n_28804), .b(FE_OFN306_n_3069), .c(n_1121), .d(FE_OFN14_n_29068), .o(n_29069) );
oa22f80 g540149 ( .a(n_29080), .b(FE_OFN412_n_28303), .c(n_1533), .d(FE_OFN329_n_4860), .o(n_29304) );
oa22f80 g540150 ( .a(n_27784), .b(FE_OFN260_n_4280), .c(n_1587), .d(FE_OFN355_n_4860), .o(n_28124) );
oa22f80 g540151 ( .a(n_28953), .b(FE_OFN256_n_4280), .c(n_1598), .d(FE_OFN358_n_4860), .o(n_29207) );
oa22f80 g540152 ( .a(n_29078), .b(FE_OFN234_n_4162), .c(n_115), .d(FE_OFN74_n_27012), .o(n_29302) );
oa22f80 g540153 ( .a(n_28952), .b(FE_OFN268_n_4280), .c(n_371), .d(FE_OFN329_n_4860), .o(n_29206) );
oa22f80 g540154 ( .a(n_28950), .b(FE_OFN254_n_4280), .c(n_732), .d(FE_OFN11_n_29204), .o(n_29205) );
oa22f80 g540155 ( .a(FE_OFN634_n_27731), .b(FE_OFN265_n_4280), .c(n_681), .d(FE_OFN11_n_29204), .o(n_27732) );
oa22f80 g540156 ( .a(n_27717), .b(x_in_20_15), .c(FE_OFN634_n_27731), .d(n_1140), .o(n_29471) );
na02f80 g540174 ( .a(n_28006), .b(n_27828), .o(n_29328) );
no02f80 g540175 ( .a(n_27963), .b(n_28120), .o(n_29231) );
na02f80 g540176 ( .a(n_28119), .b(n_27961), .o(n_29325) );
na02f80 g540177 ( .a(n_28118), .b(n_27959), .o(n_29322) );
na02f80 g540178 ( .a(n_28117), .b(n_27957), .o(n_29319) );
na02f80 g540179 ( .a(n_28005), .b(n_27823), .o(n_29229) );
na02f80 g540180 ( .a(n_28116), .b(n_27955), .o(n_29156) );
na02f80 g540181 ( .a(n_28002), .b(n_27820), .o(n_29226) );
na02f80 g540182 ( .a(n_28001), .b(n_27818), .o(n_29223) );
na02f80 g540183 ( .a(n_28115), .b(n_27953), .o(n_29220) );
na02f80 g540184 ( .a(n_28114), .b(n_27951), .o(n_29086) );
no02f80 g540185 ( .a(n_29147), .b(n_29146), .o(n_29148) );
no02f80 g540186 ( .a(n_29298), .b(n_29297), .o(n_29299) );
no02f80 g540187 ( .a(n_29295), .b(n_29294), .o(n_29296) );
no02f80 g540188 ( .a(n_29292), .b(n_29291), .o(n_29293) );
no02f80 g540189 ( .a(n_29144), .b(n_29143), .o(n_29145) );
no02f80 g540190 ( .a(n_29289), .b(n_29288), .o(n_29290) );
no02f80 g540191 ( .a(n_29434), .b(FE_OFN1224_n_29433), .o(n_29435) );
no02f80 g540192 ( .a(n_29202), .b(n_29201), .o(n_29203) );
no02f80 g540193 ( .a(n_29286), .b(n_29285), .o(n_29287) );
no02f80 g540194 ( .a(n_29283), .b(n_29282), .o(n_29284) );
no02f80 g540195 ( .a(n_29199), .b(n_29198), .o(n_29200) );
no02f80 g540196 ( .a(n_29141), .b(n_29140), .o(n_29142) );
na02f80 g540197 ( .a(n_28113), .b(n_27947), .o(n_29153) );
no02f80 g540198 ( .a(n_29280), .b(n_29279), .o(n_29281) );
na02f80 g540199 ( .a(n_28112), .b(n_27944), .o(n_29082) );
no02f80 g540200 ( .a(n_29196), .b(n_29195), .o(n_29197) );
no02f80 g540201 ( .a(n_28093), .b(n_28266), .o(n_29217) );
in01f80 g540202 ( .a(n_27867), .o(n_27868) );
na02f80 g540203 ( .a(n_27717), .b(x_in_20_14), .o(n_27867) );
no02f80 g540204 ( .a(n_27717), .b(x_in_20_14), .o(n_28177) );
no02f80 g540205 ( .a(n_29138), .b(n_29137), .o(n_29139) );
na03f80 g540206 ( .a(n_27175), .b(FE_OFN634_n_27731), .c(FE_OFN1182_rst), .o(n_27715) );
no02f80 g540207 ( .a(n_27628), .b(n_27865), .o(n_28954) );
in01f80 g540208 ( .a(n_28110), .o(n_28111) );
na02f80 g540209 ( .a(n_27801), .b(n_27996), .o(n_28110) );
na02f80 g540210 ( .a(n_28226), .b(n_28265), .o(n_29330) );
na02f80 g540211 ( .a(n_27940), .b(n_27995), .o(n_28959) );
na02f80 g540212 ( .a(n_28224), .b(n_28264), .o(n_29150) );
in01f80 g540213 ( .a(n_27705), .o(n_27706) );
no02f80 g540214 ( .a(FE_OFN634_n_27731), .b(n_28222), .o(n_27705) );
na02f80 g540215 ( .a(FE_OFN634_n_27731), .b(n_28222), .o(n_28047) );
no02f80 g540216 ( .a(n_28850), .b(n_28849), .o(n_28851) );
no02f80 g540217 ( .a(n_27863), .b(FE_OFN716_n_29187), .o(n_27864) );
in01f80 g540218 ( .a(n_27993), .o(n_27994) );
no02f80 g540219 ( .a(n_27862), .b(n_2022), .o(n_27993) );
in01f80 g540220 ( .a(n_27991), .o(n_27992) );
na02f80 g540221 ( .a(n_27862), .b(FE_OFN34_n_15183), .o(n_27991) );
no02f80 g540222 ( .a(n_27618), .b(FE_OFN368_n_26312), .o(n_27861) );
oa12f80 g540223 ( .a(FE_OFN32_n_27986), .b(n_1952), .c(FE_OFN193_n_28928), .o(n_27990) );
oa12f80 g540224 ( .a(n_27986), .b(n_726), .c(FE_OFN119_n_27449), .o(n_27987) );
no02f80 g540225 ( .a(n_28108), .b(n_29456), .o(n_28109) );
na02f80 g540226 ( .a(n_27783), .b(n_28400), .o(n_28391) );
oa22f80 g540227 ( .a(n_28745), .b(n_29194), .c(n_28944), .d(n_27231), .o(n_29386) );
oa12f80 g540228 ( .a(n_27910), .b(n_27482), .c(n_28932), .o(n_29186) );
oa12f80 g540229 ( .a(n_27363), .b(n_29117), .c(n_26919), .o(n_29316) );
oa12f80 g540230 ( .a(n_27401), .b(n_27789), .c(n_26109), .o(n_27860) );
oa12f80 g540231 ( .a(n_27692), .b(n_1550), .c(FE_OFN330_n_4860), .o(n_27694) );
oa12f80 g540232 ( .a(n_27692), .b(n_249), .c(FE_OFN288_n_29266), .o(n_27693) );
oa12f80 g540233 ( .a(n_27396), .b(n_1102), .c(FE_OFN1113_rst), .o(n_27687) );
in01f80 g540234 ( .a(n_29277), .o(n_29278) );
ao12f80 g540235 ( .a(n_29190), .b(n_29076), .c(x_in_36_12), .o(n_29277) );
in01f80 g540236 ( .a(n_28223), .o(n_28221) );
oa12f80 g540237 ( .a(FE_OFN634_n_27731), .b(n_26969), .c(n_27211), .o(n_28223) );
in01f80 g540238 ( .a(n_29425), .o(n_29577) );
no02f80 g540239 ( .a(n_29249), .b(n_29190), .o(n_29425) );
oa12f80 g540240 ( .a(n_27797), .b(n_27829), .c(n_27939), .o(n_28291) );
ao12f80 g540241 ( .a(n_28909), .b(n_28908), .c(n_28907), .o(n_29067) );
oa12f80 g540242 ( .a(n_27436), .b(n_27435), .c(x_in_58_15), .o(n_29234) );
ao12f80 g540243 ( .a(n_29019), .b(n_29018), .c(n_29017), .o(n_29134) );
ao12f80 g540244 ( .a(n_29016), .b(FE_OFN1270_n_29015), .c(n_29089), .o(n_29133) );
ao12f80 g540245 ( .a(n_29014), .b(n_29013), .c(n_29012), .o(n_29132) );
oa12f80 g540246 ( .a(n_27938), .b(n_27937), .c(FE_OFN1224_n_29433), .o(n_29547) );
ao12f80 g540247 ( .a(n_29011), .b(n_29010), .c(n_29009), .o(n_29131) );
ao12f80 g540248 ( .a(n_29008), .b(n_29007), .c(n_29006), .o(n_29130) );
ao12f80 g540249 ( .a(n_28090), .b(n_28089), .c(n_29279), .o(n_29541) );
ao12f80 g540250 ( .a(n_28906), .b(n_28905), .c(n_28904), .o(n_29061) );
oa12f80 g540251 ( .a(n_27438), .b(n_27437), .c(x_in_60_15), .o(n_29429) );
ao12f80 g540252 ( .a(n_28818), .b(n_28817), .c(n_28816), .o(n_28937) );
ao12f80 g540253 ( .a(n_28903), .b(n_28902), .c(n_28901), .o(n_29060) );
oa12f80 g540254 ( .a(n_27796), .b(n_27795), .c(n_27794), .o(n_28289) );
ao12f80 g540255 ( .a(n_28900), .b(n_28899), .c(n_28898), .o(n_29059) );
ao12f80 g540256 ( .a(n_28897), .b(n_28896), .c(n_28895), .o(n_29058) );
ao12f80 g540257 ( .a(n_28735), .b(n_28734), .c(n_28733), .o(n_28847) );
in01f80 g540258 ( .a(n_27984), .o(n_27985) );
oa12f80 g540259 ( .a(n_27623), .b(n_27622), .c(n_27857), .o(n_27984) );
ao12f80 g540260 ( .a(n_28894), .b(n_28893), .c(n_28892), .o(n_29057) );
ao12f80 g540261 ( .a(n_28891), .b(n_28890), .c(n_28889), .o(n_29056) );
ao12f80 g540262 ( .a(n_29005), .b(n_29004), .c(n_29003), .o(n_29126) );
ao12f80 g540263 ( .a(n_29002), .b(n_29001), .c(n_29000), .o(n_29125) );
ao12f80 g540264 ( .a(n_28732), .b(n_28731), .c(n_28730), .o(n_28846) );
ao12f80 g540265 ( .a(n_28999), .b(n_28998), .c(n_28997), .o(n_29124) );
ao12f80 g540266 ( .a(n_28729), .b(n_28728), .c(n_28806), .o(n_28845) );
ao12f80 g540267 ( .a(n_28888), .b(n_28887), .c(n_28886), .o(n_29055) );
ao12f80 g540268 ( .a(n_28885), .b(n_28884), .c(n_28883), .o(n_29054) );
ao12f80 g540269 ( .a(n_28882), .b(n_28881), .c(n_28880), .o(n_29053) );
in01f80 g540270 ( .a(n_27852), .o(n_27853) );
oa12f80 g540271 ( .a(n_27431), .b(n_27430), .c(n_27429), .o(n_27852) );
ao12f80 g540272 ( .a(n_28996), .b(n_28995), .c(n_28994), .o(n_29123) );
ao12f80 g540273 ( .a(n_28815), .b(n_28814), .c(n_28813), .o(n_28936) );
oa22f80 g540274 ( .a(n_26928), .b(FE_OFN308_n_3069), .c(n_18), .d(FE_OFN1114_rst), .o(n_27503) );
ao12f80 g540275 ( .a(n_28812), .b(n_28811), .c(n_28810), .o(n_28935) );
ao12f80 g540276 ( .a(n_29170), .b(n_29169), .c(n_29168), .o(n_29275) );
ao12f80 g540277 ( .a(n_28993), .b(n_28992), .c(n_28991), .o(n_29122) );
in01f80 g540278 ( .a(n_27675), .o(n_28039) );
ao12f80 g540279 ( .a(n_27215), .b(n_27214), .c(n_27213), .o(n_27675) );
ao12f80 g540280 ( .a(n_28879), .b(n_28878), .c(n_28877), .o(n_29052) );
ao12f80 g540281 ( .a(n_28990), .b(n_28989), .c(n_28988), .o(n_29121) );
ao12f80 g540282 ( .a(n_28876), .b(n_28875), .c(n_28874), .o(n_29051) );
ao12f80 g540283 ( .a(n_28987), .b(n_28986), .c(n_28985), .o(n_29120) );
ao12f80 g540284 ( .a(n_28639), .b(n_28638), .c(n_28637), .o(n_28764) );
oa12f80 g540285 ( .a(n_27403), .b(n_27624), .c(n_27402), .o(n_28079) );
ao12f80 g540286 ( .a(n_28809), .b(n_28808), .c(n_28807), .o(n_28934) );
ao22s80 g540287 ( .a(n_28023), .b(n_28932), .c(n_28022), .d(n_28709), .o(n_28933) );
oa12f80 g540288 ( .a(n_27793), .b(n_27936), .c(n_27792), .o(n_28288) );
ao12f80 g540289 ( .a(n_28984), .b(n_28983), .c(n_28982), .o(n_29119) );
ao12f80 g540290 ( .a(n_29098), .b(n_29097), .c(n_29096), .o(n_29184) );
ao12f80 g540291 ( .a(n_28727), .b(n_28726), .c(n_28725), .o(n_28844) );
oa12f80 g540292 ( .a(n_27629), .b(n_27630), .c(x_in_40_15), .o(n_29612) );
ao12f80 g540293 ( .a(n_28724), .b(n_28723), .c(n_28805), .o(n_28843) );
ao22s80 g540294 ( .a(n_29117), .b(n_27575), .c(n_28859), .d(n_27574), .o(n_29118) );
ao12f80 g540295 ( .a(n_28980), .b(n_28979), .c(n_28978), .o(n_29116) );
in01f80 g540296 ( .a(n_28254), .o(n_27851) );
ao12f80 g540297 ( .a(n_27423), .b(n_27422), .c(x_in_10_15), .o(n_28254) );
ao12f80 g540298 ( .a(n_28977), .b(n_28976), .c(n_29050), .o(n_29115) );
ao22s80 g540299 ( .a(n_28777), .b(n_27570), .c(n_29050), .d(x_in_48_13), .o(n_29276) );
oa22f80 g540300 ( .a(n_26945), .b(n_26927), .c(n_1700), .d(FE_OFN114_n_27449), .o(n_27485) );
ao12f80 g540301 ( .a(n_28975), .b(n_28974), .c(n_28973), .o(n_29114) );
in01f80 g540302 ( .a(n_28247), .o(n_27842) );
ao12f80 g540303 ( .a(n_27419), .b(n_27418), .c(x_in_42_15), .o(n_28247) );
ao12f80 g540304 ( .a(n_29095), .b(n_29094), .c(n_29093), .o(n_29183) );
ao12f80 g540305 ( .a(n_28972), .b(n_28971), .c(n_28970), .o(n_29113) );
ao12f80 g540306 ( .a(n_28520), .b(n_28519), .c(n_28518), .o(n_28666) );
oa12f80 g540307 ( .a(n_27406), .b(n_27667), .c(x_in_52_13), .o(n_28872) );
in01f80 g540308 ( .a(n_28246), .o(n_27835) );
ao12f80 g540309 ( .a(n_27416), .b(n_27415), .c(x_in_26_15), .o(n_28246) );
ao12f80 g540310 ( .a(n_27621), .b(n_27620), .c(n_27619), .o(n_27834) );
ao12f80 g540311 ( .a(n_28722), .b(n_28721), .c(n_28720), .o(n_28842) );
ao12f80 g540312 ( .a(n_28969), .b(n_28968), .c(n_28967), .o(n_29112) );
oa22f80 g540313 ( .a(n_28707), .b(n_29046), .c(n_86), .d(FE_OFN92_n_27449), .o(n_28931) );
oa22f80 g540314 ( .a(FE_OFN1136_n_28794), .b(n_29046), .c(n_791), .d(n_27449), .o(n_29049) );
oa22f80 g540315 ( .a(n_28795), .b(n_29046), .c(n_902), .d(FE_OFN326_n_4860), .o(n_29047) );
oa22f80 g540316 ( .a(n_28793), .b(FE_OFN254_n_4280), .c(n_602), .d(FE_OFN1124_rst), .o(n_29045) );
oa22f80 g540317 ( .a(n_28940), .b(FE_OFN260_n_4280), .c(n_553), .d(FE_OFN1120_rst), .o(n_29180) );
oa22f80 g540318 ( .a(n_28792), .b(FE_OFN254_n_4280), .c(n_1928), .d(FE_OFN285_n_29266), .o(n_29043) );
oa22f80 g540319 ( .a(n_28791), .b(FE_OFN166_n_29269), .c(n_662), .d(FE_OFN90_n_27449), .o(n_29042) );
oa22f80 g540320 ( .a(n_28706), .b(n_29269), .c(n_1176), .d(n_28928), .o(n_28929) );
oa22f80 g540321 ( .a(n_28630), .b(n_29046), .c(n_332), .d(n_27449), .o(n_28841) );
oa22f80 g540322 ( .a(n_28705), .b(FE_OFN269_n_4280), .c(n_1906), .d(FE_OFN1114_rst), .o(n_28926) );
oa22f80 g540323 ( .a(n_28704), .b(n_29046), .c(n_1911), .d(FE_OFN1115_rst), .o(n_28925) );
oa22f80 g540324 ( .a(FE_OFN1021_n_28703), .b(n_29046), .c(n_1806), .d(FE_OFN60_n_27012), .o(n_28923) );
oa22f80 g540325 ( .a(n_28493), .b(FE_OFN296_n_3069), .c(n_966), .d(FE_OFN352_n_4860), .o(n_28758) );
oa22f80 g540326 ( .a(n_28702), .b(FE_OFN183_n_29402), .c(n_1690), .d(FE_OFN363_n_4860), .o(n_28921) );
oa22f80 g540327 ( .a(n_28701), .b(FE_OFN296_n_3069), .c(n_885), .d(FE_OFN352_n_4860), .o(n_28920) );
oa22f80 g540328 ( .a(n_28790), .b(FE_OFN300_n_3069), .c(n_169), .d(FE_OFN329_n_4860), .o(n_29039) );
oa22f80 g540329 ( .a(n_28789), .b(FE_OFN294_n_3069), .c(n_182), .d(FE_OFN363_n_4860), .o(n_29038) );
oa22f80 g540330 ( .a(n_28491), .b(FE_OFN307_n_3069), .c(n_459), .d(FE_OFN1112_rst), .o(n_28752) );
oa22f80 g540331 ( .a(n_28788), .b(FE_OFN309_n_3069), .c(n_251), .d(FE_OFN364_n_4860), .o(n_29037) );
oa22f80 g540332 ( .a(n_28700), .b(FE_OFN293_n_3069), .c(n_1239), .d(FE_OFN64_n_27012), .o(n_28919) );
oa22f80 g540333 ( .a(n_28492), .b(FE_OFN295_n_3069), .c(n_1552), .d(FE_OFN74_n_27012), .o(n_28748) );
oa22f80 g540334 ( .a(n_28699), .b(FE_OFN266_n_4280), .c(n_1240), .d(FE_OFN114_n_27449), .o(n_28917) );
oa22f80 g540335 ( .a(n_28698), .b(FE_OFN165_n_29269), .c(n_651), .d(n_28607), .o(n_28915) );
oa22f80 g540336 ( .a(n_28787), .b(n_29269), .c(n_789), .d(FE_OFN1117_rst), .o(n_29035) );
oa22f80 g540337 ( .a(FE_OFN1131_n_28629), .b(n_29033), .c(n_805), .d(FE_OFN63_n_27012), .o(n_28830) );
oa22f80 g540338 ( .a(n_28697), .b(FE_OFN404_n_28303), .c(n_1413), .d(FE_OFN363_n_4860), .o(n_28914) );
oa22f80 g540339 ( .a(FE_OFN1132_n_28627), .b(n_29033), .c(n_67), .d(FE_OFN324_n_4860), .o(n_28827) );
oa22f80 g540340 ( .a(FE_OFN1138_n_28938), .b(n_29033), .c(n_444), .d(FE_OFN95_n_27449), .o(n_29179) );
oa22f80 g540341 ( .a(n_28786), .b(n_29033), .c(n_1194), .d(n_27449), .o(n_29034) );
oa22f80 g540342 ( .a(FE_OFN945_n_27398), .b(n_28608), .c(n_903), .d(FE_OFN95_n_27449), .o(n_27458) );
oa22f80 g540343 ( .a(n_28696), .b(n_29033), .c(n_368), .d(FE_OFN95_n_27449), .o(n_28913) );
oa22f80 g540344 ( .a(n_28785), .b(FE_OFN184_n_29402), .c(n_1653), .d(FE_OFN56_n_27012), .o(n_29031) );
oa22f80 g540345 ( .a(n_28695), .b(FE_OFN183_n_29402), .c(n_967), .d(FE_OFN80_n_27012), .o(n_28911) );
oa22f80 g540346 ( .a(n_28784), .b(FE_OFN293_n_3069), .c(n_1588), .d(FE_OFN64_n_27012), .o(n_29030) );
oa22f80 g540347 ( .a(n_28369), .b(n_29033), .c(n_1845), .d(FE_OFN63_n_27012), .o(n_28652) );
oa22f80 g540348 ( .a(n_28626), .b(n_29033), .c(n_1299), .d(FE_OFN63_n_27012), .o(n_28822) );
oa22f80 g540349 ( .a(n_28625), .b(FE_OFN253_n_4280), .c(n_1841), .d(FE_OFN138_n_27449), .o(n_28821) );
oa22f80 g540350 ( .a(n_28624), .b(FE_OFN240_n_4162), .c(n_516), .d(FE_OFN141_n_27449), .o(n_28819) );
oa22f80 g540351 ( .a(n_28783), .b(FE_OFN269_n_4280), .c(n_1749), .d(FE_OFN90_n_27449), .o(n_29029) );
oa22f80 g540352 ( .a(n_28857), .b(FE_OFN295_n_3069), .c(n_450), .d(FE_OFN130_n_27449), .o(n_29109) );
oa22f80 g540353 ( .a(n_28490), .b(FE_OFN293_n_3069), .c(n_985), .d(FE_OFN89_n_27449), .o(n_28741) );
oa22f80 g540354 ( .a(n_28489), .b(FE_OFN244_n_4162), .c(n_329), .d(FE_OFN108_n_27449), .o(n_28740) );
oa22f80 g540355 ( .a(FE_OFN1133_n_28782), .b(FE_OFN1151_n_3069), .c(n_199), .d(n_29104), .o(n_29027) );
oa22f80 g540356 ( .a(n_28780), .b(FE_OFN259_n_4280), .c(n_717), .d(FE_OFN1120_rst), .o(n_29026) );
oa22f80 g540357 ( .a(n_28779), .b(FE_OFN258_n_4280), .c(n_531), .d(FE_OFN1121_rst), .o(n_29024) );
oa22f80 g540358 ( .a(n_28775), .b(FE_OFN267_n_4280), .c(n_894), .d(FE_OFN90_n_27449), .o(n_29023) );
oa22f80 g540359 ( .a(n_28855), .b(FE_OFN265_n_4280), .c(n_563), .d(FE_OFN128_n_27449), .o(n_29106) );
oa22f80 g540360 ( .a(n_28694), .b(n_4280), .c(n_567), .d(FE_OFN100_n_27449), .o(n_28910) );
oa22f80 g540361 ( .a(n_28854), .b(FE_OFN303_n_3069), .c(n_1586), .d(n_29104), .o(n_29105) );
oa22f80 g540362 ( .a(n_28267), .b(FE_OFN295_n_3069), .c(n_506), .d(FE_OFN130_n_27449), .o(n_28527) );
oa22f80 g540363 ( .a(n_28774), .b(FE_OFN183_n_29402), .c(n_53), .d(FE_OFN101_n_27449), .o(n_29021) );
oa22f80 g540364 ( .a(n_27157), .b(FE_OFN183_n_29402), .c(n_995), .d(FE_OFN100_n_27449), .o(n_27647) );
oa22f80 g540365 ( .a(n_28488), .b(FE_OFN414_n_28303), .c(n_1908), .d(FE_OFN115_n_27449), .o(n_28736) );
oa22f80 g540366 ( .a(n_28773), .b(FE_OFN412_n_28303), .c(n_877), .d(FE_OFN119_n_27449), .o(n_29020) );
in01f80 g540444 ( .a(n_27962), .o(n_27963) );
na02f80 g540445 ( .a(n_27829), .b(x_in_60_14), .o(n_27962) );
no02f80 g540446 ( .a(n_27829), .b(x_in_60_14), .o(n_28120) );
na02f80 g540447 ( .a(n_27437), .b(x_in_60_15), .o(n_27438) );
no02f80 g540448 ( .a(n_28908), .b(n_28907), .o(n_28909) );
na02f80 g540449 ( .a(n_27435), .b(x_in_58_15), .o(n_27436) );
no02f80 g540450 ( .a(n_29018), .b(n_29017), .o(n_29019) );
na02f80 g540451 ( .a(n_27642), .b(x_in_2_14), .o(n_28006) );
in01f80 g540452 ( .a(n_27827), .o(n_27828) );
no02f80 g540453 ( .a(n_27642), .b(x_in_2_14), .o(n_27827) );
no02f80 g540454 ( .a(FE_OFN1270_n_29015), .b(n_29089), .o(n_29016) );
no02f80 g540455 ( .a(n_29013), .b(n_29012), .o(n_29014) );
na02f80 g540456 ( .a(n_27826), .b(x_in_34_14), .o(n_28119) );
in01f80 g540457 ( .a(n_27960), .o(n_27961) );
no02f80 g540458 ( .a(n_27826), .b(x_in_34_14), .o(n_27960) );
no02f80 g540459 ( .a(n_29010), .b(n_29009), .o(n_29011) );
na02f80 g540460 ( .a(n_27825), .b(x_in_18_14), .o(n_28118) );
in01f80 g540461 ( .a(n_27958), .o(n_27959) );
no02f80 g540462 ( .a(n_27825), .b(x_in_18_14), .o(n_27958) );
no02f80 g540463 ( .a(n_29007), .b(n_29006), .o(n_29008) );
na02f80 g540464 ( .a(n_27824), .b(x_in_50_14), .o(n_28117) );
in01f80 g540465 ( .a(n_27956), .o(n_27957) );
no02f80 g540466 ( .a(n_27824), .b(x_in_50_14), .o(n_27956) );
no02f80 g540467 ( .a(n_28905), .b(n_28904), .o(n_28906) );
na02f80 g540468 ( .a(n_27638), .b(x_in_10_14), .o(n_28005) );
in01f80 g540469 ( .a(n_27822), .o(n_27823) );
no02f80 g540470 ( .a(n_27638), .b(x_in_10_14), .o(n_27822) );
no02f80 g540471 ( .a(n_28817), .b(n_28816), .o(n_28818) );
na02f80 g540472 ( .a(n_27821), .b(x_in_6_14), .o(n_28116) );
no02f80 g540473 ( .a(n_28902), .b(n_28901), .o(n_28903) );
na02f80 g540474 ( .a(n_27637), .b(x_in_42_14), .o(n_28002) );
in01f80 g540475 ( .a(n_27819), .o(n_27820) );
no02f80 g540476 ( .a(n_27637), .b(x_in_42_14), .o(n_27819) );
in01f80 g540477 ( .a(n_27954), .o(n_27955) );
no02f80 g540478 ( .a(n_27821), .b(x_in_6_14), .o(n_27954) );
no02f80 g540479 ( .a(n_28899), .b(n_28898), .o(n_28900) );
na02f80 g540480 ( .a(n_27636), .b(x_in_26_14), .o(n_28001) );
in01f80 g540481 ( .a(n_27817), .o(n_27818) );
no02f80 g540482 ( .a(n_27636), .b(x_in_26_14), .o(n_27817) );
no02f80 g540483 ( .a(n_28896), .b(n_28895), .o(n_28897) );
na02f80 g540484 ( .a(n_27816), .b(x_in_58_14), .o(n_28115) );
in01f80 g540485 ( .a(n_27952), .o(n_27953) );
no02f80 g540486 ( .a(n_27816), .b(x_in_58_14), .o(n_27952) );
no02f80 g540487 ( .a(n_28734), .b(n_28733), .o(n_28735) );
na02f80 g540488 ( .a(n_27815), .b(x_in_6_13), .o(n_28114) );
in01f80 g540489 ( .a(n_27950), .o(n_27951) );
no02f80 g540490 ( .a(n_27815), .b(x_in_6_13), .o(n_27950) );
no02f80 g540491 ( .a(n_28893), .b(n_28892), .o(n_28894) );
in01f80 g540492 ( .a(n_27948), .o(n_27949) );
na02f80 g540493 ( .a(n_27384), .b(n_27814), .o(n_27948) );
no02f80 g540494 ( .a(n_28890), .b(n_28889), .o(n_28891) );
in01f80 g540495 ( .a(n_27812), .o(n_27813) );
na02f80 g540496 ( .a(n_27192), .b(n_27635), .o(n_27812) );
no02f80 g540497 ( .a(n_29004), .b(n_29003), .o(n_29005) );
no02f80 g540498 ( .a(n_29001), .b(n_29000), .o(n_29002) );
no02f80 g540499 ( .a(n_28731), .b(n_28730), .o(n_28732) );
in01f80 g540500 ( .a(n_27810), .o(n_27811) );
na02f80 g540501 ( .a(n_27190), .b(n_27634), .o(n_27810) );
no02f80 g540502 ( .a(n_28998), .b(n_28997), .o(n_28999) );
no02f80 g540503 ( .a(n_28887), .b(n_28886), .o(n_28888) );
in01f80 g540504 ( .a(n_27808), .o(n_27809) );
na02f80 g540505 ( .a(n_27188), .b(n_27633), .o(n_27808) );
no02f80 g540506 ( .a(n_28884), .b(n_28883), .o(n_28885) );
in01f80 g540507 ( .a(n_27806), .o(n_27807) );
na02f80 g540508 ( .a(n_27186), .b(n_27632), .o(n_27806) );
no02f80 g540509 ( .a(n_28728), .b(n_28806), .o(n_28729) );
no02f80 g540510 ( .a(n_28881), .b(n_28880), .o(n_28882) );
in01f80 g540511 ( .a(n_27804), .o(n_27805) );
na02f80 g540512 ( .a(n_27184), .b(n_27631), .o(n_27804) );
no02f80 g540513 ( .a(n_28995), .b(n_28994), .o(n_28996) );
na02f80 g540514 ( .a(n_27430), .b(n_27429), .o(n_27431) );
no02f80 g540515 ( .a(n_28814), .b(n_28813), .o(n_28815) );
no02f80 g540516 ( .a(n_28811), .b(n_28810), .o(n_28812) );
no02f80 g540517 ( .a(n_29169), .b(n_29168), .o(n_29170) );
no02f80 g540518 ( .a(n_28992), .b(n_28991), .o(n_28993) );
no02f80 g540519 ( .a(n_28878), .b(n_28877), .o(n_28879) );
no02f80 g540520 ( .a(n_28989), .b(n_28988), .o(n_28990) );
no02f80 g540521 ( .a(n_28875), .b(n_28874), .o(n_28876) );
no02f80 g540522 ( .a(n_28986), .b(n_28985), .o(n_28987) );
no02f80 g540523 ( .a(n_28638), .b(n_28637), .o(n_28639) );
no02f80 g540524 ( .a(n_28808), .b(n_28807), .o(n_28809) );
na02f80 g540525 ( .a(n_27803), .b(x_in_16_14), .o(n_28113) );
in01f80 g540526 ( .a(n_27946), .o(n_27947) );
no02f80 g540527 ( .a(n_27803), .b(x_in_16_14), .o(n_27946) );
no02f80 g540528 ( .a(n_28983), .b(n_28982), .o(n_28984) );
no02f80 g540529 ( .a(n_29097), .b(n_29096), .o(n_29098) );
no02f80 g540530 ( .a(n_28726), .b(n_28725), .o(n_28727) );
na02f80 g540531 ( .a(n_27802), .b(x_in_40_13), .o(n_28112) );
in01f80 g540532 ( .a(n_27943), .o(n_27944) );
no02f80 g540533 ( .a(n_27802), .b(x_in_40_13), .o(n_27943) );
in01f80 g540534 ( .a(n_27800), .o(n_27801) );
no02f80 g540535 ( .a(n_27630), .b(x_in_40_14), .o(n_27800) );
na02f80 g540536 ( .a(n_27630), .b(x_in_40_14), .o(n_27996) );
na02f80 g540537 ( .a(n_27630), .b(x_in_40_15), .o(n_27629) );
no02f80 g540538 ( .a(n_28723), .b(n_28805), .o(n_28724) );
in01f80 g540539 ( .a(n_27627), .o(n_27628) );
na02f80 g540540 ( .a(n_27426), .b(x_in_32_14), .o(n_27627) );
no02f80 g540541 ( .a(n_27426), .b(x_in_32_14), .o(n_27865) );
no02f80 g540542 ( .a(n_28979), .b(n_28978), .o(n_28980) );
no02f80 g540543 ( .a(n_27422), .b(x_in_10_15), .o(n_27423) );
no02f80 g540544 ( .a(n_28976), .b(n_29050), .o(n_28977) );
in01f80 g540545 ( .a(n_28092), .o(n_28093) );
na02f80 g540546 ( .a(n_27942), .b(x_in_48_14), .o(n_28092) );
no02f80 g540547 ( .a(n_27942), .b(x_in_48_14), .o(n_28266) );
no02f80 g540548 ( .a(n_28974), .b(n_28973), .o(n_28975) );
no02f80 g540549 ( .a(n_27418), .b(x_in_42_15), .o(n_27419) );
no02f80 g540550 ( .a(n_29094), .b(n_29093), .o(n_29095) );
no02f80 g540551 ( .a(n_28519), .b(n_28518), .o(n_28520) );
no02f80 g540552 ( .a(n_28971), .b(n_28970), .o(n_28972) );
no02f80 g540553 ( .a(n_27415), .b(x_in_26_15), .o(n_27416) );
no02f80 g540554 ( .a(n_28721), .b(n_28720), .o(n_28722) );
no02f80 g540555 ( .a(n_28968), .b(n_28967), .o(n_28969) );
no02f80 g540556 ( .a(n_27214), .b(n_27213), .o(n_27215) );
na02f80 g540557 ( .a(n_29073), .b(n_27457), .o(n_29249) );
in01f80 g540558 ( .a(n_28226), .o(n_28227) );
na02f80 g540559 ( .a(n_27746), .b(x_in_60_13), .o(n_28226) );
na02f80 g540560 ( .a(n_27745), .b(n_27562), .o(n_28265) );
in01f80 g540561 ( .a(n_27940), .o(n_27941) );
na02f80 g540562 ( .a(n_27361), .b(x_in_32_13), .o(n_27940) );
na02f80 g540563 ( .a(n_27360), .b(n_27151), .o(n_27995) );
in01f80 g540564 ( .a(n_28224), .o(n_28225) );
na02f80 g540565 ( .a(n_27737), .b(x_in_48_13), .o(n_28224) );
na02f80 g540566 ( .a(n_27736), .b(n_27547), .o(n_28264) );
na02f80 g540567 ( .a(n_27667), .b(x_in_52_13), .o(n_27406) );
na02f80 g540568 ( .a(n_27437), .b(FE_OFN290_n_27194), .o(n_27692) );
na02f80 g540569 ( .a(n_27402), .b(n_27624), .o(n_27403) );
na02f80 g540570 ( .a(n_27077), .b(n_27624), .o(n_27863) );
na02f80 g540571 ( .a(n_27939), .b(n_27829), .o(n_27797) );
na02f80 g540572 ( .a(n_27939), .b(n_27582), .o(n_28168) );
na02f80 g540573 ( .a(n_27386), .b(n_27160), .o(n_27986) );
na02f80 g540574 ( .a(n_27937), .b(FE_OFN1224_n_29433), .o(n_27938) );
no02f80 g540575 ( .a(n_28089), .b(n_29279), .o(n_28090) );
na02f80 g540576 ( .a(n_27795), .b(n_27794), .o(n_27796) );
na02f80 g540577 ( .a(n_27622), .b(n_27857), .o(n_27623) );
na02f80 g540578 ( .a(n_27936), .b(n_27792), .o(n_27793) );
na02f80 g540579 ( .a(n_27936), .b(n_27460), .o(n_28108) );
ao22s80 g540580 ( .a(n_27174), .b(n_26222), .c(x_out_42_32), .d(FE_OFN318_n_27400), .o(n_27401) );
no02f80 g540581 ( .a(n_27620), .b(n_27619), .o(n_27621) );
in01f80 g540582 ( .a(n_28104), .o(n_27618) );
na02f80 g540583 ( .a(FE_OFN945_n_27398), .b(n_27619), .o(n_28104) );
oa12f80 g540584 ( .a(n_28018), .b(n_27658), .c(n_28823), .o(n_29383) );
oa12f80 g540585 ( .a(n_27580), .b(n_27385), .c(n_26762), .o(n_27935) );
oa12f80 g540586 ( .a(n_27602), .b(n_28757), .c(n_27132), .o(n_29233) );
in01f80 g540587 ( .a(n_29327), .o(n_29248) );
oa12f80 g540588 ( .a(n_27766), .b(n_27302), .c(n_28840), .o(n_29327) );
in01f80 g540589 ( .a(n_29324), .o(n_29247) );
oa12f80 g540590 ( .a(n_27912), .b(n_27494), .c(n_28839), .o(n_29324) );
in01f80 g540591 ( .a(n_29321), .o(n_29246) );
oa12f80 g540592 ( .a(n_27601), .b(n_27127), .c(n_28838), .o(n_29321) );
in01f80 g540593 ( .a(n_29318), .o(n_29245) );
oa12f80 g540594 ( .a(n_27600), .b(n_27125), .c(n_28837), .o(n_29318) );
in01f80 g540595 ( .a(n_29228), .o(n_29166) );
oa12f80 g540596 ( .a(n_27765), .b(n_28756), .c(n_27296), .o(n_29228) );
in01f80 g540597 ( .a(n_29225), .o(n_29165) );
oa12f80 g540598 ( .a(n_27763), .b(n_28755), .c(n_27289), .o(n_29225) );
in01f80 g540599 ( .a(n_29155), .o(n_29092) );
oa12f80 g540600 ( .a(n_27764), .b(n_27294), .c(n_28659), .o(n_29155) );
in01f80 g540601 ( .a(n_29222), .o(n_29164) );
oa12f80 g540602 ( .a(n_27762), .b(n_28754), .c(n_27287), .o(n_29222) );
in01f80 g540603 ( .a(n_29219), .o(n_29163) );
oa12f80 g540604 ( .a(n_27599), .b(n_28753), .c(n_27119), .o(n_29219) );
in01f80 g540605 ( .a(n_29085), .o(n_28966) );
oa12f80 g540606 ( .a(n_27911), .b(n_27486), .c(n_28543), .o(n_29085) );
oa12f80 g540607 ( .a(n_26657), .b(n_26045), .c(n_28961), .o(n_29147) );
in01f80 g540608 ( .a(n_29162), .o(n_29381) );
oa12f80 g540609 ( .a(n_27761), .b(n_27284), .c(n_28751), .o(n_29162) );
in01f80 g540610 ( .a(n_29161), .o(n_29379) );
oa12f80 g540611 ( .a(n_27598), .b(n_27116), .c(n_28750), .o(n_29161) );
in01f80 g540612 ( .a(n_29244), .o(n_29451) );
oa12f80 g540613 ( .a(n_27382), .b(n_28836), .c(n_26907), .o(n_29244) );
oa12f80 g540614 ( .a(n_27381), .b(n_28835), .c(n_26905), .o(n_29298) );
in01f80 g540615 ( .a(n_28965), .o(n_29214) );
oa12f80 g540616 ( .a(n_27597), .b(n_27114), .c(n_28542), .o(n_28965) );
in01f80 g540617 ( .a(n_29160), .o(n_29377) );
oa12f80 g540618 ( .a(n_27595), .b(n_27110), .c(n_28749), .o(n_29160) );
in01f80 g540619 ( .a(n_29159), .o(n_29375) );
oa12f80 g540620 ( .a(n_27594), .b(n_27108), .c(n_28747), .o(n_29159) );
oa12f80 g540621 ( .a(n_27596), .b(n_28834), .c(n_27112), .o(n_29295) );
in01f80 g540622 ( .a(n_29158), .o(n_29373) );
oa12f80 g540623 ( .a(n_27593), .b(n_27106), .c(n_28746), .o(n_29158) );
oa12f80 g540624 ( .a(n_27182), .b(n_28833), .c(n_26676), .o(n_29292) );
oa12f80 g540625 ( .a(n_27181), .b(n_28657), .c(n_26598), .o(n_29144) );
oa12f80 g540626 ( .a(n_27180), .b(n_28832), .c(n_26596), .o(n_29289) );
oa12f80 g540627 ( .a(n_27760), .b(n_29036), .c(n_27280), .o(n_29434) );
oa12f80 g540628 ( .a(n_27592), .b(n_28744), .c(n_27103), .o(n_29202) );
oa12f80 g540629 ( .a(n_27179), .b(n_28831), .c(n_26594), .o(n_29286) );
oa12f80 g540630 ( .a(n_27178), .b(n_28829), .c(n_26589), .o(n_29283) );
oa12f80 g540631 ( .a(n_27591), .b(n_28743), .c(n_27101), .o(n_29199) );
oa12f80 g540632 ( .a(n_27590), .b(n_27099), .c(n_28433), .o(n_29074) );
oa12f80 g540633 ( .a(n_23241), .b(n_28956), .c(n_22586), .o(n_29141) );
in01f80 g540634 ( .a(n_29152), .o(n_29091) );
oa12f80 g540635 ( .a(n_27589), .b(n_27097), .c(n_28655), .o(n_29152) );
oa12f80 g540636 ( .a(n_27588), .b(n_28828), .c(n_27095), .o(n_29280) );
in01f80 g540637 ( .a(n_29081), .o(n_28964) );
oa12f80 g540638 ( .a(n_27759), .b(n_27277), .c(n_28541), .o(n_29081) );
oa12f80 g540639 ( .a(n_27394), .b(n_29079), .c(n_26941), .o(n_29196) );
in01f80 g540640 ( .a(n_29240), .o(n_29241) );
oa12f80 g540641 ( .a(n_27587), .b(n_28826), .c(n_27092), .o(n_29240) );
in01f80 g540642 ( .a(n_29238), .o(n_29239) );
oa12f80 g540643 ( .a(n_27586), .b(n_28825), .c(n_27090), .o(n_29238) );
oa12f80 g540644 ( .a(n_27170), .b(n_27367), .c(n_26112), .o(n_27615) );
in01f80 g540645 ( .a(n_29489), .o(n_29332) );
oa12f80 g540646 ( .a(n_28020), .b(n_28912), .c(n_27663), .o(n_29489) );
ao12f80 g540647 ( .a(n_28713), .b(n_28714), .c(n_27380), .o(n_28939) );
in01f80 g540648 ( .a(n_29236), .o(n_29237) );
oa12f80 g540649 ( .a(n_27585), .b(n_28824), .c(n_27088), .o(n_29236) );
in01f80 g540650 ( .a(n_28963), .o(n_29212) );
oa12f80 g540651 ( .a(n_27758), .b(n_28540), .c(n_27273), .o(n_28963) );
in01f80 g540652 ( .a(n_29090), .o(n_29308) );
oa12f80 g540653 ( .a(n_27362), .b(n_28951), .c(n_26890), .o(n_29090) );
oa12f80 g540654 ( .a(n_26640), .b(n_26026), .c(n_28949), .o(n_29138) );
in01f80 g540655 ( .a(n_27612), .o(n_28009) );
oa12f80 g540656 ( .a(n_12484), .b(n_27397), .c(n_13674), .o(n_27612) );
oa12f80 g540657 ( .a(n_27789), .b(n_1726), .c(FE_OFN364_n_4860), .o(n_27790) );
oa12f80 g540658 ( .a(n_27366), .b(n_27369), .c(n_26071), .o(n_27788) );
oa12f80 g540659 ( .a(n_27163), .b(n_27164), .c(n_26943), .o(n_27611) );
oa12f80 g540660 ( .a(n_27158), .b(n_1454), .c(FE_OFN100_n_27449), .o(n_27610) );
ao12f80 g540661 ( .a(n_24319), .b(n_28717), .c(n_24996), .o(n_28850) );
ao12f80 g540662 ( .a(n_26579), .b(n_28806), .c(n_27173), .o(n_29062) );
oa12f80 g540663 ( .a(n_27445), .b(n_29077), .c(n_27444), .o(n_29190) );
oa12f80 g540664 ( .a(n_27377), .b(n_27376), .c(n_29294), .o(n_29550) );
ao12f80 g540665 ( .a(n_27584), .b(n_27583), .c(n_29198), .o(n_29544) );
ao22s80 g540666 ( .a(n_28739), .b(n_27581), .c(n_29089), .d(x_in_60_13), .o(n_29314) );
ao12f80 g540667 ( .a(n_28865), .b(n_28864), .c(n_28863), .o(n_29088) );
ao22s80 g540668 ( .a(n_26976), .b(n_28961), .c(n_26975), .d(n_28658), .o(n_28962) );
oa12f80 g540669 ( .a(n_27193), .b(n_27195), .c(x_in_22_15), .o(n_29486) );
oa12f80 g540670 ( .a(n_26958), .b(n_26959), .c(x_in_54_15), .o(n_29483) );
oa12f80 g540671 ( .a(n_26956), .b(n_26957), .c(x_in_14_15), .o(n_29364) );
oa12f80 g540672 ( .a(n_26951), .b(n_26952), .c(x_in_46_15), .o(n_29480) );
oa12f80 g540673 ( .a(n_26949), .b(n_26950), .c(x_in_30_15), .o(n_29477) );
oa12f80 g540674 ( .a(n_26947), .b(n_26948), .c(x_in_62_15), .o(n_29474) );
ao12f80 g540675 ( .a(n_28803), .b(n_28802), .c(n_28801), .o(n_28958) );
oa22f80 g540676 ( .a(n_27395), .b(FE_OFN414_n_28303), .c(n_836), .d(FE_OFN115_n_27449), .o(n_27609) );
ao12f80 g540677 ( .a(n_28862), .b(n_28861), .c(n_28860), .o(n_29084) );
ao22s80 g540678 ( .a(n_28956), .b(n_23569), .c(n_28656), .d(n_23568), .o(n_28957) );
ao12f80 g540679 ( .a(n_27172), .b(n_27171), .c(n_29201), .o(n_29426) );
ao22s80 g540680 ( .a(n_28805), .b(x_in_32_13), .c(n_28432), .d(n_27159), .o(n_29075) );
ao22s80 g540681 ( .a(n_29079), .b(n_27604), .c(n_28742), .d(n_27603), .o(n_29080) );
ao12f80 g540682 ( .a(n_28634), .b(n_28717), .c(n_28633), .o(n_28804) );
ao12f80 g540683 ( .a(n_27375), .b(n_27374), .c(n_27373), .o(n_27784) );
in01f80 g540684 ( .a(n_27862), .o(n_27783) );
oa12f80 g540685 ( .a(n_27177), .b(n_27397), .c(n_27176), .o(n_27862) );
na03f80 g540686 ( .a(n_27395), .b(n_26561), .c(FE_OFN1113_rst), .o(n_27396) );
ao12f80 g540687 ( .a(n_28800), .b(n_28799), .c(n_28798), .o(n_28953) );
in01f80 g540688 ( .a(FE_OFN634_n_27731), .o(n_27717) );
ao22s80 g540689 ( .a(n_26261), .b(n_4062), .c(n_4063), .d(x_in_21_13), .o(n_27731) );
ao22s80 g540690 ( .a(n_29077), .b(n_27649), .c(n_29076), .d(n_27648), .o(n_29078) );
ao12f80 g540691 ( .a(n_28942), .b(n_28943), .c(n_28941), .o(n_29149) );
oa12f80 g540692 ( .a(n_27379), .b(n_28714), .c(n_28713), .o(n_28715) );
ao22s80 g540693 ( .a(n_28654), .b(n_27572), .c(n_28951), .d(n_27573), .o(n_28952) );
ao22s80 g540694 ( .a(n_26967), .b(n_28949), .c(n_26966), .d(n_28653), .o(n_28950) );
oa22f80 g540695 ( .a(n_28649), .b(FE_OFN400_n_28303), .c(n_1843), .d(FE_OFN347_n_4860), .o(n_28948) );
oa22f80 g540696 ( .a(n_28539), .b(FE_OFN400_n_28303), .c(n_40), .d(FE_OFN56_n_27012), .o(n_28871) );
oa22f80 g540697 ( .a(n_28537), .b(FE_OFN236_n_4162), .c(n_1498), .d(FE_OFN125_n_27449), .o(n_28870) );
oa22f80 g540698 ( .a(n_27035), .b(FE_OFN306_n_3069), .c(n_1745), .d(FE_OFN125_n_27449), .o(n_27776) );
oa22f80 g540699 ( .a(n_28341), .b(FE_OFN306_n_3069), .c(n_1445), .d(rst), .o(n_28712) );
oa22f80 g540700 ( .a(n_28647), .b(n_23291), .c(n_961), .d(FE_OFN1117_rst), .o(n_28945) );
oa22f80 g540701 ( .a(n_27254), .b(FE_OFN409_n_28303), .c(n_1975), .d(FE_OFN72_n_27012), .o(n_27913) );
oa22f80 g540702 ( .a(n_28535), .b(FE_OFN417_n_28303), .c(n_93), .d(FE_OFN108_n_27449), .o(n_28868) );
oa22f80 g540703 ( .a(n_28533), .b(FE_OFN312_n_3069), .c(n_1628), .d(FE_OFN113_n_27449), .o(n_28867) );
oa22f80 g540704 ( .a(n_28531), .b(FE_OFN296_n_3069), .c(n_1912), .d(FE_OFN108_n_27449), .o(n_28866) );
na02f80 g540733 ( .a(n_27385), .b(n_27205), .o(n_27386) );
no02f80 g540734 ( .a(n_28943), .b(x_in_36_14), .o(n_28944) );
na02f80 g540735 ( .a(n_27602), .b(n_27133), .o(n_28908) );
na02f80 g540736 ( .a(n_27766), .b(n_27303), .o(n_29018) );
na02f80 g540737 ( .a(n_27912), .b(n_27495), .o(n_29013) );
na02f80 g540738 ( .a(n_27601), .b(n_27128), .o(n_29010) );
na02f80 g540739 ( .a(n_27600), .b(n_27126), .o(n_29007) );
na02f80 g540740 ( .a(n_27765), .b(n_27297), .o(n_28905) );
na02f80 g540741 ( .a(n_27764), .b(n_27295), .o(n_28817) );
na02f80 g540742 ( .a(n_27763), .b(n_27290), .o(n_28902) );
na02f80 g540743 ( .a(n_27762), .b(n_27288), .o(n_28899) );
na02f80 g540744 ( .a(n_27599), .b(n_27120), .o(n_28896) );
na02f80 g540745 ( .a(n_27911), .b(n_27487), .o(n_28734) );
no02f80 g540746 ( .a(n_28864), .b(n_28863), .o(n_28865) );
na02f80 g540747 ( .a(n_27761), .b(n_27285), .o(n_28893) );
in01f80 g540748 ( .a(n_27383), .o(n_27384) );
no02f80 g540749 ( .a(n_27195), .b(x_in_22_14), .o(n_27383) );
na02f80 g540750 ( .a(n_27195), .b(x_in_22_14), .o(n_27814) );
na02f80 g540751 ( .a(n_27195), .b(x_in_22_15), .o(n_27193) );
na02f80 g540752 ( .a(n_27598), .b(n_27117), .o(n_28890) );
in01f80 g540753 ( .a(n_27191), .o(n_27192) );
no02f80 g540754 ( .a(n_26959), .b(x_in_54_14), .o(n_27191) );
na02f80 g540755 ( .a(n_26959), .b(x_in_54_14), .o(n_27635) );
na02f80 g540756 ( .a(n_26959), .b(x_in_54_15), .o(n_26958) );
na02f80 g540757 ( .a(n_27382), .b(n_26908), .o(n_29004) );
na02f80 g540758 ( .a(n_26906), .b(n_27381), .o(n_29001) );
na02f80 g540759 ( .a(n_27597), .b(n_27115), .o(n_28731) );
in01f80 g540760 ( .a(n_27189), .o(n_27190) );
no02f80 g540761 ( .a(n_26957), .b(x_in_14_14), .o(n_27189) );
na02f80 g540762 ( .a(n_26957), .b(x_in_14_14), .o(n_27634) );
na02f80 g540763 ( .a(n_26957), .b(x_in_14_15), .o(n_26956) );
na02f80 g540764 ( .a(n_27596), .b(n_27113), .o(n_28998) );
na02f80 g540765 ( .a(n_27595), .b(n_27111), .o(n_28887) );
in01f80 g540766 ( .a(n_27187), .o(n_27188) );
no02f80 g540767 ( .a(n_26952), .b(x_in_46_14), .o(n_27187) );
na02f80 g540768 ( .a(n_26952), .b(x_in_46_14), .o(n_27633) );
na02f80 g540769 ( .a(n_26952), .b(x_in_46_15), .o(n_26951) );
na02f80 g540770 ( .a(n_27594), .b(n_27109), .o(n_28884) );
in01f80 g540771 ( .a(n_27185), .o(n_27186) );
no02f80 g540772 ( .a(n_26950), .b(x_in_30_14), .o(n_27185) );
na02f80 g540773 ( .a(n_26950), .b(x_in_30_14), .o(n_27632) );
na02f80 g540774 ( .a(n_26950), .b(x_in_30_15), .o(n_26949) );
na02f80 g540775 ( .a(n_27593), .b(n_27107), .o(n_28881) );
na02f80 g540776 ( .a(n_26948), .b(x_in_62_14), .o(n_27631) );
in01f80 g540777 ( .a(n_27183), .o(n_27184) );
no02f80 g540778 ( .a(n_26948), .b(x_in_62_14), .o(n_27183) );
na02f80 g540779 ( .a(n_26948), .b(x_in_62_15), .o(n_26947) );
na02f80 g540780 ( .a(n_26677), .b(n_27182), .o(n_28995) );
no02f80 g540781 ( .a(n_28802), .b(n_28801), .o(n_28803) );
no02f80 g540782 ( .a(n_28861), .b(n_28860), .o(n_28862) );
no02f80 g540783 ( .a(n_28943), .b(n_28941), .o(n_28942) );
na02f80 g540784 ( .a(n_26599), .b(n_27181), .o(n_28811) );
na02f80 g540785 ( .a(n_27760), .b(n_27281), .o(n_29169) );
na02f80 g540786 ( .a(n_26597), .b(n_27180), .o(n_28992) );
na02f80 g540787 ( .a(n_27592), .b(n_27104), .o(n_28878) );
na02f80 g540788 ( .a(n_26595), .b(n_27179), .o(n_28989) );
na02f80 g540789 ( .a(n_27591), .b(n_27102), .o(n_28875) );
na02f80 g540790 ( .a(n_26590), .b(n_27178), .o(n_28986) );
na02f80 g540791 ( .a(n_27590), .b(n_27100), .o(n_28638) );
na02f80 g540792 ( .a(n_27589), .b(n_27098), .o(n_28808) );
in01f80 g540793 ( .a(n_28022), .o(n_28023) );
na02f80 g540794 ( .a(n_27910), .b(n_27483), .o(n_28022) );
na02f80 g540795 ( .a(n_27588), .b(n_27096), .o(n_28983) );
na02f80 g540796 ( .a(n_27759), .b(n_27278), .o(n_28726) );
no02f80 g540797 ( .a(n_28717), .b(n_28633), .o(n_28634) );
na02f80 g540798 ( .a(n_27397), .b(n_27176), .o(n_27177) );
na02f80 g540799 ( .a(n_27587), .b(n_27093), .o(n_28979) );
no02f80 g540800 ( .a(n_28799), .b(n_28798), .o(n_28800) );
na02f80 g540801 ( .a(n_27586), .b(n_27091), .o(n_28974) );
na02f80 g540802 ( .a(n_28020), .b(n_27664), .o(n_29094) );
na02f80 g540803 ( .a(n_27174), .b(n_26221), .o(n_27175) );
na02f80 g540804 ( .a(n_27380), .b(n_26875), .o(n_28519) );
no02f80 g540805 ( .a(n_26874), .b(x_in_52_13), .o(n_27379) );
na02f80 g540806 ( .a(n_27585), .b(n_27089), .o(n_28971) );
na02f80 g540807 ( .a(n_27758), .b(n_27274), .o(n_28721) );
na02f80 g540808 ( .a(n_28018), .b(n_27659), .o(n_28968) );
in01f80 g540809 ( .a(n_29072), .o(n_29073) );
no02f80 g540810 ( .a(n_29077), .b(n_26962), .o(n_29072) );
in01f80 g540811 ( .a(n_27908), .o(n_27909) );
na02f80 g540812 ( .a(n_27272), .b(n_27757), .o(n_27908) );
na02f80 g540813 ( .a(n_26578), .b(n_27173), .o(n_28728) );
na02f80 g540814 ( .a(n_26817), .b(FE_OFN1181_rst), .o(n_27789) );
na02f80 g540815 ( .a(n_27376), .b(n_29294), .o(n_27377) );
no02f80 g540816 ( .a(n_27583), .b(n_29198), .o(n_27584) );
ao22s80 g540817 ( .a(n_26215), .b(n_11072), .c(n_25730), .d(n_12422), .o(n_27430) );
oa12f80 g540818 ( .a(n_27754), .b(n_44), .c(FE_OFN1123_rst), .o(n_27756) );
oa12f80 g540819 ( .a(n_27754), .b(n_959), .c(FE_OFN78_n_27012), .o(n_27755) );
oa12f80 g540820 ( .a(n_27754), .b(n_1181), .c(FE_OFN78_n_27012), .o(n_27753) );
no02f80 g540821 ( .a(n_27171), .b(n_29201), .o(n_27172) );
oa12f80 g540822 ( .a(n_27904), .b(n_1816), .c(FE_OFN116_n_27449), .o(n_27907) );
oa12f80 g540823 ( .a(n_27904), .b(n_167), .c(FE_OFN353_n_4860), .o(n_27905) );
oa12f80 g540824 ( .a(n_27904), .b(n_207), .c(FE_OFN116_n_27449), .o(n_27903) );
oa12f80 g540825 ( .a(n_27904), .b(n_440), .c(FE_OFN116_n_27449), .o(n_27901) );
no02f80 g540826 ( .a(n_27374), .b(n_27373), .o(n_27375) );
no02f80 g540827 ( .a(n_27374), .b(n_27006), .o(n_28400) );
ao22s80 g540828 ( .a(n_26582), .b(n_26225), .c(x_out_41_32), .d(FE_OFN271_n_16028), .o(n_27170) );
in01f80 g540829 ( .a(n_27829), .o(n_27582) );
na02f80 g540830 ( .a(n_26872), .b(n_26515), .o(n_27829) );
oa12f80 g540831 ( .a(n_27385), .b(n_1800), .c(FE_OFN119_n_27449), .o(n_27372) );
oa12f80 g540832 ( .a(n_3247), .b(n_28628), .c(n_2196), .o(n_28814) );
in01f80 g540833 ( .a(n_28709), .o(n_28932) );
oa12f80 g540834 ( .a(n_27443), .b(n_27203), .c(n_28623), .o(n_28709) );
oa12f80 g540835 ( .a(n_28029), .b(n_28856), .c(n_27743), .o(n_29097) );
in01f80 g540836 ( .a(n_28859), .o(n_29117) );
oa12f80 g540837 ( .a(n_27364), .b(n_28781), .c(n_26921), .o(n_28859) );
ao12f80 g540838 ( .a(n_28776), .b(n_27246), .c(n_28778), .o(n_29050) );
oa12f80 g540839 ( .a(n_27750), .b(n_428), .c(FE_OFN131_n_27449), .o(n_27752) );
oa12f80 g540840 ( .a(n_27750), .b(n_1283), .c(FE_OFN361_n_4860), .o(n_27751) );
oa12f80 g540841 ( .a(n_27750), .b(n_509), .c(FE_OFN131_n_27449), .o(n_27749) );
oa12f80 g540842 ( .a(n_27894), .b(n_1308), .c(FE_OFN353_n_4860), .o(n_27897) );
oa12f80 g540843 ( .a(n_27894), .b(n_1288), .c(FE_OFN353_n_4860), .o(n_27895) );
oa12f80 g540844 ( .a(n_27894), .b(n_1719), .c(FE_OFN353_n_4860), .o(n_27893) );
oa12f80 g540845 ( .a(n_27894), .b(n_1536), .c(FE_OFN353_n_4860), .o(n_27892) );
oa12f80 g540846 ( .a(n_27369), .b(n_355), .c(FE_OFN353_n_4860), .o(n_27370) );
oa12f80 g540847 ( .a(n_27164), .b(n_256), .c(FE_OFN1114_rst), .o(n_27165) );
oa12f80 g540848 ( .a(n_27367), .b(n_698), .c(FE_OFN1120_rst), .o(n_27368) );
ao22s80 g540849 ( .a(n_26560), .b(n_26761), .c(x_out_39_32), .d(FE_OFN279_n_16656), .o(n_27366) );
ao22s80 g540850 ( .a(n_26517), .b(n_26191), .c(x_out_40_32), .d(FE_OFN318_n_27400), .o(n_27163) );
oa12f80 g540851 ( .a(n_11939), .b(n_26619), .c(n_13180), .o(n_27214) );
ao12f80 g540852 ( .a(x_in_41_15), .b(n_27162), .c(n_27161), .o(n_27630) );
oa12f80 g540853 ( .a(FE_OFN1114_rst), .b(n_26576), .c(n_26943), .o(n_26945) );
in01f80 g540854 ( .a(n_27437), .o(n_27160) );
ao12f80 g540855 ( .a(n_14082), .b(n_26218), .c(n_12822), .o(n_27437) );
in01f80 g540856 ( .a(n_27745), .o(n_27746) );
ao12f80 g540857 ( .a(n_27083), .b(n_27581), .c(n_27082), .o(n_27745) );
ao12f80 g540858 ( .a(n_28475), .b(n_28474), .c(n_28473), .o(n_28707) );
ao12f80 g540859 ( .a(n_27206), .b(x_out_47_31), .c(n_16656), .o(n_27580) );
oa12f80 g540860 ( .a(n_26278), .b(n_26277), .c(n_26276), .o(n_27435) );
ao12f80 g540861 ( .a(n_28591), .b(n_28590), .c(n_28589), .o(n_28795) );
ao12f80 g540862 ( .a(n_28594), .b(n_28593), .c(n_28592), .o(n_28794) );
oa12f80 g540863 ( .a(n_26575), .b(n_26574), .c(n_26868), .o(n_27642) );
ao12f80 g540864 ( .a(n_28588), .b(n_28587), .c(n_28586), .o(n_28793) );
oa12f80 g540865 ( .a(n_26867), .b(n_26866), .c(n_27078), .o(n_27826) );
ao12f80 g540866 ( .a(n_28767), .b(n_28766), .c(FE_OFN492_n_28765), .o(n_28940) );
ao12f80 g540867 ( .a(n_28585), .b(n_28584), .c(n_28583), .o(n_28792) );
oa12f80 g540868 ( .a(n_26865), .b(n_26864), .c(n_26863), .o(n_27825) );
ao12f80 g540869 ( .a(n_28582), .b(n_28581), .c(n_28580), .o(n_28791) );
oa12f80 g540870 ( .a(n_26862), .b(n_26861), .c(n_26860), .o(n_27824) );
ao12f80 g540871 ( .a(n_28472), .b(n_28471), .c(n_28470), .o(n_28706) );
oa12f80 g540872 ( .a(n_26573), .b(n_26572), .c(n_26859), .o(n_27638) );
ao12f80 g540873 ( .a(n_28353), .b(n_28352), .c(n_28351), .o(n_28630) );
ao12f80 g540874 ( .a(n_28469), .b(n_28468), .c(n_28467), .o(n_28705) );
in01f80 g540875 ( .a(n_27622), .o(n_27821) );
ao12f80 g540876 ( .a(n_26587), .b(n_26586), .c(n_26585), .o(n_27622) );
oa12f80 g540877 ( .a(n_26571), .b(n_26570), .c(n_26858), .o(n_27637) );
na03f80 g540878 ( .a(n_15850), .b(n_26584), .c(n_11046), .o(n_27795) );
ao12f80 g540879 ( .a(n_28466), .b(n_28465), .c(n_28464), .o(n_28704) );
oa12f80 g540880 ( .a(n_26569), .b(n_26568), .c(n_26857), .o(n_27636) );
ao12f80 g540881 ( .a(n_28463), .b(n_28462), .c(n_28461), .o(n_28703) );
oa12f80 g540882 ( .a(n_26856), .b(n_26855), .c(n_26854), .o(n_27816) );
ao12f80 g540883 ( .a(n_28257), .b(n_28256), .c(n_28255), .o(n_28493) );
oa12f80 g540884 ( .a(n_26853), .b(n_26852), .c(n_26851), .o(n_27815) );
ao12f80 g540885 ( .a(n_28460), .b(n_28459), .c(n_28458), .o(n_28702) );
ao12f80 g540886 ( .a(n_28457), .b(n_28456), .c(n_28455), .o(n_28701) );
ao12f80 g540887 ( .a(n_28579), .b(n_28578), .c(n_28577), .o(n_28790) );
ao12f80 g540888 ( .a(n_28576), .b(n_28575), .c(n_28574), .o(n_28789) );
ao12f80 g540889 ( .a(n_28250), .b(n_28249), .c(n_28248), .o(n_28492) );
ao12f80 g540890 ( .a(n_28573), .b(n_28572), .c(n_28571), .o(n_28788) );
oa12f80 g540891 ( .a(n_26600), .b(n_26743), .c(x_in_22_15), .o(n_29297) );
ao12f80 g540892 ( .a(n_28253), .b(n_28252), .c(n_28251), .o(n_28491) );
ao12f80 g540893 ( .a(n_28454), .b(n_28453), .c(n_28452), .o(n_28700) );
ao12f80 g540894 ( .a(n_28451), .b(n_28450), .c(n_28449), .o(n_28699) );
ao12f80 g540895 ( .a(n_28448), .b(n_28447), .c(n_28446), .o(n_28698) );
ao12f80 g540896 ( .a(n_28570), .b(n_28569), .c(n_28568), .o(n_28787) );
oa12f80 g540897 ( .a(n_26301), .b(n_26302), .c(x_in_54_15), .o(n_29291) );
ao22s80 g540898 ( .a(n_28628), .b(n_4051), .c(n_28339), .d(n_4050), .o(n_28629) );
ao12f80 g540899 ( .a(n_28445), .b(n_28444), .c(n_28525), .o(n_28697) );
ao12f80 g540900 ( .a(n_28350), .b(n_28349), .c(n_28348), .o(n_28627) );
oa12f80 g540901 ( .a(n_26299), .b(n_26300), .c(x_in_14_15), .o(n_29143) );
ao12f80 g540902 ( .a(n_28762), .b(n_28761), .c(n_28760), .o(n_28938) );
ao12f80 g540903 ( .a(n_28567), .b(n_28566), .c(n_28565), .o(n_28786) );
oa12f80 g540904 ( .a(n_26297), .b(n_26298), .c(x_in_46_15), .o(n_29288) );
in01f80 g540905 ( .a(FE_OFN945_n_27398), .o(n_27620) );
ao12f80 g540906 ( .a(n_26281), .b(n_26619), .c(n_26280), .o(n_27398) );
ao12f80 g540907 ( .a(n_28443), .b(n_28442), .c(n_28441), .o(n_28696) );
ao12f80 g540908 ( .a(n_28564), .b(n_28563), .c(n_28562), .o(n_28785) );
oa12f80 g540909 ( .a(n_26295), .b(n_26296), .c(x_in_30_15), .o(n_29285) );
ao12f80 g540910 ( .a(n_28440), .b(n_28439), .c(n_28438), .o(n_28695) );
ao12f80 g540911 ( .a(n_28561), .b(n_28560), .c(n_28559), .o(n_28784) );
oa12f80 g540912 ( .a(n_26293), .b(n_26294), .c(x_in_62_15), .o(n_29282) );
ao12f80 g540913 ( .a(n_28347), .b(n_28346), .c(n_28345), .o(n_28626) );
ao12f80 g540914 ( .a(n_28103), .b(n_28102), .c(n_28101), .o(n_28369) );
in01f80 g540915 ( .a(n_27360), .o(n_27361) );
ao12f80 g540916 ( .a(n_26567), .b(n_27159), .c(n_26848), .o(n_27360) );
ao12f80 g540917 ( .a(n_28344), .b(n_28343), .c(n_28342), .o(n_28625) );
oa12f80 g540918 ( .a(n_26846), .b(n_26845), .c(n_26844), .o(n_27803) );
ao22s80 g540919 ( .a(n_27646), .b(n_28623), .c(n_27645), .d(n_28338), .o(n_28624) );
ao12f80 g540920 ( .a(n_28558), .b(n_28557), .c(n_28556), .o(n_28783) );
in01f80 g540921 ( .a(n_27736), .o(n_27737) );
ao12f80 g540922 ( .a(n_27075), .b(n_27570), .c(n_27262), .o(n_27736) );
in01f80 g540923 ( .a(n_27936), .o(n_27942) );
ao12f80 g540924 ( .a(n_26871), .b(n_26870), .c(n_26869), .o(n_27936) );
ao22s80 g540925 ( .a(n_28158), .b(n_28856), .c(n_28157), .d(n_28643), .o(n_28857) );
ao12f80 g540926 ( .a(n_28245), .b(n_28244), .c(n_28243), .o(n_28490) );
oa22f80 g540927 ( .a(n_26631), .b(n_27161), .c(n_27162), .d(n_26605), .o(n_27802) );
ao12f80 g540928 ( .a(n_28242), .b(n_28241), .c(n_28240), .o(n_28489) );
ao22s80 g540929 ( .a(n_28524), .b(n_27576), .c(n_28781), .d(n_27577), .o(n_28782) );
ao12f80 g540930 ( .a(n_28555), .b(n_28554), .c(n_28553), .o(n_28780) );
oa12f80 g540931 ( .a(n_26275), .b(n_26274), .c(n_26273), .o(n_27422) );
ao22s80 g540932 ( .a(n_27442), .b(n_28778), .c(n_27441), .d(n_28523), .o(n_28779) );
oa12f80 g540933 ( .a(n_27245), .b(n_28776), .c(n_28778), .o(n_28777) );
in01f80 g540934 ( .a(n_26927), .o(n_26928) );
oa22f80 g540935 ( .a(n_25968), .b(n_15752), .c(n_4151), .d(x_in_5_15), .o(n_26927) );
ao12f80 g540936 ( .a(n_28552), .b(n_28551), .c(n_28550), .o(n_28775) );
ao12f80 g540937 ( .a(n_28665), .b(n_28664), .c(n_28663), .o(n_28855) );
oa12f80 g540938 ( .a(n_26272), .b(n_26271), .c(n_26270), .o(n_27418) );
ao12f80 g540939 ( .a(n_28437), .b(n_28436), .c(n_28435), .o(n_28694) );
na03f80 g540940 ( .a(n_26583), .b(n_27231), .c(FE_OFN1120_rst), .o(n_27158) );
ao12f80 g540941 ( .a(n_28662), .b(n_28661), .c(n_28660), .o(n_28854) );
ao12f80 g540942 ( .a(n_27970), .b(n_27969), .c(n_27968), .o(n_28267) );
oa12f80 g540943 ( .a(n_26269), .b(n_26279), .c(n_26926), .o(n_27667) );
ao12f80 g540944 ( .a(n_28549), .b(n_28548), .c(n_28547), .o(n_28774) );
ao12f80 g540945 ( .a(n_26558), .b(n_26557), .c(n_26556), .o(n_27157) );
oa12f80 g540946 ( .a(n_26268), .b(n_26267), .c(n_26266), .o(n_27415) );
ao12f80 g540947 ( .a(n_28238), .b(n_28237), .c(n_28236), .o(n_28488) );
oa12f80 g540948 ( .a(n_27084), .b(n_27086), .c(x_in_12_15), .o(n_29361) );
ao12f80 g540949 ( .a(n_28546), .b(n_28545), .c(n_28544), .o(n_28773) );
oa22f80 g540950 ( .a(n_26998), .b(FE_OFN251_n_4162), .c(n_628), .d(FE_OFN1111_rst), .o(n_27566) );
oa22f80 g540951 ( .a(n_28421), .b(FE_OFN251_n_4162), .c(n_220), .d(FE_OFN65_n_27012), .o(n_28693) );
oa22f80 g540952 ( .a(n_28420), .b(FE_OFN247_n_4162), .c(n_1795), .d(FE_OFN69_n_27012), .o(n_28691) );
oa22f80 g540953 ( .a(n_27581), .b(x_in_60_13), .c(n_26997), .d(n_27562), .o(n_29015) );
oa22f80 g540954 ( .a(n_28419), .b(FE_OFN417_n_28303), .c(n_1621), .d(FE_OFN361_n_4860), .o(n_28690) );
oa22f80 g540955 ( .a(n_28642), .b(FE_OFN234_n_4162), .c(n_1667), .d(FE_OFN360_n_4860), .o(n_28853) );
oa22f80 g540956 ( .a(n_28418), .b(FE_OFN417_n_28303), .c(n_427), .d(FE_OFN361_n_4860), .o(n_28689) );
oa22f80 g540957 ( .a(n_28417), .b(FE_OFN308_n_3069), .c(n_10), .d(FE_OFN90_n_27449), .o(n_28687) );
oa22f80 g540958 ( .a(n_28233), .b(n_28771), .c(n_1542), .d(FE_OFN358_n_4860), .o(n_28485) );
oa22f80 g540959 ( .a(n_28337), .b(FE_OFN299_n_3069), .c(n_1377), .d(FE_OFN350_n_4860), .o(n_28622) );
oa22f80 g540960 ( .a(n_28336), .b(FE_OFN308_n_3069), .c(n_876), .d(FE_OFN326_n_4860), .o(n_28619) );
oa22f80 g540961 ( .a(n_28335), .b(FE_OFN294_n_3069), .c(n_1777), .d(FE_OFN331_n_4860), .o(n_28617) );
oa22f80 g540962 ( .a(n_28334), .b(FE_OFN300_n_3069), .c(n_1864), .d(FE_OFN91_n_27449), .o(n_28616) );
oa22f80 g540963 ( .a(n_28098), .b(FE_OFN296_n_3069), .c(n_649), .d(FE_OFN1117_rst), .o(n_28368) );
oa22f80 g540964 ( .a(n_28333), .b(FE_OFN294_n_3069), .c(n_1931), .d(FE_OFN133_n_27449), .o(n_28614) );
oa22f80 g540965 ( .a(n_28415), .b(FE_OFN309_n_3069), .c(n_1929), .d(FE_OFN134_n_27449), .o(n_28686) );
oa22f80 g540966 ( .a(n_28332), .b(n_21988), .c(n_186), .d(FE_OFN68_n_27012), .o(n_28613) );
oa22f80 g540967 ( .a(n_28416), .b(n_28682), .c(n_235), .d(FE_OFN1106_rst), .o(n_28684) );
oa22f80 g540968 ( .a(n_28414), .b(n_28682), .c(n_1039), .d(FE_OFN363_n_4860), .o(n_28683) );
oa22f80 g540969 ( .a(n_28097), .b(FE_OFN409_n_28303), .c(n_770), .d(FE_OFN355_n_4860), .o(n_28367) );
oa22f80 g540970 ( .a(n_28096), .b(FE_OFN234_n_4162), .c(n_1267), .d(FE_OFN76_n_27012), .o(n_28366) );
oa22f80 g540971 ( .a(n_28331), .b(FE_OFN405_n_28303), .c(n_500), .d(FE_OFN94_n_27449), .o(n_28612) );
oa22f80 g540972 ( .a(n_28330), .b(FE_OFN4_n_28682), .c(n_1687), .d(FE_OFN56_n_27012), .o(n_28611) );
oa22f80 g540973 ( .a(n_28329), .b(n_28608), .c(n_853), .d(n_28607), .o(n_28609) );
oa22f80 g540974 ( .a(n_28413), .b(FE_OFN297_n_3069), .c(n_1043), .d(FE_OFN352_n_4860), .o(n_28681) );
oa22f80 g540975 ( .a(FE_OFN1011_n_28328), .b(n_28608), .c(n_1226), .d(FE_OFN336_n_4860), .o(n_28606) );
oa22f80 g540976 ( .a(n_28327), .b(FE_OFN294_n_3069), .c(n_187), .d(FE_OFN68_n_27012), .o(n_28604) );
oa22f80 g540977 ( .a(n_28232), .b(FE_OFN307_n_3069), .c(n_1971), .d(FE_OFN1112_rst), .o(n_28484) );
oa22f80 g540978 ( .a(n_28640), .b(FE_OFN417_n_28303), .c(n_965), .d(FE_OFN361_n_4860), .o(n_28848) );
oa22f80 g540979 ( .a(n_28412), .b(n_29033), .c(n_814), .d(FE_OFN324_n_4860), .o(n_28680) );
oa22f80 g540980 ( .a(n_26467), .b(n_29033), .c(n_1399), .d(FE_OFN1115_rst), .o(n_27154) );
oa22f80 g540981 ( .a(n_28326), .b(n_28682), .c(n_1289), .d(FE_OFN1121_rst), .o(n_28602) );
oa22f80 g540982 ( .a(n_28411), .b(FE_OFN303_n_3069), .c(n_353), .d(FE_OFN114_n_27449), .o(n_28679) );
oa22f80 g540983 ( .a(n_28325), .b(FE_OFN3_n_28682), .c(n_1792), .d(FE_OFN131_n_27449), .o(n_28601) );
oa22f80 g540984 ( .a(n_28410), .b(n_28682), .c(n_228), .d(n_27449), .o(n_28678) );
oa22f80 g540985 ( .a(n_28231), .b(FE_OFN4_n_28682), .c(n_305), .d(FE_OFN115_n_27449), .o(n_28481) );
oa22f80 g540986 ( .a(n_27945), .b(FE_OFN296_n_3069), .c(n_999), .d(FE_OFN131_n_27449), .o(n_28263) );
oa22f80 g540987 ( .a(n_28230), .b(FE_OFN294_n_3069), .c(n_1127), .d(FE_OFN138_n_27449), .o(n_28480) );
oa22f80 g540988 ( .a(FE_OFN913_n_28409), .b(n_29033), .c(n_1871), .d(FE_OFN63_n_27012), .o(n_28677) );
oa22f80 g540989 ( .a(FE_OFN879_n_28229), .b(n_29033), .c(n_1342), .d(FE_OFN63_n_27012), .o(n_28478) );
oa22f80 g540990 ( .a(n_28522), .b(FE_OFN203_n_28771), .c(n_1273), .d(FE_OFN130_n_27449), .o(n_28772) );
oa22f80 g540991 ( .a(n_28095), .b(FE_OFN312_n_3069), .c(n_1429), .d(FE_OFN64_n_27012), .o(n_28365) );
oa22f80 g540992 ( .a(n_28094), .b(FE_OFN296_n_3069), .c(n_1455), .d(n_28362), .o(n_28363) );
oa22f80 g540993 ( .a(n_27159), .b(x_in_32_13), .c(n_26849), .d(n_27151), .o(n_28723) );
oa22f80 g540994 ( .a(FE_OFN516_n_28406), .b(n_4280), .c(n_1503), .d(n_28362), .o(n_28674) );
oa22f80 g540995 ( .a(n_28408), .b(FE_OFN265_n_4280), .c(n_1540), .d(FE_OFN1143_n_27012), .o(n_28673) );
oa22f80 g540996 ( .a(n_26702), .b(FE_OFN265_n_4280), .c(n_777), .d(FE_OFN353_n_4860), .o(n_27346) );
oa22f80 g540997 ( .a(FE_OFN885_n_28405), .b(n_28608), .c(n_1153), .d(FE_OFN1108_rst), .o(n_28672) );
oa22f80 g540998 ( .a(n_27570), .b(x_in_48_13), .c(n_27263), .d(n_27547), .o(n_28976) );
oa22f80 g540999 ( .a(n_26463), .b(n_28608), .c(n_309), .d(FE_OFN190_n_28362), .o(n_27148) );
oa22f80 g541000 ( .a(n_28403), .b(FE_OFN248_n_4162), .c(n_163), .d(FE_OFN326_n_4860), .o(n_28670) );
oa22f80 g541001 ( .a(n_28323), .b(n_28597), .c(n_1440), .d(FE_OFN363_n_4860), .o(n_28598) );
oa22f80 g541002 ( .a(n_28517), .b(FE_OFN7_n_28597), .c(n_433), .d(FE_OFN1146_n_4860), .o(n_28770) );
oa22f80 g541003 ( .a(FE_OFN773_n_26698), .b(n_29033), .c(n_1357), .d(FE_OFN349_n_4860), .o(n_27344) );
oa22f80 g541004 ( .a(n_28516), .b(FE_OFN247_n_4162), .c(n_1313), .d(FE_OFN134_n_27449), .o(n_28769) );
oa22f80 g541005 ( .a(FE_OFN626_n_26697), .b(n_29033), .c(n_1158), .d(FE_OFN1108_rst), .o(n_27343) );
oa22f80 g541006 ( .a(n_27798), .b(FE_OFN7_n_28597), .c(n_1231), .d(FE_OFN130_n_27449), .o(n_28107) );
oa22f80 g541007 ( .a(n_28402), .b(FE_OFN214_n_29687), .c(n_405), .d(FE_OFN78_n_27012), .o(n_28669) );
oa22f80 g541008 ( .a(n_26695), .b(FE_OFN259_n_4280), .c(n_598), .d(FE_OFN1119_rst), .o(n_27341) );
oa22f80 g541009 ( .a(n_28091), .b(FE_OFN217_n_29687), .c(n_155), .d(FE_OFN1113_rst), .o(n_28359) );
oa22f80 g541010 ( .a(n_28322), .b(FE_OFN248_n_4162), .c(n_1518), .d(FE_OFN326_n_4860), .o(n_28595) );
oa22f80 g541011 ( .a(n_28399), .b(FE_OFN251_n_4162), .c(n_483), .d(rst), .o(n_28668) );
oa22f80 g541012 ( .a(n_27473), .b(x_in_50_15), .c(n_27474), .d(n_2), .o(n_29279) );
oa22f80 g541013 ( .a(n_27270), .b(n_1125), .c(n_27269), .d(x_in_34_15), .o(n_29433) );
in01f80 g541014 ( .a(n_27624), .o(n_27426) );
ao22s80 g541015 ( .a(n_25965), .b(n_4984), .c(n_13928), .d(x_in_33_14), .o(n_27624) );
no02f80 g541090 ( .a(n_26909), .b(n_27205), .o(n_27206) );
na02f80 g541091 ( .a(n_26909), .b(FE_OFN34_n_15183), .o(n_27385) );
na02f80 g541092 ( .a(n_26605), .b(x_in_40_13), .o(n_27382) );
in01f80 g541093 ( .a(n_26907), .o(n_26908) );
no02f80 g541094 ( .a(n_26605), .b(x_in_40_13), .o(n_26907) );
in01f80 g541095 ( .a(n_26905), .o(n_26906) );
no02f80 g541096 ( .a(n_26743), .b(x_in_22_14), .o(n_26905) );
na02f80 g541097 ( .a(n_26743), .b(x_in_22_14), .o(n_27381) );
na02f80 g541098 ( .a(n_26743), .b(x_in_22_15), .o(n_26600) );
na02f80 g541099 ( .a(n_26302), .b(x_in_54_14), .o(n_27182) );
in01f80 g541100 ( .a(n_26676), .o(n_26677) );
no02f80 g541101 ( .a(n_26302), .b(x_in_54_14), .o(n_26676) );
na02f80 g541102 ( .a(n_26302), .b(x_in_54_15), .o(n_26301) );
in01f80 g541103 ( .a(n_26598), .o(n_26599) );
no02f80 g541104 ( .a(n_26300), .b(x_in_14_14), .o(n_26598) );
na02f80 g541105 ( .a(n_26300), .b(x_in_14_14), .o(n_27181) );
na02f80 g541106 ( .a(n_26300), .b(x_in_14_15), .o(n_26299) );
in01f80 g541107 ( .a(n_26596), .o(n_26597) );
no02f80 g541108 ( .a(n_26298), .b(x_in_46_14), .o(n_26596) );
na02f80 g541109 ( .a(n_26298), .b(x_in_46_14), .o(n_27180) );
na02f80 g541110 ( .a(n_26298), .b(x_in_46_15), .o(n_26297) );
in01f80 g541111 ( .a(n_26594), .o(n_26595) );
no02f80 g541112 ( .a(n_26296), .b(x_in_30_14), .o(n_26594) );
na02f80 g541113 ( .a(n_26296), .b(x_in_30_14), .o(n_27179) );
na02f80 g541114 ( .a(n_26296), .b(x_in_30_15), .o(n_26295) );
in01f80 g541115 ( .a(n_26589), .o(n_26590) );
no02f80 g541116 ( .a(n_26294), .b(x_in_62_14), .o(n_26589) );
na02f80 g541117 ( .a(n_26294), .b(x_in_62_14), .o(n_27178) );
na02f80 g541118 ( .a(n_26294), .b(x_in_62_15), .o(n_26293) );
no02f80 g541119 ( .a(n_28474), .b(n_28473), .o(n_28475) );
na02f80 g541120 ( .a(n_26901), .b(x_in_58_14), .o(n_27602) );
in01f80 g541121 ( .a(n_27132), .o(n_27133) );
no02f80 g541122 ( .a(n_26901), .b(x_in_58_14), .o(n_27132) );
no02f80 g541123 ( .a(n_28593), .b(n_28592), .o(n_28594) );
na02f80 g541124 ( .a(n_27129), .b(x_in_2_13), .o(n_27766) );
in01f80 g541125 ( .a(n_27302), .o(n_27303) );
no02f80 g541126 ( .a(n_27129), .b(x_in_2_13), .o(n_27302) );
no02f80 g541127 ( .a(n_28590), .b(n_28589), .o(n_28591) );
no02f80 g541128 ( .a(n_28587), .b(n_28586), .o(n_28588) );
na02f80 g541129 ( .a(n_27301), .b(x_in_34_13), .o(n_27912) );
in01f80 g541130 ( .a(n_27494), .o(n_27495) );
no02f80 g541131 ( .a(n_27301), .b(x_in_34_13), .o(n_27494) );
no02f80 g541132 ( .a(n_28766), .b(FE_OFN492_n_28765), .o(n_28767) );
no02f80 g541133 ( .a(n_28584), .b(n_28583), .o(n_28585) );
na02f80 g541134 ( .a(n_26896), .b(x_in_18_13), .o(n_27601) );
in01f80 g541135 ( .a(n_27127), .o(n_27128) );
no02f80 g541136 ( .a(n_26896), .b(x_in_18_13), .o(n_27127) );
no02f80 g541137 ( .a(n_28581), .b(n_28580), .o(n_28582) );
na02f80 g541138 ( .a(n_26895), .b(x_in_50_13), .o(n_27600) );
in01f80 g541139 ( .a(n_27125), .o(n_27126) );
no02f80 g541140 ( .a(n_26895), .b(x_in_50_13), .o(n_27125) );
no02f80 g541141 ( .a(n_28471), .b(n_28470), .o(n_28472) );
na02f80 g541142 ( .a(n_27124), .b(x_in_10_13), .o(n_27765) );
in01f80 g541143 ( .a(n_27296), .o(n_27297) );
no02f80 g541144 ( .a(n_27124), .b(x_in_10_13), .o(n_27296) );
no02f80 g541145 ( .a(n_28352), .b(n_28351), .o(n_28353) );
na02f80 g541146 ( .a(n_27123), .b(x_in_6_13), .o(n_27764) );
in01f80 g541147 ( .a(n_27294), .o(n_27295) );
no02f80 g541148 ( .a(n_27123), .b(x_in_6_13), .o(n_27294) );
no02f80 g541149 ( .a(n_28468), .b(n_28467), .o(n_28469) );
na02f80 g541150 ( .a(n_27122), .b(x_in_42_13), .o(n_27763) );
in01f80 g541151 ( .a(n_27289), .o(n_27290) );
no02f80 g541152 ( .a(n_27122), .b(x_in_42_13), .o(n_27289) );
no02f80 g541153 ( .a(n_26586), .b(n_26585), .o(n_26587) );
na02f80 g541154 ( .a(n_26586), .b(n_15849), .o(n_26584) );
no02f80 g541155 ( .a(n_28465), .b(n_28464), .o(n_28466) );
na02f80 g541156 ( .a(n_27121), .b(x_in_26_13), .o(n_27762) );
in01f80 g541157 ( .a(n_27287), .o(n_27288) );
no02f80 g541158 ( .a(n_27121), .b(x_in_26_13), .o(n_27287) );
no02f80 g541159 ( .a(n_28462), .b(n_28461), .o(n_28463) );
na02f80 g541160 ( .a(n_26889), .b(x_in_58_13), .o(n_27599) );
in01f80 g541161 ( .a(n_27119), .o(n_27120) );
no02f80 g541162 ( .a(n_26889), .b(x_in_58_13), .o(n_27119) );
no02f80 g541163 ( .a(n_28256), .b(n_28255), .o(n_28257) );
na02f80 g541164 ( .a(n_27286), .b(x_in_6_12), .o(n_27911) );
in01f80 g541165 ( .a(n_27486), .o(n_27487) );
no02f80 g541166 ( .a(n_27286), .b(x_in_6_12), .o(n_27486) );
no02f80 g541167 ( .a(n_28459), .b(n_28458), .o(n_28460) );
na02f80 g541168 ( .a(n_27118), .b(x_in_22_13), .o(n_27761) );
in01f80 g541169 ( .a(n_27284), .o(n_27285) );
no02f80 g541170 ( .a(n_27118), .b(x_in_22_13), .o(n_27284) );
no02f80 g541171 ( .a(n_28456), .b(n_28455), .o(n_28457) );
na02f80 g541172 ( .a(n_26888), .b(x_in_54_13), .o(n_27598) );
in01f80 g541173 ( .a(n_27116), .o(n_27117) );
no02f80 g541174 ( .a(n_26888), .b(x_in_54_13), .o(n_27116) );
no02f80 g541175 ( .a(n_28578), .b(n_28577), .o(n_28579) );
no02f80 g541176 ( .a(n_28575), .b(n_28574), .o(n_28576) );
no02f80 g541177 ( .a(n_28252), .b(n_28251), .o(n_28253) );
na02f80 g541178 ( .a(n_26887), .b(x_in_14_13), .o(n_27597) );
in01f80 g541179 ( .a(n_27114), .o(n_27115) );
no02f80 g541180 ( .a(n_26887), .b(x_in_14_13), .o(n_27114) );
no02f80 g541181 ( .a(n_28572), .b(n_28571), .o(n_28573) );
na02f80 g541182 ( .a(n_26886), .b(x_in_2_14), .o(n_27596) );
in01f80 g541183 ( .a(n_27112), .o(n_27113) );
no02f80 g541184 ( .a(n_26886), .b(x_in_2_14), .o(n_27112) );
no02f80 g541185 ( .a(n_28453), .b(n_28452), .o(n_28454) );
na02f80 g541186 ( .a(n_26885), .b(x_in_46_13), .o(n_27595) );
in01f80 g541187 ( .a(n_27110), .o(n_27111) );
no02f80 g541188 ( .a(n_26885), .b(x_in_46_13), .o(n_27110) );
no02f80 g541189 ( .a(n_28249), .b(n_28248), .o(n_28250) );
no02f80 g541190 ( .a(n_28450), .b(n_28449), .o(n_28451) );
na02f80 g541191 ( .a(n_26884), .b(x_in_30_13), .o(n_27594) );
in01f80 g541192 ( .a(n_27108), .o(n_27109) );
no02f80 g541193 ( .a(n_26884), .b(x_in_30_13), .o(n_27108) );
no02f80 g541194 ( .a(n_28447), .b(n_28446), .o(n_28448) );
na02f80 g541195 ( .a(n_26883), .b(x_in_62_13), .o(n_27593) );
in01f80 g541196 ( .a(n_27106), .o(n_27107) );
no02f80 g541197 ( .a(n_26883), .b(x_in_62_13), .o(n_27106) );
no02f80 g541198 ( .a(n_28569), .b(n_28568), .o(n_28570) );
no02f80 g541199 ( .a(n_28444), .b(n_28525), .o(n_28445) );
no02f80 g541200 ( .a(n_28349), .b(n_28348), .o(n_28350) );
no02f80 g541201 ( .a(n_28761), .b(n_28760), .o(n_28762) );
na02f80 g541202 ( .a(n_27105), .b(x_in_34_14), .o(n_27760) );
in01f80 g541203 ( .a(n_27280), .o(n_27281) );
no02f80 g541204 ( .a(n_27105), .b(x_in_34_14), .o(n_27280) );
no02f80 g541205 ( .a(n_28566), .b(n_28565), .o(n_28567) );
no02f80 g541206 ( .a(n_28442), .b(n_28441), .o(n_28443) );
na02f80 g541207 ( .a(n_26882), .b(x_in_16_14), .o(n_27592) );
in01f80 g541208 ( .a(n_27103), .o(n_27104) );
no02f80 g541209 ( .a(n_26882), .b(x_in_16_14), .o(n_27103) );
no02f80 g541210 ( .a(n_28563), .b(n_28562), .o(n_28564) );
no02f80 g541211 ( .a(n_28439), .b(n_28438), .o(n_28440) );
na02f80 g541212 ( .a(n_26881), .b(x_in_18_14), .o(n_27591) );
in01f80 g541213 ( .a(n_27101), .o(n_27102) );
no02f80 g541214 ( .a(n_26881), .b(x_in_18_14), .o(n_27101) );
no02f80 g541215 ( .a(n_28560), .b(n_28559), .o(n_28561) );
no02f80 g541216 ( .a(n_28346), .b(n_28345), .o(n_28347) );
no02f80 g541217 ( .a(n_28102), .b(n_28101), .o(n_28103) );
na02f80 g541218 ( .a(n_26880), .b(x_in_32_12), .o(n_27590) );
in01f80 g541219 ( .a(n_27099), .o(n_27100) );
no02f80 g541220 ( .a(n_26880), .b(x_in_32_12), .o(n_27099) );
no02f80 g541221 ( .a(n_28343), .b(n_28342), .o(n_28344) );
na02f80 g541222 ( .a(n_26879), .b(x_in_16_13), .o(n_27589) );
in01f80 g541223 ( .a(n_27097), .o(n_27098) );
no02f80 g541224 ( .a(n_26879), .b(x_in_16_13), .o(n_27097) );
na02f80 g541225 ( .a(n_27279), .b(x_in_48_12), .o(n_27910) );
no02f80 g541226 ( .a(n_28557), .b(n_28556), .o(n_28558) );
in01f80 g541227 ( .a(n_27482), .o(n_27483) );
no02f80 g541228 ( .a(n_27279), .b(x_in_48_12), .o(n_27482) );
na02f80 g541229 ( .a(n_26878), .b(x_in_50_14), .o(n_27588) );
in01f80 g541230 ( .a(n_27095), .o(n_27096) );
no02f80 g541231 ( .a(n_26878), .b(x_in_50_14), .o(n_27095) );
no02f80 g541232 ( .a(n_28244), .b(n_28243), .o(n_28245) );
na02f80 g541233 ( .a(n_27094), .b(x_in_40_12), .o(n_27759) );
in01f80 g541234 ( .a(n_27277), .o(n_27278) );
no02f80 g541235 ( .a(n_27094), .b(x_in_40_12), .o(n_27277) );
no02f80 g541236 ( .a(n_28241), .b(n_28240), .o(n_28242) );
no02f80 g541237 ( .a(n_28554), .b(n_28553), .o(n_28555) );
na02f80 g541238 ( .a(n_26877), .b(x_in_10_14), .o(n_27587) );
in01f80 g541239 ( .a(n_27092), .o(n_27093) );
no02f80 g541240 ( .a(n_26877), .b(x_in_10_14), .o(n_27092) );
no02f80 g541241 ( .a(n_28664), .b(n_28663), .o(n_28665) );
no02f80 g541242 ( .a(n_28551), .b(n_28550), .o(n_28552) );
na02f80 g541243 ( .a(n_26876), .b(x_in_42_14), .o(n_27586) );
in01f80 g541244 ( .a(n_27090), .o(n_27091) );
no02f80 g541245 ( .a(n_26876), .b(x_in_42_14), .o(n_27090) );
no02f80 g541246 ( .a(n_28436), .b(n_28435), .o(n_28437) );
na02f80 g541247 ( .a(n_26582), .b(n_26224), .o(n_26583) );
no02f80 g541248 ( .a(n_28661), .b(n_28660), .o(n_28662) );
na02f80 g541249 ( .a(n_27479), .b(x_in_20_12), .o(n_28020) );
in01f80 g541250 ( .a(n_27663), .o(n_27664) );
no02f80 g541251 ( .a(n_27479), .b(x_in_20_12), .o(n_27663) );
no02f80 g541252 ( .a(n_27969), .b(n_27968), .o(n_27970) );
in01f80 g541253 ( .a(n_28713), .o(n_26875) );
no02f80 g541254 ( .a(n_26581), .b(x_in_52_12), .o(n_28713) );
in01f80 g541255 ( .a(n_27380), .o(n_26874) );
na02f80 g541256 ( .a(n_26581), .b(x_in_52_12), .o(n_27380) );
no02f80 g541257 ( .a(n_28548), .b(n_28547), .o(n_28549) );
na02f80 g541258 ( .a(n_26873), .b(x_in_26_14), .o(n_27585) );
in01f80 g541259 ( .a(n_27088), .o(n_27089) );
no02f80 g541260 ( .a(n_26873), .b(x_in_26_14), .o(n_27088) );
no02f80 g541261 ( .a(n_28237), .b(n_28236), .o(n_28238) );
na02f80 g541262 ( .a(n_27087), .b(x_in_12_13), .o(n_27758) );
in01f80 g541263 ( .a(n_27273), .o(n_27274) );
no02f80 g541264 ( .a(n_27087), .b(x_in_12_13), .o(n_27273) );
in01f80 g541265 ( .a(n_27271), .o(n_27272) );
no02f80 g541266 ( .a(n_27086), .b(x_in_12_14), .o(n_27271) );
na02f80 g541267 ( .a(n_27086), .b(x_in_12_14), .o(n_27757) );
na02f80 g541268 ( .a(n_27086), .b(x_in_12_15), .o(n_27084) );
no02f80 g541269 ( .a(n_28545), .b(n_28544), .o(n_28546) );
na02f80 g541270 ( .a(n_27475), .b(x_in_60_12), .o(n_28018) );
in01f80 g541271 ( .a(n_27658), .o(n_27659) );
no02f80 g541272 ( .a(n_27475), .b(x_in_60_12), .o(n_27658) );
oa22f80 g541273 ( .a(n_26102), .b(n_16497), .c(n_14963), .d(n_14578), .o(n_26872) );
no02f80 g541274 ( .a(n_26619), .b(n_26280), .o(n_26281) );
na03f80 g541275 ( .a(n_26638), .b(n_27270), .c(FE_OFN80_n_27012), .o(n_27750) );
na02f80 g541276 ( .a(n_27269), .b(n_4270), .o(n_27754) );
na03f80 g541277 ( .a(n_26359), .b(n_27474), .c(FE_OFN1114_rst), .o(n_27894) );
na02f80 g541278 ( .a(n_27473), .b(FE_OFN1113_rst), .o(n_27904) );
no02f80 g541279 ( .a(n_26870), .b(n_26869), .o(n_26871) );
in01f80 g541280 ( .a(n_26578), .o(n_26579) );
na02f80 g541281 ( .a(n_26279), .b(x_in_52_13), .o(n_26578) );
na02f80 g541282 ( .a(n_26577), .b(n_280), .o(n_27173) );
na02f80 g541283 ( .a(n_26464), .b(FE_OFN1113_rst), .o(n_27369) );
na02f80 g541284 ( .a(n_26576), .b(FE_OFN1114_rst), .o(n_27164) );
na02f80 g541285 ( .a(n_26462), .b(FE_OFN1109_rst), .o(n_27367) );
no02f80 g541286 ( .a(n_27581), .b(n_27082), .o(n_27083) );
no02f80 g541287 ( .a(n_27581), .b(n_26636), .o(n_27939) );
na02f80 g541288 ( .a(n_26277), .b(n_26276), .o(n_26278) );
na02f80 g541289 ( .a(n_26574), .b(n_26868), .o(n_26575) );
no02f80 g541290 ( .a(n_26886), .b(n_26868), .o(n_27376) );
na02f80 g541291 ( .a(n_26866), .b(n_27078), .o(n_26867) );
no02f80 g541292 ( .a(n_27105), .b(n_27078), .o(n_27937) );
na02f80 g541293 ( .a(n_26864), .b(n_26863), .o(n_26865) );
na02f80 g541294 ( .a(n_26864), .b(n_26361), .o(n_27583) );
na02f80 g541295 ( .a(n_26861), .b(n_26860), .o(n_26862) );
na02f80 g541296 ( .a(n_26861), .b(n_26360), .o(n_28089) );
na02f80 g541297 ( .a(n_26572), .b(n_26859), .o(n_26573) );
no02f80 g541298 ( .a(n_26877), .b(n_26859), .o(n_28036) );
na02f80 g541299 ( .a(n_26570), .b(n_26858), .o(n_26571) );
no02f80 g541300 ( .a(n_26876), .b(n_26858), .o(n_28034) );
na02f80 g541301 ( .a(n_26568), .b(n_26857), .o(n_26569) );
no02f80 g541302 ( .a(n_26873), .b(n_26857), .o(n_28032) );
na02f80 g541303 ( .a(n_26855), .b(n_26854), .o(n_26856) );
na02f80 g541304 ( .a(n_26855), .b(n_26357), .o(n_28030) );
na02f80 g541305 ( .a(n_26852), .b(n_26851), .o(n_26853) );
na02f80 g541306 ( .a(n_26852), .b(n_26354), .o(n_27857) );
no02f80 g541307 ( .a(n_27159), .b(n_26848), .o(n_26567) );
in01f80 g541308 ( .a(n_27402), .o(n_27077) );
na02f80 g541309 ( .a(n_26849), .b(n_26848), .o(n_27402) );
oa12f80 g541310 ( .a(FE_OFN42_n_26563), .b(n_1238), .c(FE_OFN142_n_27449), .o(n_26566) );
oa12f80 g541311 ( .a(FE_OFN42_n_26563), .b(n_1389), .c(FE_OFN142_n_27449), .o(n_26564) );
oa12f80 g541312 ( .a(FE_OFN42_n_26563), .b(n_1736), .c(FE_OFN77_n_27012), .o(n_26562) );
na02f80 g541313 ( .a(n_26845), .b(n_26844), .o(n_26846) );
na02f80 g541314 ( .a(n_26845), .b(n_26353), .o(n_27171) );
no02f80 g541315 ( .a(n_27570), .b(n_27262), .o(n_27075) );
in01f80 g541316 ( .a(n_27792), .o(n_27460) );
na02f80 g541317 ( .a(n_27263), .b(n_27262), .o(n_27792) );
na02f80 g541318 ( .a(n_26560), .b(n_26559), .o(n_26561) );
na02f80 g541319 ( .a(n_26274), .b(n_26273), .o(n_26275) );
oa12f80 g541320 ( .a(n_27071), .b(n_1099), .c(FE_OFN78_n_27012), .o(n_27074) );
oa12f80 g541321 ( .a(n_27071), .b(n_1608), .c(FE_OFN78_n_27012), .o(n_27072) );
na02f80 g541322 ( .a(n_26271), .b(n_26270), .o(n_26272) );
na02f80 g541323 ( .a(n_26279), .b(n_26926), .o(n_26269) );
na02f80 g541324 ( .a(n_26267), .b(n_26266), .o(n_26268) );
no02f80 g541325 ( .a(n_26557), .b(n_26556), .o(n_26558) );
no02f80 g541326 ( .a(n_26557), .b(n_26067), .o(n_27619) );
in01f80 g541327 ( .a(n_28907), .o(n_28757) );
oa12f80 g541328 ( .a(n_26807), .b(n_28385), .c(n_26430), .o(n_28907) );
in01f80 g541329 ( .a(n_29017), .o(n_28840) );
oa12f80 g541330 ( .a(n_26804), .b(n_26428), .c(n_28510), .o(n_29017) );
ao12f80 g541331 ( .a(n_28738), .b(n_27250), .c(n_28737), .o(n_29089) );
in01f80 g541332 ( .a(n_29012), .o(n_28839) );
oa12f80 g541333 ( .a(n_27026), .b(n_26668), .c(n_28509), .o(n_29012) );
in01f80 g541334 ( .a(n_29009), .o(n_28838) );
oa12f80 g541335 ( .a(n_27025), .b(n_26666), .c(n_28508), .o(n_29009) );
in01f80 g541336 ( .a(n_29006), .o(n_28837) );
oa12f80 g541337 ( .a(n_27024), .b(n_26664), .c(n_28507), .o(n_29006) );
in01f80 g541338 ( .a(n_28904), .o(n_28756) );
oa12f80 g541339 ( .a(n_26801), .b(n_28384), .c(n_26421), .o(n_28904) );
in01f80 g541340 ( .a(n_28816), .o(n_28659) );
oa12f80 g541341 ( .a(n_27023), .b(n_26662), .c(n_28281), .o(n_28816) );
in01f80 g541342 ( .a(n_28901), .o(n_28755) );
oa12f80 g541343 ( .a(n_26798), .b(n_28383), .c(n_26418), .o(n_28901) );
in01f80 g541344 ( .a(n_28898), .o(n_28754) );
oa12f80 g541345 ( .a(n_26797), .b(n_28382), .c(n_26416), .o(n_28898) );
in01f80 g541346 ( .a(n_28895), .o(n_28753) );
oa12f80 g541347 ( .a(n_27022), .b(n_28381), .c(n_26660), .o(n_28895) );
in01f80 g541348 ( .a(n_28733), .o(n_28543) );
oa12f80 g541349 ( .a(n_27021), .b(n_26658), .c(n_28142), .o(n_28733) );
oa12f80 g541350 ( .a(n_25499), .b(n_24844), .c(n_28648), .o(n_28864) );
in01f80 g541351 ( .a(n_28658), .o(n_28961) );
oa12f80 g541352 ( .a(n_25777), .b(n_25128), .c(n_28538), .o(n_28658) );
in01f80 g541353 ( .a(n_28892), .o(n_28751) );
oa12f80 g541354 ( .a(n_27020), .b(n_26655), .c(n_28379), .o(n_28892) );
in01f80 g541355 ( .a(n_28889), .o(n_28750) );
oa12f80 g541356 ( .a(n_26795), .b(n_26410), .c(n_28378), .o(n_28889) );
in01f80 g541357 ( .a(n_29003), .o(n_28836) );
oa12f80 g541358 ( .a(n_27019), .b(n_26653), .c(n_28506), .o(n_29003) );
in01f80 g541359 ( .a(n_29000), .o(n_28835) );
oa12f80 g541360 ( .a(n_27018), .b(n_26651), .c(n_28505), .o(n_29000) );
in01f80 g541361 ( .a(n_28730), .o(n_28542) );
oa12f80 g541362 ( .a(n_26792), .b(n_26406), .c(n_28141), .o(n_28730) );
in01f80 g541363 ( .a(n_28997), .o(n_28834) );
oa12f80 g541364 ( .a(n_26793), .b(n_26404), .c(n_28504), .o(n_28997) );
in01f80 g541365 ( .a(n_28886), .o(n_28749) );
oa12f80 g541366 ( .a(n_26791), .b(n_26402), .c(n_28376), .o(n_28886) );
oa12f80 g541367 ( .a(n_26235), .b(n_28140), .c(n_25890), .o(n_28806) );
in01f80 g541368 ( .a(n_28883), .o(n_28747) );
oa12f80 g541369 ( .a(n_26789), .b(n_26400), .c(n_28377), .o(n_28883) );
in01f80 g541370 ( .a(n_28880), .o(n_28746) );
oa12f80 g541371 ( .a(n_26788), .b(n_26398), .c(n_28375), .o(n_28880) );
in01f80 g541372 ( .a(n_28994), .o(n_28833) );
oa12f80 g541373 ( .a(n_26787), .b(n_26395), .c(n_28503), .o(n_28994) );
oa12f80 g541374 ( .a(n_3341), .b(n_28536), .c(n_2227), .o(n_28802) );
na03f80 g541375 ( .a(n_27241), .b(n_28745), .c(n_28650), .o(n_28943) );
in01f80 g541376 ( .a(n_28810), .o(n_28657) );
oa12f80 g541377 ( .a(n_26786), .b(n_26393), .c(n_28278), .o(n_28810) );
in01f80 g541378 ( .a(n_29168), .o(n_29036) );
oa12f80 g541379 ( .a(n_27017), .b(n_26649), .c(n_28710), .o(n_29168) );
in01f80 g541380 ( .a(n_28991), .o(n_28832) );
oa12f80 g541381 ( .a(n_26784), .b(n_26390), .c(n_28502), .o(n_28991) );
in01f80 g541382 ( .a(n_28877), .o(n_28744) );
oa12f80 g541383 ( .a(n_26781), .b(n_26388), .c(n_28373), .o(n_28877) );
in01f80 g541384 ( .a(n_28988), .o(n_28831) );
oa12f80 g541385 ( .a(n_26780), .b(n_26386), .c(n_28501), .o(n_28988) );
in01f80 g541386 ( .a(n_28874), .o(n_28743) );
oa12f80 g541387 ( .a(n_26779), .b(n_26384), .c(n_28372), .o(n_28874) );
in01f80 g541388 ( .a(n_28985), .o(n_28829) );
oa12f80 g541389 ( .a(n_26778), .b(n_26382), .c(n_28500), .o(n_28985) );
in01f80 g541390 ( .a(n_28637), .o(n_28433) );
oa12f80 g541391 ( .a(n_26777), .b(n_26379), .c(n_28017), .o(n_28637) );
in01f80 g541392 ( .a(n_28656), .o(n_28956) );
oa12f80 g541393 ( .a(n_27016), .b(n_28277), .c(n_26647), .o(n_28656) );
in01f80 g541394 ( .a(n_28807), .o(n_28655) );
oa12f80 g541395 ( .a(n_27015), .b(n_26645), .c(n_28276), .o(n_28807) );
in01f80 g541396 ( .a(n_28982), .o(n_28828) );
oa12f80 g541397 ( .a(n_26776), .b(n_26376), .c(n_28499), .o(n_28982) );
in01f80 g541398 ( .a(n_28725), .o(n_28541) );
oa12f80 g541399 ( .a(n_27247), .b(n_26972), .c(n_28139), .o(n_28725) );
ao12f80 g541400 ( .a(n_28431), .b(n_26520), .c(n_28430), .o(n_28805) );
oa12f80 g541401 ( .a(n_25584), .b(n_28340), .c(n_24974), .o(n_28717) );
in01f80 g541402 ( .a(n_28742), .o(n_29079) );
oa12f80 g541403 ( .a(n_26551), .b(n_28646), .c(n_26196), .o(n_28742) );
ao12f80 g541404 ( .a(n_13618), .b(n_26549), .c(n_14649), .o(n_27397) );
in01f80 g541405 ( .a(n_28978), .o(n_28826) );
oa12f80 g541406 ( .a(n_26775), .b(n_28498), .c(n_26374), .o(n_28978) );
oa12f80 g541407 ( .a(n_25764), .b(n_25110), .c(n_28534), .o(n_28799) );
in01f80 g541408 ( .a(n_28973), .o(n_28825) );
oa12f80 g541409 ( .a(n_26772), .b(n_28497), .c(n_26372), .o(n_28973) );
oa12f80 g541410 ( .a(n_10768), .b(FE_OFN636_n_26260), .c(n_8994), .o(n_26261) );
in01f80 g541411 ( .a(n_29076), .o(n_29077) );
oa12f80 g541412 ( .a(n_27439), .b(n_27199), .c(n_28370), .o(n_29076) );
in01f80 g541413 ( .a(n_27651), .o(n_27652) );
oa12f80 g541414 ( .a(n_27457), .b(n_27456), .c(x_in_36_13), .o(n_27651) );
in01f80 g541415 ( .a(n_29093), .o(n_28912) );
oa12f80 g541416 ( .a(n_27644), .b(n_27392), .c(n_28631), .o(n_29093) );
in01f80 g541417 ( .a(n_28518), .o(n_28714) );
oa12f80 g541418 ( .a(n_26518), .b(n_27900), .c(n_26107), .o(n_28518) );
in01f80 g541419 ( .a(n_28970), .o(n_28824) );
oa12f80 g541420 ( .a(n_26768), .b(n_28496), .c(n_26370), .o(n_28970) );
in01f80 g541421 ( .a(n_28720), .o(n_28540) );
oa12f80 g541422 ( .a(n_27013), .b(n_26641), .c(n_28138), .o(n_28720) );
oa12f80 g541423 ( .a(n_27440), .b(n_28632), .c(n_27201), .o(n_29129) );
in01f80 g541424 ( .a(n_28654), .o(n_28951) );
ao12f80 g541425 ( .a(n_26471), .b(n_28532), .c(n_26832), .o(n_28654) );
in01f80 g541426 ( .a(n_28653), .o(n_28949) );
oa12f80 g541427 ( .a(n_25761), .b(n_25106), .c(n_28530), .o(n_28653) );
in01f80 g541428 ( .a(n_28967), .o(n_28823) );
oa12f80 g541429 ( .a(n_27244), .b(n_26964), .c(n_28495), .o(n_28967) );
oa12f80 g541430 ( .a(n_27434), .b(n_27432), .c(n_25987), .o(n_27650) );
oa12f80 g541431 ( .a(n_27450), .b(n_372), .c(n_27452), .o(n_27453) );
oa12f80 g541432 ( .a(n_27450), .b(n_216), .c(FE_OFN134_n_27449), .o(n_27451) );
oa12f80 g541433 ( .a(n_27450), .b(n_217), .c(FE_OFN134_n_27449), .o(n_27448) );
oa12f80 g541434 ( .a(n_27240), .b(n_27236), .c(n_25752), .o(n_27447) );
oa12f80 g541435 ( .a(n_27051), .b(n_944), .c(FE_OFN1117_rst), .o(n_27054) );
oa12f80 g541436 ( .a(n_27051), .b(n_1343), .c(FE_OFN1117_rst), .o(n_27052) );
oa12f80 g541437 ( .a(n_27051), .b(n_775), .c(FE_OFN102_n_27449), .o(n_27050) );
oa12f80 g541438 ( .a(n_27044), .b(n_937), .c(FE_OFN1121_rst), .o(n_27048) );
oa12f80 g541439 ( .a(n_27044), .b(n_317), .c(FE_OFN1121_rst), .o(n_27045) );
oa12f80 g541440 ( .a(n_26256), .b(n_124), .c(FE_OFN1117_rst), .o(n_26258) );
oa12f80 g541441 ( .a(n_26256), .b(n_968), .c(FE_OFN102_n_27449), .o(n_26257) );
oa12f80 g541442 ( .a(n_26256), .b(n_745), .c(FE_OFN102_n_27449), .o(n_26255) );
in01f80 g541443 ( .a(n_27648), .o(n_27649) );
oa12f80 g541444 ( .a(n_27445), .b(n_27456), .c(x_in_36_12), .o(n_27648) );
oa12f80 g541445 ( .a(n_28650), .b(n_26960), .c(n_28374), .o(n_28861) );
ao12f80 g541446 ( .a(n_26743), .b(n_26544), .c(n_26543), .o(n_27195) );
ao12f80 g541447 ( .a(n_26302), .b(n_26253), .c(n_26252), .o(n_26959) );
ao12f80 g541448 ( .a(n_26300), .b(n_26251), .c(n_26250), .o(n_26957) );
ao12f80 g541449 ( .a(n_26298), .b(n_26249), .c(n_26248), .o(n_26952) );
ao12f80 g541450 ( .a(n_26296), .b(n_26247), .c(n_26246), .o(n_26950) );
ao12f80 g541451 ( .a(n_26294), .b(n_26245), .c(n_26244), .o(n_26948) );
ao12f80 g541452 ( .a(n_26508), .b(n_5605), .c(n_3641), .o(n_27395) );
in01f80 g541453 ( .a(n_27174), .o(n_26817) );
ao12f80 g541454 ( .a(n_25973), .b(FE_OFN636_n_26260), .c(n_25972), .o(n_27174) );
oa12f80 g541455 ( .a(n_27249), .b(n_28738), .c(n_28737), .o(n_28739) );
ao22s80 g541456 ( .a(n_25779), .b(n_28648), .c(n_25778), .d(n_28380), .o(n_28649) );
ao22s80 g541457 ( .a(n_26005), .b(n_28538), .c(n_26004), .d(n_28280), .o(n_28539) );
ao22s80 g541458 ( .a(n_28536), .b(n_3711), .c(n_28279), .d(n_3710), .o(n_28537) );
oa12f80 g541459 ( .a(n_26529), .b(n_26764), .c(x_in_18_15), .o(n_29198) );
ao22s80 g541460 ( .a(n_28646), .b(n_26835), .c(n_28371), .d(n_26834), .o(n_28647) );
oa12f80 g541461 ( .a(n_26519), .b(n_28431), .c(n_28430), .o(n_28432) );
ao22s80 g541462 ( .a(n_28340), .b(n_25859), .c(n_28016), .d(n_25858), .o(n_28341) );
ao12f80 g541463 ( .a(n_27009), .b(n_27008), .c(n_27007), .o(n_27254) );
in01f80 g541464 ( .a(n_27374), .o(n_27035) );
oa12f80 g541465 ( .a(n_26227), .b(n_26549), .c(n_26226), .o(n_27374) );
ao22s80 g541466 ( .a(n_25998), .b(n_28534), .c(n_25997), .d(n_28275), .o(n_28535) );
ao22s80 g541467 ( .a(n_27456), .b(x_in_36_15), .c(n_27444), .d(n_27230), .o(n_29675) );
ao22s80 g541468 ( .a(n_28532), .b(n_27064), .c(n_28274), .d(n_27063), .o(n_28533) );
ao22s80 g541469 ( .a(n_25993), .b(n_28530), .c(n_25992), .d(n_28273), .o(n_28531) );
oa22f80 g541470 ( .a(FE_OFN791_n_28272), .b(n_29033), .c(n_268), .d(FE_OFN96_n_27449), .o(n_28529) );
oa22f80 g541471 ( .a(n_28137), .b(FE_OFN303_n_3069), .c(n_1119), .d(FE_OFN114_n_27449), .o(n_28429) );
oa22f80 g541472 ( .a(n_28135), .b(FE_OFN306_n_3069), .c(n_1956), .d(FE_OFN93_n_27449), .o(n_28427) );
oa22f80 g541473 ( .a(FE_OFN666_n_26759), .b(n_28608), .c(n_1061), .d(FE_OFN96_n_27449), .o(n_26816) );
oa22f80 g541474 ( .a(n_28270), .b(FE_OFN249_n_4162), .c(n_1246), .d(FE_OFN124_n_27449), .o(n_28528) );
oa22f80 g541475 ( .a(FE_OFN662_n_27899), .b(n_28608), .c(n_767), .d(FE_OFN96_n_27449), .o(n_28235) );
oa22f80 g541476 ( .a(n_26328), .b(FE_OFN306_n_3069), .c(n_1885), .d(FE_OFN355_n_4860), .o(n_27029) );
oa22f80 g541477 ( .a(n_28133), .b(FE_OFN296_n_3069), .c(n_941), .d(FE_OFN358_n_4860), .o(n_28425) );
oa22f80 g541478 ( .a(n_28131), .b(FE_OFN312_n_3069), .c(n_1002), .d(FE_OFN113_n_27449), .o(n_28424) );
oa22f80 g541479 ( .a(n_28129), .b(FE_OFN296_n_3069), .c(n_947), .d(FE_OFN80_n_27012), .o(n_28422) );
oa22f80 g541480 ( .a(n_27444), .b(n_29194), .c(n_27456), .d(x_in_36_14), .o(n_29576) );
na02f80 g541506 ( .a(n_26764), .b(x_in_18_15), .o(n_26529) );
na02f80 g541507 ( .a(n_26807), .b(n_26431), .o(n_28474) );
na02f80 g541508 ( .a(n_27250), .b(n_26977), .o(n_28590) );
na02f80 g541509 ( .a(n_26804), .b(n_26429), .o(n_28593) );
no02f80 g541510 ( .a(FE_OFN636_n_26260), .b(n_25972), .o(n_25973) );
na02f80 g541511 ( .a(n_27026), .b(n_26669), .o(n_28587) );
na02f80 g541512 ( .a(n_27025), .b(n_26667), .o(n_28584) );
na02f80 g541513 ( .a(n_27024), .b(n_26665), .o(n_28581) );
na02f80 g541514 ( .a(n_26801), .b(n_26422), .o(n_28471) );
na02f80 g541515 ( .a(n_27023), .b(n_26663), .o(n_28352) );
no02f80 g541516 ( .a(n_26978), .b(x_in_60_13), .o(n_27249) );
na02f80 g541517 ( .a(n_26798), .b(n_26419), .o(n_28468) );
na02f80 g541518 ( .a(n_26797), .b(n_26417), .o(n_28465) );
na02f80 g541519 ( .a(n_27022), .b(n_26661), .o(n_28462) );
na02f80 g541520 ( .a(n_27021), .b(n_26659), .o(n_28256) );
na02f80 g541521 ( .a(n_27020), .b(n_26656), .o(n_28459) );
na02f80 g541522 ( .a(n_26795), .b(n_26411), .o(n_28456) );
na02f80 g541523 ( .a(n_27019), .b(n_26654), .o(n_28578) );
na02f80 g541524 ( .a(n_27018), .b(n_26652), .o(n_28575) );
na02f80 g541525 ( .a(n_26793), .b(n_26405), .o(n_28572) );
na02f80 g541526 ( .a(n_26792), .b(n_26407), .o(n_28252) );
na02f80 g541527 ( .a(n_26791), .b(n_26403), .o(n_28453) );
na02f80 g541528 ( .a(n_26235), .b(n_25891), .o(n_28249) );
na02f80 g541529 ( .a(n_26789), .b(n_26401), .o(n_28450) );
na02f80 g541530 ( .a(n_26788), .b(n_26399), .o(n_28447) );
na02f80 g541531 ( .a(n_26787), .b(n_26396), .o(n_28569) );
na02f80 g541532 ( .a(n_25729), .b(n_25728), .o(n_25730) );
na02f80 g541533 ( .a(n_26786), .b(n_26394), .o(n_28349) );
na02f80 g541534 ( .a(n_27017), .b(n_26650), .o(n_28761) );
na02f80 g541535 ( .a(n_26784), .b(n_26391), .o(n_28566) );
na02f80 g541536 ( .a(n_26781), .b(n_26389), .o(n_28442) );
na02f80 g541537 ( .a(n_26780), .b(n_26387), .o(n_28563) );
na02f80 g541538 ( .a(n_26779), .b(n_26385), .o(n_28439) );
na02f80 g541539 ( .a(n_26778), .b(n_26383), .o(n_28560) );
na02f80 g541540 ( .a(n_26648), .b(n_27016), .o(n_28346) );
na02f80 g541541 ( .a(n_26777), .b(n_26380), .o(n_28102) );
na02f80 g541542 ( .a(n_27015), .b(n_26646), .o(n_28343) );
na02f80 g541543 ( .a(n_26776), .b(n_26377), .o(n_28557) );
in01f80 g541544 ( .a(n_27645), .o(n_27646) );
na02f80 g541545 ( .a(n_27443), .b(n_27204), .o(n_27645) );
na02f80 g541546 ( .a(n_27247), .b(n_26973), .o(n_28244) );
na02f80 g541547 ( .a(n_26520), .b(n_26117), .o(n_28241) );
no02f80 g541548 ( .a(n_26118), .b(x_in_32_13), .o(n_26519) );
na02f80 g541549 ( .a(n_26549), .b(n_26226), .o(n_26227) );
na02f80 g541550 ( .a(n_26775), .b(n_26375), .o(n_28554) );
in01f80 g541551 ( .a(n_27441), .o(n_27442) );
na02f80 g541552 ( .a(n_27246), .b(n_26970), .o(n_27441) );
no02f80 g541553 ( .a(n_26971), .b(x_in_48_13), .o(n_27245) );
na02f80 g541554 ( .a(n_27202), .b(n_27440), .o(n_28664) );
na02f80 g541555 ( .a(n_26772), .b(n_26373), .o(n_28551) );
na02f80 g541556 ( .a(n_27439), .b(n_27200), .o(n_28436) );
no02f80 g541557 ( .a(n_26224), .b(FE_OFN368_n_26312), .o(n_26225) );
na02f80 g541558 ( .a(n_27644), .b(n_27393), .o(n_28661) );
no02f80 g541559 ( .a(n_26221), .b(FE_OFN23_n_26609), .o(n_26222) );
na02f80 g541560 ( .a(n_26518), .b(n_26108), .o(n_27969) );
na02f80 g541561 ( .a(n_26768), .b(n_26371), .o(n_28548) );
na02f80 g541562 ( .a(n_27013), .b(n_26642), .o(n_28237) );
in01f80 g541563 ( .a(n_27830), .o(n_27831) );
na02f80 g541564 ( .a(n_27388), .b(n_27643), .o(n_27830) );
na02f80 g541565 ( .a(n_27244), .b(n_26965), .o(n_28545) );
na03f80 g541566 ( .a(n_25226), .b(n_26368), .c(FE_OFN80_n_27012), .o(n_27450) );
na02f80 g541567 ( .a(n_27456), .b(x_in_36_13), .o(n_27457) );
na03f80 g541568 ( .a(n_24860), .b(FE_OFN901_n_26098), .c(FE_OFN421_n_16909), .o(n_27044) );
na02f80 g541569 ( .a(n_26099), .b(FE_OFN290_n_27194), .o(n_27071) );
na02f80 g541570 ( .a(n_26961), .b(n_28650), .o(n_28444) );
na02f80 g541571 ( .a(n_27456), .b(x_in_36_12), .o(n_27445) );
na02f80 g541572 ( .a(n_25626), .b(n_4270), .o(n_26256) );
no02f80 g541573 ( .a(n_25866), .b(n_26609), .o(n_26517) );
na02f80 g541574 ( .a(n_26764), .b(n_4270), .o(n_27051) );
in01f80 g541575 ( .a(n_27474), .o(n_27473) );
ao22s80 g541576 ( .a(n_26020), .b(n_9719), .c(n_25821), .d(n_12353), .o(n_27474) );
na02f80 g541577 ( .a(n_26762), .b(FE_OFN330_n_4860), .o(n_27205) );
no02f80 g541578 ( .a(n_26559), .b(FE_OFN23_n_26609), .o(n_26761) );
ao12f80 g541579 ( .a(n_10323), .b(n_25267), .c(n_9372), .o(n_26743) );
ao12f80 g541580 ( .a(n_10324), .b(n_24963), .c(n_9369), .o(n_26302) );
ao12f80 g541581 ( .a(n_10322), .b(n_24961), .c(n_9384), .o(n_26300) );
ao12f80 g541582 ( .a(n_10321), .b(n_24959), .c(n_9381), .o(n_26298) );
ao12f80 g541583 ( .a(n_10320), .b(n_24955), .c(n_9378), .o(n_26296) );
ao12f80 g541584 ( .a(n_10319), .b(n_24953), .c(n_9375), .o(n_26294) );
oa12f80 g541585 ( .a(n_11338), .b(n_26217), .c(n_12825), .o(n_26218) );
oa12f80 g541586 ( .a(n_26515), .b(n_26217), .c(n_25910), .o(n_26909) );
in01f80 g541587 ( .a(n_28339), .o(n_28628) );
oa12f80 g541588 ( .a(n_2158), .b(n_28234), .c(n_3267), .o(n_28339) );
in01f80 g541589 ( .a(n_26605), .o(n_27161) );
oa12f80 g541590 ( .a(n_3485), .b(n_25264), .c(n_9709), .o(n_26605) );
no02f80 g541591 ( .a(n_27008), .b(n_27007), .o(n_27009) );
in01f80 g541592 ( .a(n_27006), .o(n_27373) );
na02f80 g541593 ( .a(n_26759), .b(n_27007), .o(n_27006) );
na02f80 g541594 ( .a(n_28525), .b(n_26963), .o(n_28745) );
oa12f80 g541595 ( .a(n_27340), .b(n_28641), .c(n_26841), .o(n_28766) );
oa12f80 g541596 ( .a(n_15834), .b(n_26216), .c(n_16493), .o(n_26586) );
na03f80 g541597 ( .a(n_25728), .b(n_25729), .c(n_12421), .o(n_26215) );
oa12f80 g541598 ( .a(n_27241), .b(n_32744), .c(x_in_36_13), .o(n_28860) );
in01f80 g541599 ( .a(n_28338), .o(n_28623) );
oa12f80 g541600 ( .a(n_26613), .b(n_26001), .c(n_28228), .o(n_28338) );
in01f80 g541601 ( .a(n_28643), .o(n_28856) );
oa12f80 g541602 ( .a(n_27499), .b(n_28521), .c(n_27067), .o(n_28643) );
in01f80 g541603 ( .a(n_28524), .o(n_28781) );
ao12f80 g541604 ( .a(n_27130), .b(n_28407), .c(n_27578), .o(n_28524) );
in01f80 g541605 ( .a(n_28523), .o(n_28778) );
oa12f80 g541606 ( .a(n_26612), .b(n_25999), .c(n_28404), .o(n_28523) );
ao22s80 g541607 ( .a(n_26611), .b(n_26637), .c(x_out_49_30), .d(FE_OFN280_n_16656), .o(n_27434) );
ao22s80 g541608 ( .a(n_26314), .b(n_26358), .c(x_out_51_29), .d(FE_OFN274_n_16893), .o(n_27240) );
oa12f80 g541609 ( .a(n_27432), .b(n_556), .c(FE_OFN131_n_27449), .o(n_27433) );
oa12f80 g541610 ( .a(n_27236), .b(n_935), .c(FE_OFN353_n_4860), .o(n_27237) );
oa12f80 g541611 ( .a(n_27639), .b(n_287), .c(FE_OFN20_n_27452), .o(n_27641) );
oa12f80 g541612 ( .a(n_27639), .b(n_109), .c(FE_OFN329_n_4860), .o(n_27640) );
oa12f80 g541613 ( .a(FE_OFN316_n_26999), .b(n_1321), .c(FE_OFN134_n_27449), .o(n_27001) );
oa12f80 g541614 ( .a(FE_OFN316_n_26999), .b(n_432), .c(FE_OFN134_n_27449), .o(n_27000) );
ao12f80 g541615 ( .a(n_9183), .b(n_25937), .c(n_10961), .o(n_25968) );
no03m80 g541616 ( .a(n_10962), .b(n_25689), .c(n_3820), .o(n_26508) );
ao12f80 g541617 ( .a(n_14089), .b(n_25966), .c(n_15025), .o(n_26619) );
ao12f80 g541618 ( .a(FE_OFN542_n_23570), .b(n_26694), .c(n_26693), .o(n_27086) );
oa12f80 g541619 ( .a(n_11469), .b(n_26501), .c(n_11857), .o(n_26870) );
oa12f80 g541620 ( .a(n_25627), .b(n_24871), .c(n_25516), .o(n_26563) );
oa12f80 g541621 ( .a(n_14290), .b(n_25964), .c(n_15106), .o(n_25965) );
ao12f80 g541622 ( .a(n_28205), .b(n_28204), .c(n_28203), .o(n_28421) );
in01f80 g541623 ( .a(n_26855), .o(n_26901) );
ao12f80 g541624 ( .a(n_25687), .b(n_25963), .c(n_25686), .o(n_26855) );
ao12f80 g541625 ( .a(n_26367), .b(n_26366), .c(n_26365), .o(n_26998) );
oa12f80 g541626 ( .a(n_15572), .b(n_25963), .c(n_15837), .o(n_26277) );
ao12f80 g541627 ( .a(n_28202), .b(n_28201), .c(n_28200), .o(n_28420) );
oa12f80 g541628 ( .a(n_26093), .b(n_26092), .c(n_26091), .o(n_27129) );
in01f80 g541629 ( .a(n_27581), .o(n_26997) );
oa12f80 g541630 ( .a(n_26105), .b(n_26104), .c(n_26103), .o(n_27581) );
ao12f80 g541631 ( .a(n_28197), .b(n_28196), .c(n_28195), .o(n_28419) );
oa12f80 g541632 ( .a(n_26364), .b(n_26363), .c(n_26362), .o(n_27301) );
ao22s80 g541633 ( .a(n_27532), .b(n_28641), .c(n_27531), .d(n_28268), .o(n_28642) );
ao12f80 g541634 ( .a(n_28194), .b(n_28193), .c(n_28192), .o(n_28418) );
oa12f80 g541635 ( .a(n_25865), .b(n_25864), .c(n_26090), .o(n_26896) );
ao12f80 g541636 ( .a(n_28191), .b(n_28190), .c(n_28189), .o(n_28417) );
oa12f80 g541637 ( .a(n_25863), .b(n_25862), .c(n_26089), .o(n_26895) );
ao12f80 g541638 ( .a(n_27925), .b(n_27924), .c(n_27923), .o(n_28233) );
ao12f80 g541639 ( .a(n_28078), .b(n_28077), .c(n_28076), .o(n_28337) );
oa12f80 g541640 ( .a(n_26088), .b(n_26087), .c(n_26086), .o(n_27124) );
in01f80 g541641 ( .a(n_26852), .o(n_27123) );
ao12f80 g541642 ( .a(n_25906), .b(n_26216), .c(n_25905), .o(n_26852) );
ao12f80 g541643 ( .a(n_28075), .b(n_28074), .c(n_28073), .o(n_28336) );
oa12f80 g541644 ( .a(n_26085), .b(n_26084), .c(n_26083), .o(n_27122) );
ao12f80 g541645 ( .a(n_28072), .b(n_28071), .c(n_28070), .o(n_28335) );
oa12f80 g541646 ( .a(n_26082), .b(n_26081), .c(n_26080), .o(n_27121) );
ao12f80 g541647 ( .a(n_28069), .b(n_28068), .c(n_28067), .o(n_28334) );
oa12f80 g541648 ( .a(n_25861), .b(n_25860), .c(n_26079), .o(n_26889) );
ao12f80 g541649 ( .a(n_27787), .b(n_27786), .c(n_27785), .o(n_28098) );
oa12f80 g541650 ( .a(n_26356), .b(n_26420), .c(n_26355), .o(n_27286) );
ao12f80 g541651 ( .a(n_28066), .b(n_28065), .c(n_28064), .o(n_28333) );
oa22f80 g541652 ( .a(n_26544), .b(n_25760), .c(n_26408), .d(n_26543), .o(n_27118) );
ao12f80 g541653 ( .a(n_28063), .b(n_28062), .c(n_28061), .o(n_28332) );
oa22f80 g541654 ( .a(n_26253), .b(n_25447), .c(n_26131), .d(n_26252), .o(n_26888) );
ao12f80 g541655 ( .a(n_28188), .b(n_28187), .c(n_28186), .o(n_28416) );
ao12f80 g541656 ( .a(n_28180), .b(n_28179), .c(n_28178), .o(n_28415) );
ao12f80 g541657 ( .a(n_28185), .b(n_28184), .c(n_28183), .o(n_28414) );
ao12f80 g541658 ( .a(n_27782), .b(n_27781), .c(n_27780), .o(n_28097) );
oa22f80 g541659 ( .a(n_26251), .b(n_25446), .c(n_26130), .d(n_26250), .o(n_26887) );
in01f80 g541660 ( .a(n_26574), .o(n_26886) );
ao12f80 g541661 ( .a(n_25630), .b(n_25629), .c(n_25628), .o(n_26574) );
ao12f80 g541662 ( .a(n_27779), .b(n_27778), .c(n_27777), .o(n_28096) );
ao12f80 g541663 ( .a(n_28059), .b(n_28058), .c(n_28057), .o(n_28331) );
oa22f80 g541664 ( .a(n_26249), .b(n_25449), .c(n_26129), .d(n_26248), .o(n_26885) );
ao12f80 g541665 ( .a(n_28056), .b(n_28055), .c(n_28054), .o(n_28330) );
in01f80 g541666 ( .a(n_26279), .o(n_26577) );
oa12f80 g541667 ( .a(n_25358), .b(n_25357), .c(n_25356), .o(n_26279) );
oa22f80 g541668 ( .a(n_26247), .b(n_25445), .c(n_26126), .d(n_26246), .o(n_26884) );
ao12f80 g541669 ( .a(n_28053), .b(n_28052), .c(n_28051), .o(n_28329) );
oa22f80 g541670 ( .a(n_26245), .b(n_25444), .c(n_26124), .d(n_26244), .o(n_26883) );
ao12f80 g541671 ( .a(n_28176), .b(n_28175), .c(n_28174), .o(n_28413) );
ao12f80 g541672 ( .a(n_28025), .b(n_28234), .c(n_28024), .o(n_28328) );
ao12f80 g541673 ( .a(n_28050), .b(n_28049), .c(n_28048), .o(n_28327) );
oa22f80 g541674 ( .a(n_32744), .b(x_in_36_15), .c(n_27231), .d(n_27230), .o(n_29385) );
ao12f80 g541675 ( .a(n_27922), .b(n_27921), .c(n_27920), .o(n_28232) );
ao12f80 g541676 ( .a(n_28388), .b(n_28387), .c(n_28386), .o(n_28640) );
ao12f80 g541677 ( .a(n_28172), .b(n_28171), .c(n_28170), .o(n_28412) );
in01f80 g541678 ( .a(n_26866), .o(n_27105) );
ao12f80 g541679 ( .a(n_25872), .b(n_25871), .c(n_25870), .o(n_26866) );
in01f80 g541680 ( .a(n_26557), .o(n_26467) );
oa12f80 g541681 ( .a(n_25632), .b(n_25966), .c(n_25631), .o(n_26557) );
ao12f80 g541682 ( .a(n_28045), .b(n_28044), .c(n_28043), .o(n_28326) );
in01f80 g541683 ( .a(n_26845), .o(n_26882) );
ao12f80 g541684 ( .a(n_25661), .b(n_25660), .c(n_25659), .o(n_26845) );
ao12f80 g541685 ( .a(n_28167), .b(n_28166), .c(n_28165), .o(n_28411) );
ao12f80 g541686 ( .a(n_28042), .b(n_28041), .c(n_28040), .o(n_28325) );
in01f80 g541687 ( .a(n_26864), .o(n_26881) );
ao12f80 g541688 ( .a(n_25635), .b(n_25634), .c(n_25633), .o(n_26864) );
ao12f80 g541689 ( .a(n_28164), .b(n_28163), .c(n_28162), .o(n_28410) );
ao12f80 g541690 ( .a(n_27919), .b(n_27918), .c(n_27917), .o(n_28231) );
ao12f80 g541691 ( .a(n_27607), .b(n_27606), .c(n_27605), .o(n_27945) );
oa12f80 g541692 ( .a(n_25857), .b(n_26078), .c(n_25856), .o(n_26880) );
ao12f80 g541693 ( .a(n_27916), .b(n_27915), .c(n_27914), .o(n_28230) );
oa12f80 g541694 ( .a(n_25855), .b(n_25854), .c(n_26077), .o(n_26879) );
ao22s80 g541695 ( .a(n_26939), .b(n_28228), .c(n_26938), .d(n_27740), .o(n_28229) );
ao12f80 g541696 ( .a(n_28161), .b(n_28160), .c(n_28159), .o(n_28409) );
oa12f80 g541697 ( .a(n_26352), .b(n_26351), .c(n_26632), .o(n_27279) );
in01f80 g541698 ( .a(n_26861), .o(n_26878) );
ao12f80 g541699 ( .a(n_25606), .b(n_25605), .c(n_25604), .o(n_26861) );
in01f80 g541700 ( .a(n_27570), .o(n_27263) );
oa12f80 g541701 ( .a(n_26101), .b(n_26501), .c(n_26100), .o(n_27570) );
ao22s80 g541702 ( .a(n_27680), .b(n_28521), .c(n_27679), .d(n_28125), .o(n_28522) );
ao12f80 g541703 ( .a(n_27775), .b(n_27774), .c(n_27773), .o(n_28095) );
oa12f80 g541704 ( .a(n_26076), .b(n_26075), .c(n_26350), .o(n_27094) );
ao12f80 g541705 ( .a(n_27772), .b(n_27771), .c(n_27770), .o(n_28094) );
in01f80 g541706 ( .a(n_27159), .o(n_26849) );
oa12f80 g541707 ( .a(n_25613), .b(n_25964), .c(n_25612), .o(n_27159) );
ao22s80 g541708 ( .a(n_27742), .b(n_28407), .c(n_27741), .d(n_28008), .o(n_28408) );
ao12f80 g541709 ( .a(n_28156), .b(n_28155), .c(n_28154), .o(n_28406) );
ao12f80 g541710 ( .a(n_26074), .b(n_26073), .c(n_26072), .o(n_26702) );
in01f80 g541711 ( .a(n_26560), .o(n_26464) );
ao12f80 g541712 ( .a(n_25655), .b(n_25688), .c(n_25654), .o(n_26560) );
in01f80 g541713 ( .a(n_26572), .o(n_26877) );
ao12f80 g541714 ( .a(n_25622), .b(n_25938), .c(n_25621), .o(n_26572) );
oa12f80 g541715 ( .a(n_15508), .b(n_25938), .c(n_15847), .o(n_26274) );
ao22s80 g541716 ( .a(n_26937), .b(n_28404), .c(n_26936), .d(n_28007), .o(n_28405) );
ao12f80 g541717 ( .a(n_28287), .b(n_28286), .c(n_28285), .o(n_28517) );
ao12f80 g541718 ( .a(n_25869), .b(n_25868), .c(n_25867), .o(n_26463) );
in01f80 g541719 ( .a(n_26191), .o(n_26576) );
ao22s80 g541720 ( .a(n_25937), .b(n_11601), .c(n_24939), .d(n_11600), .o(n_26191) );
ao12f80 g541721 ( .a(n_28028), .b(n_28027), .c(n_28026), .o(n_28323) );
ao12f80 g541722 ( .a(n_28153), .b(n_28152), .c(n_28151), .o(n_28403) );
in01f80 g541723 ( .a(n_26570), .o(n_26876) );
ao12f80 g541724 ( .a(n_25620), .b(n_25936), .c(n_25619), .o(n_26570) );
oa12f80 g541725 ( .a(n_15499), .b(n_25936), .c(n_15775), .o(n_26271) );
ao12f80 g541726 ( .a(n_26114), .b(n_26443), .c(n_26113), .o(n_26698) );
in01f80 g541727 ( .a(n_26582), .o(n_26462) );
ao12f80 g541728 ( .a(n_25603), .b(n_25602), .c(n_25601), .o(n_26582) );
ao12f80 g541729 ( .a(n_28284), .b(n_28283), .c(n_28282), .o(n_28516) );
oa12f80 g541730 ( .a(n_26630), .b(n_26629), .c(n_27211), .o(n_27479) );
ao12f80 g541731 ( .a(n_26111), .b(n_26459), .c(n_26110), .o(n_26697) );
ao12f80 g541732 ( .a(n_28150), .b(n_28149), .c(n_28148), .o(n_28402) );
ao12f80 g541733 ( .a(n_27391), .b(n_27390), .c(n_27389), .o(n_27798) );
oa12f80 g541734 ( .a(n_25570), .b(n_25847), .c(n_25569), .o(n_26581) );
in01f80 g541735 ( .a(n_26568), .o(n_26873) );
ao12f80 g541736 ( .a(n_25608), .b(n_25935), .c(n_25607), .o(n_26568) );
ao12f80 g541737 ( .a(n_26070), .b(n_26069), .c(n_26068), .o(n_26695) );
oa12f80 g541738 ( .a(n_15486), .b(n_25935), .c(n_15762), .o(n_26267) );
ao12f80 g541739 ( .a(n_27769), .b(n_27768), .c(n_27767), .o(n_28091) );
oa22f80 g541740 ( .a(n_26694), .b(n_25759), .c(n_26381), .d(n_26693), .o(n_27087) );
oa12f80 g541741 ( .a(n_27196), .b(n_27197), .c(x_in_44_15), .o(n_29422) );
ao12f80 g541742 ( .a(n_28147), .b(n_28146), .c(n_28145), .o(n_28399) );
ao12f80 g541743 ( .a(n_28082), .b(n_28081), .c(n_28080), .o(n_28322) );
oa12f80 g541744 ( .a(n_26628), .b(n_26670), .c(n_26627), .o(n_27475) );
oa22f80 g541745 ( .a(n_26459), .b(FE_OFN247_n_4162), .c(n_219), .d(FE_OFN1181_rst), .o(n_26460) );
oa22f80 g541746 ( .a(FE_OFN1055_n_25805), .b(FE_OFN312_n_3069), .c(n_205), .d(n_29264), .o(n_26688) );
oa22f80 g541747 ( .a(FE_OFN1039_n_27890), .b(FE_OFN312_n_3069), .c(n_730), .d(n_29264), .o(n_28321) );
oa22f80 g541748 ( .a(FE_OFN438_n_27889), .b(n_28608), .c(n_1015), .d(n_29264), .o(n_28320) );
oa22f80 g541749 ( .a(FE_OFN730_n_27888), .b(n_27933), .c(n_276), .d(FE_OFN1108_rst), .o(n_28319) );
oa22f80 g541750 ( .a(FE_OFN746_n_26604), .b(n_28608), .c(n_680), .d(FE_OFN336_n_4860), .o(n_27399) );
oa22f80 g541751 ( .a(n_28123), .b(FE_OFN259_n_4280), .c(n_949), .d(FE_OFN130_n_27449), .o(n_28515) );
oa22f80 g541752 ( .a(n_27571), .b(FE_OFN256_n_4280), .c(n_625), .d(FE_OFN102_n_27449), .o(n_28088) );
oa22f80 g541753 ( .a(n_27887), .b(FE_OFN313_n_3069), .c(n_1044), .d(FE_OFN131_n_27449), .o(n_28318) );
oa22f80 g541754 ( .a(n_27886), .b(FE_OFN269_n_4280), .c(n_1319), .d(FE_OFN90_n_27449), .o(n_28317) );
oa22f80 g541755 ( .a(n_26308), .b(n_4162), .c(n_806), .d(FE_OFN116_n_27449), .o(n_27209) );
oa22f80 g541756 ( .a(n_27738), .b(FE_OFN239_n_4162), .c(n_57), .d(FE_OFN135_n_27449), .o(n_28220) );
oa22f80 g541757 ( .a(FE_OFN937_n_27359), .b(n_27933), .c(n_1058), .d(FE_OFN1109_rst), .o(n_27934) );
oa22f80 g541758 ( .a(n_27735), .b(FE_OFN217_n_29687), .c(n_284), .d(FE_OFN1114_rst), .o(n_28219) );
oa22f80 g541759 ( .a(n_27734), .b(n_29687), .c(n_561), .d(FE_OFN101_n_27449), .o(n_28218) );
oa22f80 g541760 ( .a(n_26094), .b(FE_OFN1176_n_28597), .c(n_946), .d(FE_OFN1111_rst), .o(n_26452) );
oa22f80 g541761 ( .a(n_27733), .b(FE_OFN1177_n_28597), .c(n_1731), .d(FE_OFN113_n_27449), .o(n_28217) );
oa22f80 g541762 ( .a(n_27358), .b(FE_OFN6_n_28597), .c(n_889), .d(FE_OFN285_n_29266), .o(n_27932) );
oa22f80 g541763 ( .a(n_27730), .b(FE_OFN240_n_4162), .c(n_1416), .d(FE_OFN133_n_27449), .o(n_28216) );
oa22f80 g541764 ( .a(n_27729), .b(FE_OFN230_n_4162), .c(n_1891), .d(FE_OFN101_n_27449), .o(n_28215) );
oa22f80 g541765 ( .a(n_27884), .b(FE_OFN253_n_4280), .c(n_290), .d(FE_OFN21_n_27452), .o(n_28316) );
oa22f80 g541766 ( .a(n_27883), .b(FE_OFN312_n_3069), .c(n_584), .d(FE_OFN357_n_4860), .o(n_28315) );
oa22f80 g541767 ( .a(n_27885), .b(FE_OFN309_n_3069), .c(n_842), .d(FE_OFN364_n_4860), .o(n_28314) );
oa22f80 g541768 ( .a(n_27357), .b(FE_OFN409_n_28303), .c(n_154), .d(FE_OFN72_n_27012), .o(n_27931) );
oa22f80 g541769 ( .a(FE_OFN851_n_27728), .b(n_29664), .c(n_46), .d(FE_OFN347_n_4860), .o(n_28214) );
oa22f80 g541770 ( .a(n_27727), .b(FE_OFN411_n_28303), .c(n_1851), .d(FE_OFN335_n_4860), .o(n_28213) );
oa22f80 g541771 ( .a(n_27726), .b(n_28303), .c(n_1860), .d(n_27449), .o(n_28212) );
oa22f80 g541772 ( .a(n_27882), .b(FE_OFN258_n_4280), .c(n_1868), .d(FE_OFN1117_rst), .o(n_28312) );
oa22f80 g541773 ( .a(FE_OFN1009_n_27881), .b(n_22960), .c(n_458), .d(FE_OFN114_n_27449), .o(n_28310) );
oa22f80 g541774 ( .a(n_25848), .b(FE_OFN265_n_4280), .c(n_476), .d(FE_OFN115_n_27449), .o(n_26178) );
oa22f80 g541775 ( .a(n_25600), .b(FE_OFN235_n_4162), .c(n_1347), .d(n_29264), .o(n_25931) );
oa22f80 g541776 ( .a(n_27725), .b(FE_OFN294_n_3069), .c(n_445), .d(FE_OFN100_n_27449), .o(n_28210) );
oa22f80 g541777 ( .a(n_26443), .b(FE_OFN295_n_3069), .c(n_1372), .d(FE_OFN360_n_4860), .o(n_26444) );
oa22f80 g541778 ( .a(n_27231), .b(FE_OFN295_n_3069), .c(n_981), .d(FE_OFN100_n_27449), .o(n_27208) );
oa22f80 g541779 ( .a(n_28121), .b(FE_OFN313_n_3069), .c(n_843), .d(FE_OFN361_n_4860), .o(n_28513) );
oa22f80 g541780 ( .a(n_27569), .b(FE_OFN307_n_3069), .c(n_1672), .d(FE_OFN355_n_4860), .o(n_28087) );
oa22f80 g541781 ( .a(FE_OFN853_n_27880), .b(n_21076), .c(n_1306), .d(n_27449), .o(n_28308) );
oa22f80 g541782 ( .a(n_25846), .b(FE_OFN239_n_4162), .c(n_691), .d(FE_OFN350_n_4860), .o(n_26170) );
oa22f80 g541783 ( .a(n_27724), .b(FE_OFN240_n_4162), .c(n_1492), .d(FE_OFN352_n_4860), .o(n_28209) );
oa22f80 g541784 ( .a(n_27723), .b(FE_OFN417_n_28303), .c(n_1510), .d(FE_OFN131_n_27449), .o(n_28208) );
oa22f80 g541785 ( .a(n_27879), .b(FE_OFN235_n_4162), .c(n_700), .d(FE_OFN114_n_27449), .o(n_28306) );
oa22f80 g541786 ( .a(n_27878), .b(n_28303), .c(n_1152), .d(n_27449), .o(n_28304) );
oa22f80 g541787 ( .a(n_27568), .b(n_4162), .c(n_559), .d(FE_OFN353_n_4860), .o(n_28086) );
oa22f80 g541788 ( .a(n_27156), .b(FE_OFN417_n_28303), .c(n_1850), .d(FE_OFN361_n_4860), .o(n_27791) );
oa22f80 g541789 ( .a(n_27567), .b(FE_OFN240_n_4162), .c(n_608), .d(FE_OFN133_n_27449), .o(n_28085) );
oa22f80 g541790 ( .a(n_27877), .b(FE_OFN414_n_28303), .c(n_385), .d(FE_OFN326_n_4860), .o(n_28302) );
oa22f80 g541791 ( .a(n_25803), .b(FE_OFN253_n_4280), .c(n_997), .d(FE_OFN141_n_27449), .o(n_26679) );
oa22f80 g541792 ( .a(n_27564), .b(FE_OFN258_n_4280), .c(n_606), .d(FE_OFN141_n_27449), .o(n_28083) );
oa22f80 g541793 ( .a(n_28004), .b(FE_OFN410_n_28303), .c(n_620), .d(n_29204), .o(n_28398) );
oa22f80 g541794 ( .a(n_27356), .b(FE_OFN7_n_28597), .c(n_316), .d(FE_OFN11_n_29204), .o(n_27930) );
oa22f80 g541795 ( .a(n_27355), .b(n_28597), .c(n_311), .d(FE_OFN98_n_27449), .o(n_27928) );
oa22f80 g541796 ( .a(n_27876), .b(FE_OFN310_n_3069), .c(n_434), .d(FE_OFN115_n_27449), .o(n_28301) );
oa22f80 g541797 ( .a(n_27874), .b(FE_OFN299_n_3069), .c(n_543), .d(FE_OFN74_n_27012), .o(n_28299) );
oa22f80 g541798 ( .a(n_25528), .b(FE_OFN310_n_3069), .c(n_1660), .d(FE_OFN1143_n_27012), .o(n_26437) );
oa22f80 g541799 ( .a(n_27873), .b(FE_OFN297_n_3069), .c(n_1374), .d(FE_OFN285_n_29266), .o(n_28298) );
oa22f80 g541800 ( .a(n_28000), .b(FE_OFN311_n_3069), .c(n_213), .d(FE_OFN1171_n_4860), .o(n_28397) );
oa22f80 g541801 ( .a(n_25527), .b(FE_OFN150_n_25677), .c(n_783), .d(FE_OFN114_n_27449), .o(n_26436) );
oa22f80 g541802 ( .a(n_27871), .b(FE_OFN414_n_28303), .c(n_224), .d(FE_OFN90_n_27449), .o(n_28297) );
oa22f80 g541803 ( .a(n_27869), .b(n_4280), .c(n_121), .d(FE_OFN286_n_29266), .o(n_28295) );
oa22f80 g541804 ( .a(n_25802), .b(FE_OFN295_n_3069), .c(n_692), .d(FE_OFN100_n_27449), .o(n_26675) );
oa22f80 g541805 ( .a(n_27722), .b(FE_OFN203_n_28771), .c(n_84), .d(FE_OFN100_n_27449), .o(n_28207) );
oa22f80 g541806 ( .a(n_25801), .b(FE_OFN309_n_3069), .c(n_81), .d(FE_OFN128_n_27449), .o(n_26672) );
oa22f80 g541807 ( .a(n_27999), .b(FE_OFN311_n_3069), .c(n_263), .d(FE_OFN134_n_27449), .o(n_28396) );
oa22f80 g541808 ( .a(n_27870), .b(FE_OFN412_n_28303), .c(n_197), .d(FE_OFN119_n_27449), .o(n_28294) );
oa22f80 g541809 ( .a(n_25525), .b(FE_OFN259_n_4280), .c(n_723), .d(FE_OFN136_n_27449), .o(n_26434) );
oa22f80 g541810 ( .a(n_26925), .b(FE_OFN7_n_28597), .c(n_66), .d(FE_OFN360_n_4860), .o(n_27614) );
oa22f80 g541811 ( .a(n_27354), .b(FE_OFN7_n_28597), .c(n_998), .d(FE_OFN134_n_27449), .o(n_27927) );
oa22f80 g541812 ( .a(n_27721), .b(FE_OFN156_n_28014), .c(n_243), .d(FE_OFN91_n_27449), .o(n_28206) );
oa22f80 g541813 ( .a(n_32744), .b(x_in_36_14), .c(n_27231), .d(n_29194), .o(n_28941) );
in01f80 g541814 ( .a(n_27270), .o(n_27269) );
oa22f80 g541815 ( .a(n_25807), .b(n_13763), .c(n_13351), .d(n_13350), .o(n_27270) );
no02f80 g541904 ( .a(n_25688), .b(n_10963), .o(n_25689) );
no02f80 g541905 ( .a(n_28081), .b(n_28080), .o(n_28082) );
na02f80 g541906 ( .a(n_26146), .b(x_in_58_13), .o(n_26807) );
in01f80 g541907 ( .a(n_26430), .o(n_26431) );
no02f80 g541908 ( .a(n_26146), .b(x_in_58_13), .o(n_26430) );
no02f80 g541909 ( .a(n_25963), .b(n_25686), .o(n_25687) );
no02f80 g541910 ( .a(n_28204), .b(n_28203), .o(n_28205) );
in01f80 g541911 ( .a(n_27250), .o(n_26978) );
na02f80 g541912 ( .a(n_26670), .b(x_in_60_12), .o(n_27250) );
no02f80 g541913 ( .a(n_28201), .b(n_28200), .o(n_28202) );
na02f80 g541914 ( .a(n_26144), .b(x_in_2_12), .o(n_26804) );
in01f80 g541915 ( .a(n_26428), .o(n_26429) );
no02f80 g541916 ( .a(n_26144), .b(x_in_2_12), .o(n_26428) );
in01f80 g541917 ( .a(n_28738), .o(n_26977) );
no02f80 g541918 ( .a(n_26670), .b(x_in_60_12), .o(n_28738) );
no02f80 g541919 ( .a(n_28196), .b(n_28195), .o(n_28197) );
na02f80 g541920 ( .a(n_26426), .b(x_in_34_12), .o(n_27026) );
in01f80 g541921 ( .a(n_26668), .o(n_26669) );
no02f80 g541922 ( .a(n_26426), .b(x_in_34_12), .o(n_26668) );
na02f80 g541923 ( .a(n_26217), .b(n_25910), .o(n_26515) );
no02f80 g541924 ( .a(n_28193), .b(n_28192), .o(n_28194) );
na02f80 g541925 ( .a(n_26424), .b(x_in_18_12), .o(n_27025) );
in01f80 g541926 ( .a(n_26666), .o(n_26667) );
no02f80 g541927 ( .a(n_26424), .b(x_in_18_12), .o(n_26666) );
no02f80 g541928 ( .a(n_28190), .b(n_28189), .o(n_28191) );
na02f80 g541929 ( .a(n_26423), .b(x_in_50_12), .o(n_27024) );
in01f80 g541930 ( .a(n_26664), .o(n_26665) );
no02f80 g541931 ( .a(n_26423), .b(x_in_50_12), .o(n_26664) );
no02f80 g541932 ( .a(n_28077), .b(n_28076), .o(n_28078) );
na02f80 g541933 ( .a(n_26142), .b(x_in_10_12), .o(n_26801) );
in01f80 g541934 ( .a(n_26421), .o(n_26422) );
no02f80 g541935 ( .a(n_26142), .b(x_in_10_12), .o(n_26421) );
no02f80 g541936 ( .a(n_27924), .b(n_27923), .o(n_27925) );
na02f80 g541937 ( .a(n_26420), .b(x_in_6_12), .o(n_27023) );
in01f80 g541938 ( .a(n_26662), .o(n_26663) );
no02f80 g541939 ( .a(n_26420), .b(x_in_6_12), .o(n_26662) );
no02f80 g541940 ( .a(n_26216), .b(n_25905), .o(n_25906) );
no02f80 g541941 ( .a(n_28074), .b(n_28073), .o(n_28075) );
na02f80 g541942 ( .a(n_26140), .b(x_in_42_12), .o(n_26798) );
in01f80 g541943 ( .a(n_26418), .o(n_26419) );
no02f80 g541944 ( .a(n_26140), .b(x_in_42_12), .o(n_26418) );
no02f80 g541945 ( .a(n_28071), .b(n_28070), .o(n_28072) );
na02f80 g541946 ( .a(n_26139), .b(x_in_26_12), .o(n_26797) );
in01f80 g541947 ( .a(n_26416), .o(n_26417) );
no02f80 g541948 ( .a(n_26139), .b(x_in_26_12), .o(n_26416) );
no02f80 g541949 ( .a(n_28068), .b(n_28067), .o(n_28069) );
na02f80 g541950 ( .a(n_26414), .b(x_in_58_12), .o(n_27022) );
in01f80 g541951 ( .a(n_26660), .o(n_26661) );
no02f80 g541952 ( .a(n_26414), .b(x_in_58_12), .o(n_26660) );
no02f80 g541953 ( .a(n_27786), .b(n_27785), .o(n_27787) );
na02f80 g541954 ( .a(n_26413), .b(x_in_6_11), .o(n_27021) );
in01f80 g541955 ( .a(n_26658), .o(n_26659) );
no02f80 g541956 ( .a(n_26413), .b(x_in_6_11), .o(n_26658) );
in01f80 g541957 ( .a(n_26975), .o(n_26976) );
na02f80 g541958 ( .a(n_26657), .b(n_26046), .o(n_26975) );
no02f80 g541959 ( .a(n_28065), .b(n_28064), .o(n_28066) );
na02f80 g541960 ( .a(n_26412), .b(x_in_22_12), .o(n_27020) );
in01f80 g541961 ( .a(n_26655), .o(n_26656) );
no02f80 g541962 ( .a(n_26412), .b(x_in_22_12), .o(n_26655) );
no02f80 g541963 ( .a(n_28062), .b(n_28061), .o(n_28063) );
na02f80 g541964 ( .a(n_26138), .b(x_in_54_12), .o(n_26795) );
in01f80 g541965 ( .a(n_26410), .o(n_26411) );
no02f80 g541966 ( .a(n_26138), .b(x_in_54_12), .o(n_26410) );
no02f80 g541967 ( .a(n_28187), .b(n_28186), .o(n_28188) );
na02f80 g541968 ( .a(n_26409), .b(x_in_40_12), .o(n_27019) );
in01f80 g541969 ( .a(n_26653), .o(n_26654) );
no02f80 g541970 ( .a(n_26409), .b(x_in_40_12), .o(n_26653) );
no02f80 g541971 ( .a(n_28184), .b(n_28183), .o(n_28185) );
na02f80 g541972 ( .a(n_26408), .b(x_in_22_13), .o(n_27018) );
in01f80 g541973 ( .a(n_26651), .o(n_26652) );
no02f80 g541974 ( .a(n_26408), .b(x_in_22_13), .o(n_26651) );
no02f80 g541975 ( .a(n_28179), .b(n_28178), .o(n_28180) );
na02f80 g541976 ( .a(n_26136), .b(x_in_2_13), .o(n_26793) );
no02f80 g541977 ( .a(n_27781), .b(n_27780), .o(n_27782) );
na02f80 g541978 ( .a(n_26137), .b(x_in_14_12), .o(n_26792) );
in01f80 g541979 ( .a(n_26406), .o(n_26407) );
no02f80 g541980 ( .a(n_26137), .b(x_in_14_12), .o(n_26406) );
in01f80 g541981 ( .a(n_26404), .o(n_26405) );
no02f80 g541982 ( .a(n_26136), .b(x_in_2_13), .o(n_26404) );
no02f80 g541983 ( .a(n_27778), .b(n_27777), .o(n_27779) );
na02f80 g541984 ( .a(n_25847), .b(x_in_52_12), .o(n_26235) );
no02f80 g541985 ( .a(n_28058), .b(n_28057), .o(n_28059) );
na02f80 g541986 ( .a(n_26135), .b(x_in_46_12), .o(n_26791) );
in01f80 g541987 ( .a(n_26402), .o(n_26403) );
no02f80 g541988 ( .a(n_26135), .b(x_in_46_12), .o(n_26402) );
in01f80 g541989 ( .a(n_25890), .o(n_25891) );
no02f80 g541990 ( .a(n_25847), .b(x_in_52_12), .o(n_25890) );
no02f80 g541991 ( .a(n_28055), .b(n_28054), .o(n_28056) );
na02f80 g541992 ( .a(n_26133), .b(x_in_30_12), .o(n_26789) );
in01f80 g541993 ( .a(n_26400), .o(n_26401) );
no02f80 g541994 ( .a(n_26133), .b(x_in_30_12), .o(n_26400) );
na02f80 g541995 ( .a(n_25357), .b(n_25356), .o(n_25358) );
no02f80 g541996 ( .a(n_28052), .b(n_28051), .o(n_28053) );
na02f80 g541997 ( .a(n_26132), .b(x_in_62_12), .o(n_26788) );
in01f80 g541998 ( .a(n_26398), .o(n_26399) );
no02f80 g541999 ( .a(n_26132), .b(x_in_62_12), .o(n_26398) );
no02f80 g542000 ( .a(n_28175), .b(n_28174), .o(n_28176) );
na02f80 g542001 ( .a(n_26131), .b(x_in_54_13), .o(n_26787) );
in01f80 g542002 ( .a(n_26395), .o(n_26396) );
no02f80 g542003 ( .a(n_26131), .b(x_in_54_13), .o(n_26395) );
na02f80 g542004 ( .a(n_25357), .b(n_15840), .o(n_25729) );
no02f80 g542005 ( .a(n_28049), .b(n_28048), .o(n_28050) );
no02f80 g542006 ( .a(n_27921), .b(n_27920), .o(n_27922) );
na02f80 g542007 ( .a(n_26130), .b(x_in_14_13), .o(n_26786) );
in01f80 g542008 ( .a(n_26393), .o(n_26394) );
no02f80 g542009 ( .a(n_26130), .b(x_in_14_13), .o(n_26393) );
no02f80 g542010 ( .a(n_28387), .b(n_28386), .o(n_28388) );
na02f80 g542011 ( .a(n_26392), .b(x_in_34_13), .o(n_27017) );
in01f80 g542012 ( .a(n_26649), .o(n_26650) );
no02f80 g542013 ( .a(n_26392), .b(x_in_34_13), .o(n_26649) );
no02f80 g542014 ( .a(n_28171), .b(n_28170), .o(n_28172) );
na02f80 g542015 ( .a(n_26129), .b(x_in_46_13), .o(n_26784) );
in01f80 g542016 ( .a(n_26390), .o(n_26391) );
no02f80 g542017 ( .a(n_26129), .b(x_in_46_13), .o(n_26390) );
no02f80 g542018 ( .a(n_28044), .b(n_28043), .o(n_28045) );
na02f80 g542019 ( .a(n_26128), .b(x_in_16_13), .o(n_26781) );
in01f80 g542020 ( .a(n_26388), .o(n_26389) );
no02f80 g542021 ( .a(n_26128), .b(x_in_16_13), .o(n_26388) );
no02f80 g542022 ( .a(n_25660), .b(n_25659), .o(n_25661) );
no02f80 g542023 ( .a(n_28166), .b(n_28165), .o(n_28167) );
na02f80 g542024 ( .a(n_26126), .b(x_in_30_13), .o(n_26780) );
in01f80 g542025 ( .a(n_26386), .o(n_26387) );
no02f80 g542026 ( .a(n_26126), .b(x_in_30_13), .o(n_26386) );
no02f80 g542027 ( .a(n_28041), .b(n_28040), .o(n_28042) );
na02f80 g542028 ( .a(n_26125), .b(x_in_18_13), .o(n_26779) );
in01f80 g542029 ( .a(n_26384), .o(n_26385) );
no02f80 g542030 ( .a(n_26125), .b(x_in_18_13), .o(n_26384) );
no02f80 g542031 ( .a(n_28163), .b(n_28162), .o(n_28164) );
na02f80 g542032 ( .a(n_26124), .b(x_in_62_13), .o(n_26778) );
in01f80 g542033 ( .a(n_26382), .o(n_26383) );
no02f80 g542034 ( .a(n_26124), .b(x_in_62_13), .o(n_26382) );
no02f80 g542035 ( .a(n_27918), .b(n_27917), .o(n_27919) );
in01f80 g542036 ( .a(n_26647), .o(n_26648) );
no02f80 g542037 ( .a(n_26381), .b(x_in_12_13), .o(n_26647) );
no02f80 g542038 ( .a(n_27606), .b(n_27605), .o(n_27607) );
na02f80 g542039 ( .a(n_26381), .b(x_in_12_13), .o(n_27016) );
na02f80 g542040 ( .a(n_26123), .b(x_in_32_11), .o(n_26777) );
in01f80 g542041 ( .a(n_26379), .o(n_26380) );
no02f80 g542042 ( .a(n_26123), .b(x_in_32_11), .o(n_26379) );
no02f80 g542043 ( .a(n_27915), .b(n_27914), .o(n_27916) );
na02f80 g542044 ( .a(n_26378), .b(x_in_16_12), .o(n_27015) );
in01f80 g542045 ( .a(n_26645), .o(n_26646) );
no02f80 g542046 ( .a(n_26378), .b(x_in_16_12), .o(n_26645) );
no02f80 g542047 ( .a(n_28160), .b(n_28159), .o(n_28161) );
na02f80 g542048 ( .a(n_26119), .b(x_in_50_13), .o(n_26776) );
in01f80 g542049 ( .a(n_26376), .o(n_26377) );
no02f80 g542050 ( .a(n_26119), .b(x_in_50_13), .o(n_26376) );
na02f80 g542051 ( .a(n_26974), .b(x_in_48_11), .o(n_27443) );
in01f80 g542052 ( .a(n_27203), .o(n_27204) );
no02f80 g542053 ( .a(n_26974), .b(x_in_48_11), .o(n_27203) );
in01f80 g542054 ( .a(n_28157), .o(n_28158) );
na02f80 g542055 ( .a(n_28029), .b(n_27744), .o(n_28157) );
no02f80 g542056 ( .a(n_27774), .b(n_27773), .o(n_27775) );
na02f80 g542057 ( .a(n_26644), .b(x_in_40_11), .o(n_27247) );
in01f80 g542058 ( .a(n_26972), .o(n_26973) );
no02f80 g542059 ( .a(n_26644), .b(x_in_40_11), .o(n_26972) );
no02f80 g542060 ( .a(n_27771), .b(n_27770), .o(n_27772) );
in01f80 g542061 ( .a(n_26520), .o(n_26118) );
na02f80 g542062 ( .a(n_26078), .b(x_in_32_12), .o(n_26520) );
in01f80 g542063 ( .a(n_28431), .o(n_26117) );
no02f80 g542064 ( .a(n_26078), .b(x_in_32_12), .o(n_28431) );
in01f80 g542065 ( .a(n_27603), .o(n_27604) );
na02f80 g542066 ( .a(n_26942), .b(n_27394), .o(n_27603) );
no02f80 g542067 ( .a(n_28155), .b(n_28154), .o(n_28156) );
na02f80 g542068 ( .a(n_26116), .b(x_in_10_13), .o(n_26775) );
in01f80 g542069 ( .a(n_26374), .o(n_26375) );
no02f80 g542070 ( .a(n_26116), .b(x_in_10_13), .o(n_26374) );
no02f80 g542071 ( .a(n_25688), .b(n_25654), .o(n_25655) );
in01f80 g542072 ( .a(n_27246), .o(n_26971) );
na02f80 g542073 ( .a(n_26643), .b(x_in_48_12), .o(n_27246) );
in01f80 g542074 ( .a(n_28776), .o(n_26970) );
no02f80 g542075 ( .a(n_26643), .b(x_in_48_12), .o(n_28776) );
no02f80 g542076 ( .a(n_28286), .b(n_28285), .o(n_28287) );
in01f80 g542077 ( .a(n_27201), .o(n_27202) );
no02f80 g542078 ( .a(n_26969), .b(x_in_20_12), .o(n_27201) );
no02f80 g542079 ( .a(n_28152), .b(n_28151), .o(n_28153) );
na02f80 g542080 ( .a(n_26115), .b(x_in_42_13), .o(n_26772) );
na02f80 g542081 ( .a(n_26969), .b(x_in_20_12), .o(n_27440) );
in01f80 g542082 ( .a(n_26372), .o(n_26373) );
no02f80 g542083 ( .a(n_26115), .b(x_in_42_13), .o(n_26372) );
no02f80 g542084 ( .a(n_28027), .b(n_28026), .o(n_28028) );
na02f80 g542085 ( .a(n_26968), .b(x_in_36_11), .o(n_27439) );
in01f80 g542086 ( .a(n_27199), .o(n_27200) );
no02f80 g542087 ( .a(n_26968), .b(x_in_36_11), .o(n_27199) );
no02f80 g542088 ( .a(n_26443), .b(n_26113), .o(n_26114) );
in01f80 g542089 ( .a(n_26224), .o(n_26112) );
no02f80 g542090 ( .a(n_25526), .b(n_26113), .o(n_26224) );
no02f80 g542091 ( .a(n_28283), .b(n_28282), .o(n_28284) );
na02f80 g542092 ( .a(n_27198), .b(x_in_20_11), .o(n_27644) );
in01f80 g542093 ( .a(n_27392), .o(n_27393) );
no02f80 g542094 ( .a(n_27198), .b(x_in_20_11), .o(n_27392) );
no02f80 g542095 ( .a(n_26459), .b(n_26110), .o(n_26111) );
in01f80 g542096 ( .a(n_26221), .o(n_26109) );
no02f80 g542097 ( .a(n_25529), .b(n_26110), .o(n_26221) );
no02f80 g542098 ( .a(n_27390), .b(n_27389), .o(n_27391) );
na02f80 g542099 ( .a(n_25873), .b(x_in_52_11), .o(n_26518) );
in01f80 g542100 ( .a(n_26107), .o(n_26108) );
no02f80 g542101 ( .a(n_25873), .b(x_in_52_11), .o(n_26107) );
no02f80 g542102 ( .a(n_28149), .b(n_28148), .o(n_28150) );
na02f80 g542103 ( .a(n_26106), .b(x_in_26_13), .o(n_26768) );
in01f80 g542104 ( .a(n_26370), .o(n_26371) );
no02f80 g542105 ( .a(n_26106), .b(x_in_26_13), .o(n_26370) );
no02f80 g542106 ( .a(n_27768), .b(n_27767), .o(n_27769) );
na02f80 g542107 ( .a(n_26369), .b(x_in_12_12), .o(n_27013) );
in01f80 g542108 ( .a(n_26641), .o(n_26642) );
no02f80 g542109 ( .a(n_26369), .b(x_in_12_12), .o(n_26641) );
in01f80 g542110 ( .a(n_27387), .o(n_27388) );
no02f80 g542111 ( .a(n_27197), .b(x_in_44_14), .o(n_27387) );
na02f80 g542112 ( .a(n_27197), .b(x_in_44_14), .o(n_27643) );
na02f80 g542113 ( .a(n_27197), .b(x_in_44_15), .o(n_27196) );
in01f80 g542114 ( .a(n_26966), .o(n_26967) );
na02f80 g542115 ( .a(n_26640), .b(n_26027), .o(n_26966) );
no02f80 g542116 ( .a(n_28146), .b(n_28145), .o(n_28147) );
na02f80 g542117 ( .a(n_26639), .b(x_in_60_11), .o(n_27244) );
in01f80 g542118 ( .a(n_26964), .o(n_26965) );
no02f80 g542119 ( .a(n_26639), .b(x_in_60_11), .o(n_26964) );
no02f80 g542120 ( .a(n_25634), .b(n_25633), .o(n_25635) );
na02f80 g542121 ( .a(n_27231), .b(n_26962), .o(n_26963) );
oa22f80 g542122 ( .a(n_24562), .b(n_12664), .c(n_24183), .d(n_12056), .o(n_26260) );
na02f80 g542123 ( .a(n_26104), .b(n_26103), .o(n_26105) );
no02f80 g542124 ( .a(n_26104), .b(n_16496), .o(n_26102) );
na02f80 g542125 ( .a(n_25966), .b(n_25631), .o(n_25632) );
no02f80 g542126 ( .a(n_25629), .b(n_25628), .o(n_25630) );
in01f80 g542127 ( .a(n_25626), .o(n_25627) );
ao12f80 g542128 ( .a(n_24594), .b(n_24197), .c(n_9339), .o(n_25626) );
no02f80 g542129 ( .a(n_25871), .b(n_25870), .o(n_25872) );
na02f80 g542130 ( .a(n_32744), .b(x_in_36_13), .o(n_27241) );
na02f80 g542131 ( .a(n_26501), .b(n_26100), .o(n_26101) );
no02f80 g542132 ( .a(n_25938), .b(n_25621), .o(n_25622) );
no02f80 g542133 ( .a(n_25936), .b(n_25619), .o(n_25620) );
no02f80 g542134 ( .a(n_28234), .b(n_28024), .o(n_28025) );
na02f80 g542135 ( .a(n_26637), .b(n_26610), .o(n_26638) );
in01f80 g542136 ( .a(n_26960), .o(n_26961) );
no02f80 g542137 ( .a(n_32744), .b(x_in_36_12), .o(n_26960) );
na02f80 g542138 ( .a(n_32744), .b(x_in_36_12), .o(n_28650) );
na02f80 g542139 ( .a(n_25964), .b(n_25612), .o(n_25613) );
no02f80 g542140 ( .a(n_25935), .b(n_25607), .o(n_25608) );
no02f80 g542141 ( .a(n_25605), .b(n_25604), .o(n_25606) );
no02f80 g542142 ( .a(n_25602), .b(n_25601), .o(n_25603) );
in01f80 g542143 ( .a(n_26764), .o(n_26368) );
no02f80 g542144 ( .a(n_25534), .b(n_25532), .o(n_26764) );
no02f80 g542145 ( .a(n_25868), .b(n_25867), .o(n_25869) );
in01f80 g542146 ( .a(n_26943), .o(n_25866) );
na02f80 g542147 ( .a(n_25600), .b(n_25867), .o(n_26943) );
in01f80 g542148 ( .a(FE_OFN901_n_26098), .o(n_26099) );
oa12f80 g542149 ( .a(n_25228), .b(n_2871), .c(x_in_49_14), .o(n_26098) );
na02f80 g542150 ( .a(n_26307), .b(FE_OFN1124_rst), .o(n_27432) );
na02f80 g542151 ( .a(n_26018), .b(FE_OFN1114_rst), .o(n_27236) );
na02f80 g542152 ( .a(n_27197), .b(FE_OFN290_n_27194), .o(n_27639) );
in01f80 g542153 ( .a(n_26636), .o(n_27082) );
na02f80 g542154 ( .a(n_26019), .b(n_26627), .o(n_26636) );
no02f80 g542155 ( .a(n_26366), .b(n_26365), .o(n_26367) );
na02f80 g542156 ( .a(n_26094), .b(n_26365), .o(n_26762) );
na02f80 g542157 ( .a(n_26092), .b(n_26091), .o(n_26093) );
na02f80 g542158 ( .a(n_26092), .b(n_25441), .o(n_26868) );
na02f80 g542159 ( .a(n_26363), .b(n_26362), .o(n_26364) );
na02f80 g542160 ( .a(n_26363), .b(n_25756), .o(n_27078) );
na02f80 g542161 ( .a(n_25864), .b(n_26090), .o(n_25865) );
in01f80 g542162 ( .a(n_26361), .o(n_26863) );
no02f80 g542163 ( .a(n_26125), .b(n_26090), .o(n_26361) );
na02f80 g542164 ( .a(n_25862), .b(n_26089), .o(n_25863) );
in01f80 g542165 ( .a(n_26360), .o(n_26860) );
no02f80 g542166 ( .a(n_26119), .b(n_26089), .o(n_26360) );
na02f80 g542167 ( .a(n_26358), .b(n_26313), .o(n_26359) );
na02f80 g542168 ( .a(n_26087), .b(n_26086), .o(n_26088) );
na02f80 g542169 ( .a(n_26087), .b(n_25437), .o(n_26859) );
na02f80 g542170 ( .a(n_26084), .b(n_26083), .o(n_26085) );
na02f80 g542171 ( .a(n_26084), .b(n_25436), .o(n_26858) );
na02f80 g542172 ( .a(n_26081), .b(n_26080), .o(n_26082) );
na02f80 g542173 ( .a(n_26081), .b(n_25435), .o(n_26857) );
na02f80 g542174 ( .a(n_25860), .b(n_26079), .o(n_25861) );
in01f80 g542175 ( .a(n_26357), .o(n_26854) );
no02f80 g542176 ( .a(n_26146), .b(n_26079), .o(n_26357) );
na02f80 g542177 ( .a(n_26420), .b(n_26355), .o(n_26356) );
in01f80 g542178 ( .a(n_26851), .o(n_26354) );
na02f80 g542179 ( .a(n_25804), .b(n_26355), .o(n_26851) );
oa12f80 g542180 ( .a(n_26953), .b(n_1695), .c(FE_OFN60_n_27012), .o(n_26955) );
oa12f80 g542181 ( .a(n_26953), .b(n_172), .c(FE_OFN129_n_27449), .o(n_26954) );
na02f80 g542182 ( .a(n_26078), .b(n_25856), .o(n_25857) );
no02f80 g542183 ( .a(n_26078), .b(n_25433), .o(n_26848) );
na02f80 g542184 ( .a(n_25854), .b(n_26077), .o(n_25855) );
in01f80 g542185 ( .a(n_26353), .o(n_26844) );
no02f80 g542186 ( .a(n_26128), .b(n_26077), .o(n_26353) );
oa12f80 g542187 ( .a(n_26633), .b(n_1939), .c(FE_OFN138_n_27449), .o(n_26635) );
oa12f80 g542188 ( .a(n_26633), .b(n_301), .c(FE_OFN78_n_27012), .o(n_26634) );
na02f80 g542189 ( .a(n_26351), .b(n_26632), .o(n_26352) );
no02f80 g542190 ( .a(n_26643), .b(n_26632), .o(n_27262) );
na02f80 g542191 ( .a(n_26075), .b(n_26350), .o(n_26076) );
in01f80 g542192 ( .a(n_27162), .o(n_26631) );
no02f80 g542193 ( .a(n_26409), .b(n_26350), .o(n_27162) );
no02f80 g542194 ( .a(n_26073), .b(n_26072), .o(n_26074) );
in01f80 g542195 ( .a(n_26071), .o(n_26559) );
na02f80 g542196 ( .a(n_25848), .b(n_26072), .o(n_26071) );
na02f80 g542197 ( .a(n_26629), .b(n_27211), .o(n_26630) );
na02f80 g542198 ( .a(n_25847), .b(n_25569), .o(n_25570) );
no02f80 g542199 ( .a(n_25847), .b(n_25145), .o(n_26926) );
no02f80 g542200 ( .a(n_26069), .b(n_26068), .o(n_26070) );
in01f80 g542201 ( .a(n_26067), .o(n_26556) );
na02f80 g542202 ( .a(n_25846), .b(n_26068), .o(n_26067) );
na02f80 g542203 ( .a(n_26670), .b(n_26627), .o(n_26628) );
in01f80 g542204 ( .a(n_28473), .o(n_28385) );
oa12f80 g542205 ( .a(n_26025), .b(n_27850), .c(n_25511), .o(n_28473) );
in01f80 g542206 ( .a(n_28589), .o(n_28737) );
oa12f80 g542207 ( .a(n_26616), .b(n_26010), .c(n_27983), .o(n_28589) );
in01f80 g542208 ( .a(n_28592), .o(n_28510) );
oa12f80 g542209 ( .a(n_26326), .b(n_25790), .c(n_27982), .o(n_28592) );
oa12f80 g542210 ( .a(n_26624), .b(n_1466), .c(FE_OFN134_n_27449), .o(n_26626) );
oa12f80 g542211 ( .a(n_26624), .b(n_1387), .c(FE_OFN134_n_27449), .o(n_26625) );
in01f80 g542212 ( .a(n_28586), .o(n_28509) );
oa12f80 g542213 ( .a(n_26615), .b(n_26008), .c(n_27981), .o(n_28586) );
in01f80 g542214 ( .a(n_28583), .o(n_28508) );
oa12f80 g542215 ( .a(n_26049), .b(n_25508), .c(n_27980), .o(n_28583) );
oa12f80 g542216 ( .a(n_25816), .b(n_26021), .c(n_24807), .o(n_26349) );
in01f80 g542217 ( .a(n_28580), .o(n_28507) );
oa12f80 g542218 ( .a(n_26048), .b(n_25506), .c(n_27979), .o(n_28580) );
in01f80 g542219 ( .a(n_28470), .o(n_28384) );
oa12f80 g542220 ( .a(n_26324), .b(n_27849), .c(n_25787), .o(n_28470) );
in01f80 g542221 ( .a(n_28351), .o(n_28281) );
oa12f80 g542222 ( .a(n_26325), .b(n_25785), .c(n_27671), .o(n_28351) );
in01f80 g542223 ( .a(n_28467), .o(n_28383) );
oa12f80 g542224 ( .a(n_26323), .b(n_27848), .c(n_25783), .o(n_28467) );
in01f80 g542225 ( .a(n_28464), .o(n_28382) );
oa12f80 g542226 ( .a(n_26322), .b(n_27847), .c(n_25781), .o(n_28464) );
in01f80 g542227 ( .a(n_28461), .o(n_28381) );
oa12f80 g542228 ( .a(n_26047), .b(n_27846), .c(n_25500), .o(n_28461) );
in01f80 g542229 ( .a(n_28255), .o(n_28142) );
oa12f80 g542230 ( .a(n_26614), .b(n_26006), .c(n_27484), .o(n_28255) );
in01f80 g542231 ( .a(n_28380), .o(n_28648) );
oa12f80 g542232 ( .a(n_25076), .b(n_24392), .c(n_28271), .o(n_28380) );
in01f80 g542233 ( .a(n_28280), .o(n_28538) );
oa12f80 g542234 ( .a(n_25075), .b(n_24390), .c(n_28136), .o(n_28280) );
in01f80 g542235 ( .a(n_28458), .o(n_28379) );
oa12f80 g542236 ( .a(n_26321), .b(n_25775), .c(n_27844), .o(n_28458) );
in01f80 g542237 ( .a(n_28455), .o(n_28378) );
oa12f80 g542238 ( .a(n_26044), .b(n_25496), .c(n_27843), .o(n_28455) );
in01f80 g542239 ( .a(n_28449), .o(n_28377) );
oa12f80 g542240 ( .a(n_26030), .b(n_25485), .c(n_27840), .o(n_28449) );
in01f80 g542241 ( .a(n_28577), .o(n_28506) );
oa12f80 g542242 ( .a(n_26320), .b(n_25773), .c(n_27978), .o(n_28577) );
in01f80 g542243 ( .a(n_28574), .o(n_28505) );
ao12f80 g542244 ( .a(n_25493), .b(n_26042), .c(n_27977), .o(n_28574) );
in01f80 g542245 ( .a(n_28571), .o(n_28504) );
oa12f80 g542246 ( .a(n_26043), .b(n_25491), .c(n_27976), .o(n_28571) );
in01f80 g542247 ( .a(n_28251), .o(n_28141) );
oa12f80 g542248 ( .a(n_26041), .b(n_25489), .c(n_27480), .o(n_28251) );
in01f80 g542249 ( .a(n_28452), .o(n_28376) );
oa12f80 g542250 ( .a(n_26040), .b(n_25487), .c(n_27841), .o(n_28452) );
in01f80 g542251 ( .a(n_28248), .o(n_28140) );
oa12f80 g542252 ( .a(n_25829), .b(n_27481), .c(n_25217), .o(n_28248) );
in01f80 g542253 ( .a(n_28446), .o(n_28375) );
oa12f80 g542254 ( .a(n_26039), .b(n_25483), .c(n_27839), .o(n_28446) );
in01f80 g542255 ( .a(n_28568), .o(n_28503) );
ao12f80 g542256 ( .a(n_25212), .b(n_25828), .c(n_27975), .o(n_28568) );
in01f80 g542257 ( .a(n_28279), .o(n_28536) );
oa12f80 g542258 ( .a(n_23994), .b(n_28134), .c(n_23365), .o(n_28279) );
in01f80 g542259 ( .a(n_28525), .o(n_28374) );
oa12f80 g542260 ( .a(n_26940), .b(n_26303), .c(n_27838), .o(n_28525) );
in01f80 g542261 ( .a(n_28348), .o(n_28278) );
ao12f80 g542262 ( .a(n_25210), .b(n_25827), .c(n_27668), .o(n_28348) );
in01f80 g542263 ( .a(n_28760), .o(n_28710) );
oa12f80 g542264 ( .a(n_26318), .b(n_25771), .c(n_28239), .o(n_28760) );
in01f80 g542265 ( .a(n_28565), .o(n_28502) );
oa12f80 g542266 ( .a(n_25826), .b(n_25208), .c(n_27974), .o(n_28565) );
in01f80 g542267 ( .a(n_28441), .o(n_28373) );
oa12f80 g542268 ( .a(n_26038), .b(n_25481), .c(n_27837), .o(n_28441) );
in01f80 g542269 ( .a(n_28562), .o(n_28501) );
ao12f80 g542270 ( .a(n_25205), .b(n_25825), .c(n_27973), .o(n_28562) );
in01f80 g542271 ( .a(n_28438), .o(n_28372) );
oa12f80 g542272 ( .a(n_26037), .b(n_25479), .c(n_27836), .o(n_28438) );
in01f80 g542273 ( .a(n_28559), .o(n_28500) );
oa12f80 g542274 ( .a(n_25824), .b(n_25202), .c(n_27972), .o(n_28559) );
in01f80 g542275 ( .a(n_28101), .o(n_28017) );
oa12f80 g542276 ( .a(n_26317), .b(n_25769), .c(n_27276), .o(n_28101) );
in01f80 g542277 ( .a(n_28345), .o(n_28277) );
ao12f80 g542278 ( .a(n_25477), .b(n_26036), .c(n_27666), .o(n_28345) );
in01f80 g542279 ( .a(n_28342), .o(n_28276) );
oa12f80 g542280 ( .a(n_26035), .b(n_25474), .c(n_27665), .o(n_28342) );
in01f80 g542281 ( .a(n_28556), .o(n_28499) );
oa12f80 g542282 ( .a(n_26034), .b(n_25472), .c(n_27971), .o(n_28556) );
in01f80 g542283 ( .a(n_28243), .o(n_28139) );
oa12f80 g542284 ( .a(n_26316), .b(n_25766), .c(n_27478), .o(n_28243) );
in01f80 g542285 ( .a(n_28240), .o(n_28430) );
oa12f80 g542286 ( .a(n_26033), .b(n_25469), .c(n_27477), .o(n_28240) );
in01f80 g542287 ( .a(n_28371), .o(n_28646) );
oa12f80 g542288 ( .a(n_25929), .b(n_28269), .c(n_25303), .o(n_28371) );
in01f80 g542289 ( .a(n_28016), .o(n_28340) );
ao12f80 g542290 ( .a(n_23971), .b(n_27898), .c(n_24659), .o(n_28016) );
oa12f80 g542291 ( .a(n_11818), .b(n_25839), .c(n_13121), .o(n_26549) );
in01f80 g542292 ( .a(n_28553), .o(n_28498) );
oa12f80 g542293 ( .a(n_26032), .b(n_27967), .c(n_25467), .o(n_28553) );
in01f80 g542294 ( .a(n_28275), .o(n_28534) );
oa12f80 g542295 ( .a(n_24756), .b(n_24111), .c(n_28132), .o(n_28275) );
in01f80 g542296 ( .a(n_28663), .o(n_28632) );
oa12f80 g542297 ( .a(n_26935), .b(n_26291), .c(n_28100), .o(n_28663) );
in01f80 g542298 ( .a(n_28550), .o(n_28497) );
oa12f80 g542299 ( .a(n_26031), .b(n_27966), .c(n_25465), .o(n_28550) );
in01f80 g542300 ( .a(n_28435), .o(n_28370) );
oa12f80 g542301 ( .a(n_26934), .b(n_26289), .c(n_27832), .o(n_28435) );
in01f80 g542302 ( .a(n_28660), .o(n_28631) );
oa12f80 g542303 ( .a(n_26933), .b(n_26287), .c(n_28099), .o(n_28660) );
in01f80 g542304 ( .a(n_27968), .o(n_27900) );
oa12f80 g542305 ( .a(n_26028), .b(n_27085), .c(n_25457), .o(n_27968) );
in01f80 g542306 ( .a(n_28547), .o(n_28496) );
oa12f80 g542307 ( .a(n_26029), .b(n_27965), .c(n_25455), .o(n_28547) );
in01f80 g542308 ( .a(n_28236), .o(n_28138) );
oa12f80 g542309 ( .a(n_26315), .b(n_25762), .c(n_27476), .o(n_28236) );
in01f80 g542310 ( .a(n_28274), .o(n_28532) );
oa12f80 g542311 ( .a(n_26171), .b(n_28130), .c(n_25571), .o(n_28274) );
in01f80 g542312 ( .a(n_28273), .o(n_28530) );
oa12f80 g542313 ( .a(n_25055), .b(n_24372), .c(n_28128), .o(n_28273) );
oa12f80 g542314 ( .a(n_26017), .b(n_26309), .c(n_25050), .o(n_26621) );
in01f80 g542315 ( .a(n_28544), .o(n_28495) );
oa12f80 g542316 ( .a(n_26932), .b(n_26282), .c(n_27964), .o(n_28544) );
oa12f80 g542317 ( .a(n_26329), .b(n_1729), .c(FE_OFN100_n_27449), .o(n_26331) );
oa12f80 g542318 ( .a(n_26329), .b(n_264), .c(FE_OFN100_n_27449), .o(n_26330) );
oa12f80 g542319 ( .a(n_25517), .b(n_25536), .c(n_24137), .o(n_26051) );
oa12f80 g542320 ( .a(n_27166), .b(n_204), .c(FE_OFN98_n_27449), .o(n_27169) );
oa12f80 g542321 ( .a(n_27166), .b(n_1483), .c(FE_OFN329_n_4860), .o(n_27167) );
oa12f80 g542322 ( .a(n_24849), .b(n_25757), .c(n_26016), .o(n_26999) );
ao22s80 g542323 ( .a(n_25397), .b(n_27845), .c(n_25398), .d(n_28271), .o(n_28272) );
ao22s80 g542324 ( .a(n_25396), .b(n_28136), .c(n_25395), .d(n_27670), .o(n_28137) );
ao12f80 g542325 ( .a(n_25818), .b(n_28863), .c(n_25817), .o(n_29146) );
ao22s80 g542326 ( .a(n_27669), .b(n_24260), .c(n_28134), .d(n_24261), .o(n_28135) );
ao22s80 g542327 ( .a(n_28269), .b(n_26175), .c(n_27833), .d(n_26174), .o(n_28270) );
ao22s80 g542328 ( .a(n_27898), .b(n_24977), .c(n_27275), .d(n_24976), .o(n_27899) );
oa12f80 g542329 ( .a(n_26617), .b(n_26618), .c(x_in_44_15), .o(n_29195) );
ao12f80 g542330 ( .a(n_25815), .b(n_25814), .c(n_25813), .o(n_26328) );
in01f80 g542331 ( .a(n_26759), .o(n_27008) );
ao12f80 g542332 ( .a(n_25545), .b(n_25839), .c(n_25544), .o(n_26759) );
ao22s80 g542333 ( .a(n_25059), .b(n_28132), .c(n_25058), .d(n_27662), .o(n_28133) );
in01f80 g542334 ( .a(n_27456), .o(n_27444) );
no02f80 g542335 ( .a(n_32744), .b(n_25986), .o(n_27456) );
ao22s80 g542336 ( .a(n_28130), .b(n_26442), .c(n_27661), .d(n_26441), .o(n_28131) );
ao22s80 g542337 ( .a(n_25385), .b(n_28128), .c(n_25384), .d(n_27660), .o(n_28129) );
ao12f80 g542338 ( .a(n_25542), .b(n_28798), .c(n_25541), .o(n_29137) );
oa22f80 g542339 ( .a(n_27657), .b(FE_OFN266_n_4280), .c(n_1704), .d(FE_OFN347_n_4860), .o(n_28127) );
oa22f80 g542340 ( .a(n_27472), .b(FE_OFN157_n_28014), .c(n_412), .d(FE_OFN96_n_27449), .o(n_28015) );
oa22f80 g542341 ( .a(n_27470), .b(FE_OFN409_n_28303), .c(n_1754), .d(FE_OFN93_n_27449), .o(n_28013) );
oa22f80 g542342 ( .a(n_25423), .b(FE_OFN409_n_28303), .c(n_473), .d(FE_OFN72_n_27012), .o(n_26327) );
oa22f80 g542343 ( .a(n_27268), .b(FE_OFN260_n_4280), .c(n_663), .d(FE_OFN1120_rst), .o(n_27891) );
oa22f80 g542344 ( .a(n_27081), .b(FE_OFN410_n_28303), .c(n_1111), .d(FE_OFN76_n_27012), .o(n_27748) );
oa22f80 g542345 ( .a(n_27655), .b(FE_OFN312_n_3069), .c(n_551), .d(FE_OFN60_n_27012), .o(n_28126) );
oa22f80 g542346 ( .a(n_27080), .b(FE_OFN306_n_3069), .c(n_159), .d(FE_OFN93_n_27449), .o(n_27747) );
oa22f80 g542347 ( .a(n_25744), .b(FE_OFN409_n_28303), .c(n_830), .d(FE_OFN355_n_4860), .o(n_26620) );
oa22f80 g542348 ( .a(n_27468), .b(FE_OFN296_n_3069), .c(n_1707), .d(FE_OFN358_n_4860), .o(n_28012) );
oa22f80 g542349 ( .a(n_27466), .b(FE_OFN312_n_3069), .c(n_1884), .d(FE_OFN329_n_4860), .o(n_28011) );
oa22f80 g542350 ( .a(n_27464), .b(FE_OFN296_n_3069), .c(n_1170), .d(FE_OFN1123_rst), .o(n_28010) );
oa22f80 g542351 ( .a(n_26024), .b(n_1029), .c(n_26319), .d(x_in_2_15), .o(n_29294) );
in01f80 g542375 ( .a(n_26941), .o(n_26942) );
no02f80 g542376 ( .a(n_26618), .b(x_in_44_14), .o(n_26941) );
na02f80 g542377 ( .a(n_26618), .b(x_in_44_14), .o(n_27394) );
na02f80 g542378 ( .a(n_26618), .b(x_in_44_15), .o(n_26617) );
na02f80 g542379 ( .a(n_26616), .b(n_26011), .o(n_28204) );
na02f80 g542380 ( .a(n_26326), .b(n_25791), .o(n_28201) );
na02f80 g542381 ( .a(n_26615), .b(n_26009), .o(n_28196) );
na02f80 g542382 ( .a(n_26049), .b(n_25509), .o(n_28193) );
na02f80 g542383 ( .a(n_26048), .b(n_25507), .o(n_28190) );
na02f80 g542384 ( .a(n_26325), .b(n_25786), .o(n_27924) );
na02f80 g542385 ( .a(n_26324), .b(n_25788), .o(n_28077) );
na02f80 g542386 ( .a(n_26323), .b(n_25784), .o(n_28074) );
na02f80 g542387 ( .a(n_26322), .b(n_25782), .o(n_28071) );
na02f80 g542388 ( .a(n_26047), .b(n_25501), .o(n_28068) );
na02f80 g542389 ( .a(n_26614), .b(n_26007), .o(n_27786) );
na02f80 g542390 ( .a(n_25830), .b(x_in_38_14), .o(n_26657) );
in01f80 g542391 ( .a(n_26045), .o(n_26046) );
no02f80 g542392 ( .a(n_25830), .b(x_in_38_14), .o(n_26045) );
na02f80 g542393 ( .a(n_26321), .b(n_25776), .o(n_28065) );
na02f80 g542394 ( .a(n_26044), .b(n_25497), .o(n_28062) );
na02f80 g542395 ( .a(n_26320), .b(n_25774), .o(n_28187) );
na02f80 g542396 ( .a(n_26043), .b(n_25492), .o(n_28179) );
na02f80 g542397 ( .a(n_26042), .b(n_25494), .o(n_28184) );
na02f80 g542398 ( .a(n_25829), .b(n_25218), .o(n_27778) );
na02f80 g542399 ( .a(n_26041), .b(n_25490), .o(n_27781) );
na02f80 g542400 ( .a(n_26040), .b(n_25488), .o(n_28058) );
na02f80 g542401 ( .a(n_26039), .b(n_25484), .o(n_28052) );
na02f80 g542402 ( .a(n_25828), .b(n_25213), .o(n_28175) );
na02f80 g542403 ( .a(n_26319), .b(n_27194), .o(n_26953) );
na02f80 g542404 ( .a(n_26940), .b(n_26304), .o(n_28049) );
na02f80 g542405 ( .a(n_25827), .b(n_25211), .o(n_27921) );
na02f80 g542406 ( .a(n_26318), .b(n_25772), .o(n_28387) );
na02f80 g542407 ( .a(n_25826), .b(n_25209), .o(n_28171) );
na02f80 g542408 ( .a(n_26038), .b(n_25482), .o(n_28044) );
na02f80 g542409 ( .a(n_25825), .b(n_25206), .o(n_28166) );
na02f80 g542410 ( .a(n_26037), .b(n_25480), .o(n_28041) );
na02f80 g542411 ( .a(n_25824), .b(n_25203), .o(n_28163) );
na02f80 g542412 ( .a(n_26036), .b(n_25478), .o(n_27918) );
na02f80 g542413 ( .a(n_26317), .b(n_25770), .o(n_27606) );
na02f80 g542414 ( .a(n_26035), .b(n_25475), .o(n_27915) );
na02f80 g542415 ( .a(n_26034), .b(n_25473), .o(n_28160) );
in01f80 g542416 ( .a(n_26938), .o(n_26939) );
na02f80 g542417 ( .a(n_26613), .b(n_26002), .o(n_26938) );
na02f80 g542418 ( .a(n_27579), .b(x_in_8_14), .o(n_28029) );
in01f80 g542419 ( .a(n_27743), .o(n_27744) );
no02f80 g542420 ( .a(n_27579), .b(x_in_8_14), .o(n_27743) );
na02f80 g542421 ( .a(n_26316), .b(n_25767), .o(n_27774) );
na02f80 g542422 ( .a(n_26033), .b(n_25470), .o(n_27771) );
no02f80 g542423 ( .a(n_25839), .b(n_25544), .o(n_25545) );
in01f80 g542424 ( .a(n_27741), .o(n_27742) );
na02f80 g542425 ( .a(n_27578), .b(n_27131), .o(n_27741) );
in01f80 g542426 ( .a(n_27576), .o(n_27577) );
na02f80 g542427 ( .a(n_26922), .b(n_27364), .o(n_27576) );
in01f80 g542428 ( .a(n_27574), .o(n_27575) );
na02f80 g542429 ( .a(n_26920), .b(n_27363), .o(n_27574) );
na02f80 g542430 ( .a(n_26032), .b(n_25468), .o(n_28155) );
in01f80 g542431 ( .a(n_26936), .o(n_26937) );
na02f80 g542432 ( .a(n_26612), .b(n_26000), .o(n_26936) );
na02f80 g542433 ( .a(n_26935), .b(n_26292), .o(n_28286) );
na02f80 g542434 ( .a(n_26031), .b(n_25466), .o(n_28152) );
na02f80 g542435 ( .a(n_26934), .b(n_26290), .o(n_28027) );
na02f80 g542436 ( .a(n_26933), .b(n_26288), .o(n_28283) );
na02f80 g542437 ( .a(n_26030), .b(n_25486), .o(n_28055) );
na02f80 g542438 ( .a(n_26029), .b(n_25456), .o(n_28149) );
na02f80 g542439 ( .a(n_26028), .b(n_25458), .o(n_27390) );
na02f80 g542440 ( .a(n_26315), .b(n_25763), .o(n_27768) );
in01f80 g542441 ( .a(n_27572), .o(n_27573) );
na02f80 g542442 ( .a(n_27362), .b(n_26891), .o(n_27572) );
na02f80 g542443 ( .a(n_25822), .b(x_in_28_14), .o(n_26640) );
in01f80 g542444 ( .a(n_26026), .o(n_26027) );
no02f80 g542445 ( .a(n_25822), .b(x_in_28_14), .o(n_26026) );
na02f80 g542446 ( .a(n_26025), .b(n_25512), .o(n_28081) );
na02f80 g542447 ( .a(n_26932), .b(n_26283), .o(n_28146) );
na02f80 g542448 ( .a(n_25820), .b(n_25819), .o(n_25821) );
no02f80 g542449 ( .a(n_26610), .b(FE_OFN23_n_26609), .o(n_26611) );
na02f80 g542450 ( .a(n_26618), .b(FE_OFN290_n_27194), .o(n_27166) );
no02f80 g542451 ( .a(n_28798), .b(n_25541), .o(n_25542) );
no02f80 g542452 ( .a(n_28863), .b(n_25817), .o(n_25818) );
no02f80 g542453 ( .a(n_26313), .b(FE_OFN369_n_26312), .o(n_26314) );
na02f80 g542454 ( .a(n_25138), .b(FE_OFN290_n_27194), .o(n_26329) );
oa12f80 g542455 ( .a(n_26024), .b(FE_OFN40_n_25450), .c(n_25424), .o(n_26624) );
oa12f80 g542456 ( .a(n_26929), .b(n_1448), .c(FE_OFN360_n_4860), .o(n_26931) );
oa12f80 g542457 ( .a(n_26929), .b(n_1415), .c(FE_OFN75_n_27012), .o(n_26930) );
ao22s80 g542458 ( .a(n_24847), .b(FE_OFN606_n_25225), .c(x_out_50_30), .d(FE_OFN1162_n_5003), .o(n_25816) );
oa12f80 g542459 ( .a(n_25740), .b(n_25513), .c(n_24814), .o(n_26311) );
na02f80 g542460 ( .a(n_25514), .b(n_25137), .o(n_26633) );
oa12f80 g542461 ( .a(n_26606), .b(n_847), .c(FE_OFN360_n_4860), .o(n_26608) );
oa12f80 g542462 ( .a(n_26606), .b(n_1311), .c(FE_OFN360_n_4860), .o(n_26607) );
no02f80 g542463 ( .a(n_25814), .b(n_25813), .o(n_25815) );
no02f80 g542464 ( .a(n_25814), .b(n_25100), .o(n_27007) );
ao12f80 g542465 ( .a(n_15811), .b(n_24966), .c(n_16498), .o(n_25963) );
na02f80 g542466 ( .a(n_25425), .b(n_25451), .o(n_26023) );
ao12f80 g542467 ( .a(n_14403), .b(n_25269), .c(n_15174), .o(n_26217) );
in01f80 g542468 ( .a(n_28268), .o(n_28641) );
oa12f80 g542469 ( .a(n_27002), .b(n_28122), .c(n_26447), .o(n_28268) );
ao12f80 g542470 ( .a(n_15424), .b(n_25268), .c(n_16121), .o(n_26216) );
oa12f80 g542471 ( .a(n_15420), .b(n_25266), .c(n_15843), .o(n_25267) );
oa12f80 g542472 ( .a(n_14937), .b(n_24640), .c(n_15546), .o(n_25357) );
oa12f80 g542473 ( .a(n_15357), .b(n_24962), .c(n_15838), .o(n_24963) );
oa12f80 g542474 ( .a(n_15402), .b(n_24960), .c(n_15835), .o(n_24961) );
oa12f80 g542475 ( .a(n_15392), .b(n_24958), .c(n_15828), .o(n_24959) );
ao12f80 g542476 ( .a(n_12264), .b(n_24956), .c(n_12465), .o(n_25660) );
oa12f80 g542477 ( .a(n_15380), .b(n_24954), .c(n_15825), .o(n_24955) );
oa12f80 g542478 ( .a(n_15362), .b(n_24952), .c(n_15822), .o(n_24953) );
in01f80 g542479 ( .a(n_27740), .o(n_28228) );
oa12f80 g542480 ( .a(n_25981), .b(n_25722), .c(n_27563), .o(n_27740) );
in01f80 g542481 ( .a(n_28125), .o(n_28521) );
oa12f80 g542482 ( .a(n_26837), .b(n_26478), .c(n_28003), .o(n_28125) );
in01f80 g542483 ( .a(n_28008), .o(n_28407) );
oa12f80 g542484 ( .a(n_26833), .b(n_26476), .c(n_27875), .o(n_28008) );
ao12f80 g542485 ( .a(n_11797), .b(n_24947), .c(n_13114), .o(n_25688) );
in01f80 g542486 ( .a(n_28007), .o(n_28404) );
oa12f80 g542487 ( .a(n_25736), .b(n_25388), .c(n_27872), .o(n_28007) );
oa12f80 g542488 ( .a(FE_OFN44_n_25810), .b(n_1261), .c(FE_OFN91_n_27449), .o(n_25812) );
oa12f80 g542489 ( .a(FE_OFN44_n_25810), .b(n_552), .c(FE_OFN91_n_27449), .o(n_25811) );
oa12f80 g542490 ( .a(n_25142), .b(n_25143), .c(n_23829), .o(n_25809) );
oa12f80 g542491 ( .a(FE_OFN44_n_25810), .b(n_1678), .c(FE_OFN12_n_29204), .o(n_25808) );
oa12f80 g542492 ( .a(n_26021), .b(n_1589), .c(FE_OFN1123_rst), .o(n_26022) );
oa12f80 g542493 ( .a(n_25536), .b(n_487), .c(FE_OFN104_n_27449), .o(n_25537) );
oa12f80 g542494 ( .a(n_26309), .b(n_71), .c(FE_OFN108_n_27449), .o(n_26310) );
ao12f80 g542495 ( .a(n_16486), .b(n_24943), .c(n_16984), .o(n_25634) );
ao12f80 g542496 ( .a(n_15181), .b(n_25535), .c(n_15861), .o(n_26104) );
na03f80 g542497 ( .a(n_25819), .b(n_25820), .c(n_12352), .o(n_26020) );
ao12f80 g542498 ( .a(n_13139), .b(n_25263), .c(n_14295), .o(n_25264) );
oa12f80 g542499 ( .a(n_26262), .b(n_27739), .c(n_26214), .o(n_28234) );
oa12f80 g542500 ( .a(n_12266), .b(n_24942), .c(n_12942), .o(n_25966) );
ao12f80 g542501 ( .a(n_14884), .b(n_25806), .c(n_15137), .o(n_25807) );
oa12f80 g542502 ( .a(n_15763), .b(n_24941), .c(n_16490), .o(n_25629) );
oa12f80 g542503 ( .a(n_15831), .b(n_25262), .c(n_16487), .o(n_25871) );
oa12f80 g542504 ( .a(n_9450), .b(n_25531), .c(n_25530), .o(n_25534) );
in01f80 g542505 ( .a(n_24939), .o(n_25937) );
oa12f80 g542506 ( .a(n_11786), .b(n_24627), .c(n_13109), .o(n_24939) );
ao12f80 g542507 ( .a(n_13633), .b(n_25533), .c(n_14325), .o(n_26501) );
ao12f80 g542508 ( .a(n_15784), .b(n_24938), .c(n_16473), .o(n_25938) );
ao12f80 g542509 ( .a(n_15777), .b(n_24937), .c(n_16470), .o(n_25936) );
no02f80 g542510 ( .a(n_26618), .b(n_25944), .o(n_27197) );
ao12f80 g542511 ( .a(n_14923), .b(n_24936), .c(n_15493), .o(n_25964) );
ao12f80 g542512 ( .a(n_15768), .b(n_24935), .c(n_16469), .o(n_25935) );
oa12f80 g542513 ( .a(n_15806), .b(n_24934), .c(n_16483), .o(n_25605) );
ao12f80 g542514 ( .a(n_11779), .b(n_24931), .c(n_13108), .o(n_25602) );
ao12f80 g542515 ( .a(n_9331), .b(n_25531), .c(n_25530), .o(n_25532) );
in01f80 g542516 ( .a(n_25860), .o(n_26146) );
ao12f80 g542517 ( .a(n_24560), .b(n_24966), .c(n_24559), .o(n_25860) );
ao12f80 g542518 ( .a(n_25172), .b(n_25171), .c(n_25170), .o(n_25805) );
ao12f80 g542519 ( .a(n_27541), .b(n_27540), .c(n_27539), .o(n_27890) );
ao12f80 g542520 ( .a(n_27538), .b(n_27537), .c(n_27536), .o(n_27889) );
in01f80 g542521 ( .a(n_26019), .o(n_26670) );
ao12f80 g542522 ( .a(n_25186), .b(n_25535), .c(n_25185), .o(n_26019) );
oa12f80 g542523 ( .a(n_24870), .b(n_24869), .c(n_25169), .o(n_26144) );
in01f80 g542524 ( .a(n_25529), .o(n_26459) );
oa12f80 g542525 ( .a(n_24558), .b(n_24561), .c(n_24557), .o(n_25529) );
ao12f80 g542526 ( .a(n_27535), .b(n_27534), .c(n_27533), .o(n_27888) );
oa12f80 g542527 ( .a(n_25168), .b(n_25167), .c(n_25439), .o(n_26426) );
ao12f80 g542528 ( .a(n_25990), .b(n_25989), .c(n_25988), .o(n_26604) );
ao22s80 g542529 ( .a(n_27238), .b(n_27653), .c(n_27239), .d(n_28122), .o(n_28123) );
ao12f80 g542530 ( .a(n_27145), .b(n_27144), .c(n_27143), .o(n_27571) );
ao12f80 g542531 ( .a(n_27530), .b(n_27529), .c(n_27528), .o(n_27887) );
oa12f80 g542532 ( .a(n_25166), .b(n_25165), .c(n_25164), .o(n_26424) );
ao12f80 g542533 ( .a(n_26915), .b(n_26914), .c(n_26913), .o(n_27359) );
ao12f80 g542534 ( .a(n_27527), .b(n_27526), .c(n_27525), .o(n_27886) );
oa12f80 g542535 ( .a(n_25163), .b(n_25162), .c(n_25161), .o(n_26423) );
ao12f80 g542536 ( .a(n_25755), .b(n_25754), .c(n_25753), .o(n_26308) );
ao12f80 g542537 ( .a(n_27339), .b(n_27338), .c(n_27337), .o(n_27738) );
oa12f80 g542538 ( .a(n_24868), .b(n_24867), .c(n_25160), .o(n_26142) );
in01f80 g542539 ( .a(n_25804), .o(n_26420) );
ao12f80 g542540 ( .a(n_24899), .b(n_25268), .c(n_24898), .o(n_25804) );
ao12f80 g542541 ( .a(n_27336), .b(n_27335), .c(n_27334), .o(n_27735) );
oa12f80 g542542 ( .a(n_24866), .b(n_24865), .c(n_25159), .o(n_26140) );
ao12f80 g542543 ( .a(n_27333), .b(n_27332), .c(n_27331), .o(n_27734) );
oa12f80 g542544 ( .a(n_24864), .b(n_24863), .c(n_25158), .o(n_26139) );
in01f80 g542545 ( .a(n_26094), .o(n_26366) );
ao12f80 g542546 ( .a(n_24897), .b(n_25269), .c(n_24896), .o(n_26094) );
ao12f80 g542547 ( .a(n_27330), .b(n_27329), .c(n_27328), .o(n_27733) );
oa12f80 g542548 ( .a(n_25157), .b(n_25156), .c(n_25155), .o(n_26414) );
oa12f80 g542549 ( .a(n_25154), .b(n_25153), .c(n_25434), .o(n_26413) );
ao12f80 g542550 ( .a(n_26918), .b(n_26917), .c(n_26916), .o(n_27358) );
ao12f80 g542551 ( .a(n_27327), .b(n_27326), .c(n_27325), .o(n_27730) );
oa12f80 g542552 ( .a(n_25182), .b(n_25221), .c(n_25448), .o(n_26412) );
ao12f80 g542553 ( .a(n_27324), .b(n_27323), .c(n_27322), .o(n_27729) );
oa12f80 g542554 ( .a(n_24878), .b(n_24892), .c(n_25181), .o(n_26138) );
ao12f80 g542555 ( .a(n_27521), .b(n_27520), .c(n_27519), .o(n_27885) );
ao12f80 g542556 ( .a(n_27518), .b(n_27517), .c(n_27516), .o(n_27884) );
ao12f80 g542557 ( .a(n_27524), .b(n_27523), .c(n_27522), .o(n_27883) );
in01f80 g542558 ( .a(n_26544), .o(n_26408) );
ao12f80 g542559 ( .a(n_24895), .b(n_25266), .c(n_24894), .o(n_26544) );
ao12f80 g542560 ( .a(n_26912), .b(n_26911), .c(n_26910), .o(n_27357) );
in01f80 g542561 ( .a(n_26092), .o(n_26136) );
ao12f80 g542562 ( .a(n_24545), .b(n_24941), .c(n_24544), .o(n_26092) );
oa12f80 g542563 ( .a(n_24877), .b(n_24891), .c(n_25180), .o(n_26137) );
ao12f80 g542564 ( .a(n_27321), .b(n_27320), .c(n_27319), .o(n_27728) );
oa12f80 g542565 ( .a(n_24202), .b(n_24640), .c(n_24201), .o(n_25847) );
oa12f80 g542566 ( .a(n_24876), .b(n_24890), .c(n_25183), .o(n_26135) );
ao12f80 g542567 ( .a(n_27318), .b(n_27317), .c(n_27316), .o(n_27727) );
ao12f80 g542568 ( .a(n_27315), .b(n_27314), .c(n_27313), .o(n_27726) );
ao12f80 g542569 ( .a(n_27515), .b(n_27514), .c(n_27513), .o(n_27882) );
oa12f80 g542570 ( .a(n_24875), .b(n_24888), .c(n_25178), .o(n_26132) );
in01f80 g542571 ( .a(n_26253), .o(n_26131) );
ao12f80 g542572 ( .a(n_24698), .b(n_24962), .c(n_24697), .o(n_26253) );
ao12f80 g542573 ( .a(n_27617), .b(n_27616), .c(n_27739), .o(n_27881) );
ao12f80 g542574 ( .a(n_27312), .b(n_27311), .c(n_27310), .o(n_27725) );
ao12f80 g542575 ( .a(n_27142), .b(n_27141), .c(n_27140), .o(n_27569) );
in01f80 g542576 ( .a(n_26251), .o(n_26130) );
ao12f80 g542577 ( .a(n_24649), .b(n_24960), .c(n_24648), .o(n_26251) );
ao12f80 g542578 ( .a(n_27856), .b(n_27855), .c(n_27854), .o(n_28121) );
in01f80 g542579 ( .a(n_25846), .o(n_26069) );
ao12f80 g542580 ( .a(n_24547), .b(n_24942), .c(n_24546), .o(n_25846) );
in01f80 g542581 ( .a(n_26363), .o(n_26392) );
ao12f80 g542582 ( .a(n_24880), .b(n_25262), .c(n_24879), .o(n_26363) );
ao12f80 g542583 ( .a(n_27512), .b(n_27511), .c(n_27510), .o(n_27880) );
in01f80 g542584 ( .a(n_26249), .o(n_26129) );
ao12f80 g542585 ( .a(n_24564), .b(n_24958), .c(n_24563), .o(n_26249) );
ao12f80 g542586 ( .a(n_27309), .b(n_27308), .c(n_27307), .o(n_27724) );
in01f80 g542587 ( .a(n_25854), .o(n_26128) );
ao12f80 g542588 ( .a(n_24506), .b(n_24956), .c(n_24505), .o(n_25854) );
in01f80 g542589 ( .a(n_26637), .o(n_26307) );
ao12f80 g542590 ( .a(n_25453), .b(n_25806), .c(n_25452), .o(n_26637) );
ao12f80 g542591 ( .a(n_27509), .b(n_27508), .c(n_27507), .o(n_27879) );
in01f80 g542592 ( .a(n_26247), .o(n_26126) );
ao12f80 g542593 ( .a(n_24555), .b(n_24954), .c(n_24554), .o(n_26247) );
ao12f80 g542594 ( .a(n_27306), .b(n_27305), .c(n_27304), .o(n_27723) );
in01f80 g542595 ( .a(n_25864), .o(n_26125) );
ao12f80 g542596 ( .a(n_24549), .b(n_24943), .c(n_24548), .o(n_25864) );
ao12f80 g542597 ( .a(n_27506), .b(n_27505), .c(n_27504), .o(n_27878) );
in01f80 g542598 ( .a(n_26245), .o(n_26124) );
ao12f80 g542599 ( .a(n_24553), .b(n_24952), .c(n_24552), .o(n_26245) );
ao12f80 g542600 ( .a(n_27139), .b(n_27138), .c(n_27137), .o(n_27568) );
in01f80 g542601 ( .a(n_26694), .o(n_26381) );
oa12f80 g542602 ( .a(n_24885), .b(n_24884), .c(n_24883), .o(n_26694) );
oa12f80 g542603 ( .a(n_24862), .b(n_24861), .c(n_25152), .o(n_26123) );
ao12f80 g542604 ( .a(n_26593), .b(n_26592), .c(n_26591), .o(n_27156) );
ao12f80 g542605 ( .a(n_27136), .b(n_27135), .c(n_27134), .o(n_27567) );
oa12f80 g542606 ( .a(n_25151), .b(n_25150), .c(n_25149), .o(n_26378) );
oa12f80 g542607 ( .a(n_24874), .b(n_24889), .c(n_25179), .o(n_26133) );
ao12f80 g542608 ( .a(n_27502), .b(n_27501), .c(n_27500), .o(n_27877) );
in01f80 g542609 ( .a(n_25862), .o(n_26119) );
ao12f80 g542610 ( .a(n_24535), .b(n_24934), .c(n_24534), .o(n_25862) );
oa12f80 g542611 ( .a(n_25751), .b(n_25750), .c(n_25749), .o(n_26974) );
in01f80 g542612 ( .a(n_26351), .o(n_26643) );
ao12f80 g542613 ( .a(n_25176), .b(n_25533), .c(n_25175), .o(n_26351) );
ao12f80 g542614 ( .a(n_25148), .b(n_25147), .c(n_25146), .o(n_25803) );
ao22s80 g542615 ( .a(n_26265), .b(n_27563), .c(n_26264), .d(n_26830), .o(n_27564) );
ao22s80 g542616 ( .a(n_27070), .b(n_28003), .c(n_27069), .d(n_27459), .o(n_28004) );
in01f80 g542617 ( .a(n_26358), .o(n_26018) );
ao12f80 g542618 ( .a(n_25174), .b(n_25184), .c(n_25173), .o(n_26358) );
ao12f80 g542619 ( .a(n_27283), .b(n_27282), .c(FE_OFN492_n_28765), .o(n_29096) );
ao12f80 g542620 ( .a(n_26904), .b(n_26903), .c(n_26902), .o(n_27356) );
ao12f80 g542621 ( .a(n_27678), .b(n_27677), .c(n_27676), .o(n_28000) );
oa12f80 g542622 ( .a(n_25432), .b(n_25431), .c(n_25430), .o(n_26644) );
in01f80 g542623 ( .a(n_26075), .o(n_26409) );
ao12f80 g542624 ( .a(n_24882), .b(n_25263), .c(n_24881), .o(n_26075) );
oa12f80 g542625 ( .a(n_24539), .b(n_24936), .c(n_24538), .o(n_26078) );
ao12f80 g542626 ( .a(n_26900), .b(n_26899), .c(n_26898), .o(n_27355) );
oa22f80 g542627 ( .a(n_24196), .b(n_24195), .c(n_5782), .d(n_8453), .o(n_24594) );
ao22s80 g542628 ( .a(n_27066), .b(n_27875), .c(n_27065), .d(n_27259), .o(n_27876) );
oa12f80 g542629 ( .a(n_26601), .b(n_26602), .c(x_in_56_15), .o(n_29315) );
ao12f80 g542630 ( .a(n_27498), .b(n_27497), .c(n_27496), .o(n_27874) );
ao12f80 g542631 ( .a(n_24858), .b(n_24857), .c(n_24856), .o(n_25528) );
in01f80 g542632 ( .a(n_26087), .o(n_26116) );
ao12f80 g542633 ( .a(n_24543), .b(n_24938), .c(n_24542), .o(n_26087) );
in01f80 g542634 ( .a(n_25848), .o(n_26073) );
ao12f80 g542635 ( .a(n_24551), .b(n_24947), .c(n_24550), .o(n_25848) );
ao22s80 g542636 ( .a(n_25979), .b(n_27872), .c(n_25978), .d(n_27258), .o(n_27873) );
ao12f80 g542637 ( .a(n_24873), .b(n_25253), .c(n_24872), .o(n_25527) );
in01f80 g542638 ( .a(n_25600), .o(n_25868) );
ao12f80 g542639 ( .a(n_24199), .b(n_24627), .c(n_24198), .o(n_25600) );
in01f80 g542640 ( .a(n_26629), .o(n_26969) );
oa12f80 g542641 ( .a(n_25464), .b(n_25463), .c(n_25462), .o(n_26629) );
ao12f80 g542642 ( .a(n_27493), .b(n_27492), .c(n_27491), .o(n_27871) );
in01f80 g542643 ( .a(n_26084), .o(n_26115) );
ao12f80 g542644 ( .a(n_24541), .b(n_24937), .c(n_24540), .o(n_26084) );
oa12f80 g542645 ( .a(n_25748), .b(n_25747), .c(n_25985), .o(n_26968) );
oa12f80 g542647 ( .a(n_25461), .b(n_25460), .c(n_25459), .o(n_32744) );
ao12f80 g542648 ( .a(n_25195), .b(n_25194), .c(n_25193), .o(n_25802) );
in01f80 g542649 ( .a(n_25526), .o(n_26443) );
oa12f80 g542650 ( .a(n_24533), .b(n_24931), .c(n_24532), .o(n_25526) );
ao12f80 g542651 ( .a(n_27300), .b(n_27299), .c(n_27298), .o(n_27722) );
oa12f80 g542652 ( .a(n_25984), .b(n_25983), .c(n_25982), .o(n_27198) );
ao12f80 g542653 ( .a(n_27544), .b(n_27543), .c(n_27542), .o(n_27870) );
ao12f80 g542654 ( .a(n_25192), .b(n_25191), .c(n_25190), .o(n_25801) );
ao12f80 g542655 ( .a(n_27490), .b(n_27489), .c(n_27488), .o(n_27869) );
ao12f80 g542656 ( .a(n_27674), .b(n_27673), .c(n_27672), .o(n_27999) );
oa12f80 g542657 ( .a(n_24530), .b(n_24529), .c(n_24855), .o(n_25873) );
in01f80 g542658 ( .a(n_26081), .o(n_26106) );
ao12f80 g542659 ( .a(n_24537), .b(n_24935), .c(n_24536), .o(n_26081) );
ao12f80 g542660 ( .a(n_24854), .b(n_24853), .c(n_24852), .o(n_25525) );
ao12f80 g542661 ( .a(n_26286), .b(n_26285), .c(n_26284), .o(n_26925) );
ao12f80 g542662 ( .a(n_26894), .b(n_26893), .c(n_26892), .o(n_27354) );
oa12f80 g542663 ( .a(n_25177), .b(n_25201), .c(n_25443), .o(n_26369) );
ao12f80 g542664 ( .a(n_27293), .b(n_27292), .c(n_27291), .o(n_27721) );
ao22s80 g542665 ( .a(n_26016), .b(n_25442), .c(x_out_46_31), .d(FE_OFN1162_n_5003), .o(n_26017) );
oa12f80 g542666 ( .a(n_25429), .b(n_25428), .c(n_25746), .o(n_26639) );
oa22f80 g542667 ( .a(n_25098), .b(FE_OFN314_n_3069), .c(n_1199), .d(FE_OFN119_n_27449), .o(n_26014) );
oa22f80 g542668 ( .a(n_27062), .b(FE_OFN156_n_28014), .c(n_831), .d(FE_OFN330_n_4860), .o(n_27720) );
oa22f80 g542669 ( .a(n_24886), .b(FE_OFN157_n_28014), .c(n_1382), .d(FE_OFN128_n_27449), .o(n_25255) );
oa22f80 g542670 ( .a(n_27061), .b(FE_OFN402_n_28303), .c(n_413), .d(FE_OFN69_n_27012), .o(n_27719) );
oa22f80 g542671 ( .a(FE_OFN744_n_25732), .b(n_22960), .c(n_1968), .d(n_29204), .o(n_26603) );
oa22f80 g542672 ( .a(n_27257), .b(FE_OFN402_n_28303), .c(n_570), .d(FE_OFN11_n_29204), .o(n_27866) );
oa22f80 g542673 ( .a(n_27060), .b(FE_OFN417_n_28303), .c(n_1367), .d(FE_OFN361_n_4860), .o(n_27716) );
oa22f80 g542674 ( .a(n_27455), .b(FE_OFN234_n_4162), .c(n_957), .d(FE_OFN76_n_27012), .o(n_27998) );
oa22f80 g542675 ( .a(n_25097), .b(FE_OFN311_n_3069), .c(n_1650), .d(FE_OFN134_n_27449), .o(n_26013) );
oa22f80 g542676 ( .a(n_27059), .b(FE_OFN244_n_4162), .c(n_239), .d(FE_OFN131_n_27449), .o(n_27713) );
oa22f80 g542677 ( .a(n_24831), .b(n_4162), .c(n_136), .d(FE_OFN116_n_27449), .o(n_25800) );
oa22f80 g542678 ( .a(n_27058), .b(FE_OFN248_n_4162), .c(n_1376), .d(FE_OFN90_n_27449), .o(n_27711) );
oa22f80 g542679 ( .a(n_26829), .b(FE_OFN239_n_4162), .c(n_600), .d(FE_OFN135_n_27449), .o(n_27561) );
oa22f80 g542680 ( .a(n_26828), .b(FE_OFN308_n_3069), .c(n_837), .d(FE_OFN90_n_27449), .o(n_27560) );
oa22f80 g542681 ( .a(n_24830), .b(FE_OFN314_n_3069), .c(n_1717), .d(FE_OFN119_n_27449), .o(n_25799) );
oa22f80 g542682 ( .a(n_26548), .b(FE_OFN400_n_28303), .c(n_1232), .d(n_29264), .o(n_27353) );
oa22f80 g542683 ( .a(n_26827), .b(FE_OFN257_n_4280), .c(n_1139), .d(n_27709), .o(n_27559) );
oa22f80 g542684 ( .a(FE_OFN1047_n_27057), .b(FE_OFN400_n_28303), .c(n_1534), .d(n_27709), .o(n_27710) );
oa22f80 g542685 ( .a(n_27056), .b(FE_OFN247_n_4162), .c(n_250), .d(FE_OFN128_n_27449), .o(n_27708) );
oa22f80 g542686 ( .a(n_26826), .b(FE_OFN248_n_4162), .c(n_771), .d(FE_OFN113_n_27449), .o(n_27557) );
oa22f80 g542687 ( .a(n_26547), .b(FE_OFN230_n_4162), .c(n_307), .d(FE_OFN1108_rst), .o(n_27352) );
oa22f80 g542688 ( .a(n_27055), .b(FE_OFN404_n_28303), .c(n_1727), .d(FE_OFN350_n_4860), .o(n_27704) );
oa22f80 g542689 ( .a(n_26825), .b(FE_OFN240_n_4162), .c(n_537), .d(FE_OFN17_n_29617), .o(n_27556) );
oa22f80 g542690 ( .a(n_26824), .b(FE_OFN230_n_4162), .c(n_1936), .d(n_29617), .o(n_27554) );
oa22f80 g542691 ( .a(n_27040), .b(FE_OFN249_n_4162), .c(n_5), .d(FE_OFN98_n_27449), .o(n_27702) );
oa22f80 g542692 ( .a(n_26259), .b(FE_OFN211_n_29661), .c(n_1069), .d(FE_OFN355_n_4860), .o(n_27155) );
oa22f80 g542693 ( .a(n_27053), .b(FE_OFN208_n_29661), .c(n_1055), .d(FE_OFN101_n_27449), .o(n_27701) );
oa22f80 g542694 ( .a(n_26823), .b(FE_OFN405_n_28303), .c(n_1316), .d(FE_OFN94_n_27449), .o(n_27553) );
oa22f80 g542695 ( .a(n_26822), .b(FE_OFN411_n_28303), .c(n_370), .d(FE_OFN335_n_4860), .o(n_27552) );
oa22f80 g542696 ( .a(n_26821), .b(FE_OFN405_n_28303), .c(n_381), .d(FE_OFN357_n_4860), .o(n_27551) );
oa22f80 g542697 ( .a(n_27047), .b(FE_OFN4_n_28682), .c(n_16), .d(FE_OFN115_n_27449), .o(n_27700) );
oa22f80 g542698 ( .a(n_24499), .b(FE_OFN4_n_28682), .c(n_960), .d(FE_OFN115_n_27449), .o(n_25524) );
oa22f80 g542699 ( .a(FE_OFN558_n_26546), .b(n_29698), .c(n_281), .d(n_27449), .o(n_27351) );
oa22f80 g542700 ( .a(n_25253), .b(FE_OFN400_n_28303), .c(n_396), .d(FE_OFN20_n_27452), .o(n_25254) );
oa22f80 g542701 ( .a(n_27446), .b(FE_OFN417_n_28303), .c(n_447), .d(n_28928), .o(n_27989) );
oa22f80 g542702 ( .a(n_24887), .b(FE_OFN410_n_28303), .c(n_1048), .d(FE_OFN100_n_27449), .o(n_25249) );
oa22f80 g542703 ( .a(n_26820), .b(n_29691), .c(n_38), .d(FE_OFN101_n_27449), .o(n_27550) );
oa22f80 g542704 ( .a(n_27043), .b(FE_OFN405_n_28303), .c(n_1708), .d(n_27449), .o(n_27699) );
oa22f80 g542705 ( .a(n_24507), .b(FE_OFN299_n_3069), .c(n_1212), .d(FE_OFN74_n_27012), .o(n_25523) );
oa22f80 g542706 ( .a(n_26819), .b(FE_OFN413_n_28303), .c(n_88), .d(FE_OFN133_n_27449), .o(n_27549) );
oa22f80 g542707 ( .a(n_26254), .b(FE_OFN259_n_4280), .c(n_1644), .d(FE_OFN1120_rst), .o(n_27153) );
oa22f80 g542708 ( .a(n_26545), .b(FE_OFN414_n_28303), .c(n_1317), .d(FE_OFN1113_rst), .o(n_27350) );
oa22f80 g542709 ( .a(n_25758), .b(FE_OFN254_n_4280), .c(n_776), .d(FE_OFN361_n_4860), .o(n_26012) );
oa22f80 g542710 ( .a(n_26818), .b(FE_OFN254_n_4280), .c(n_1244), .d(FE_OFN361_n_4860), .o(n_27548) );
oa22f80 g542711 ( .a(n_27042), .b(FE_OFN411_n_28303), .c(n_1947), .d(FE_OFN114_n_27449), .o(n_27698) );
oa22f80 g542712 ( .a(n_27041), .b(n_28303), .c(n_1854), .d(FE_OFN357_n_4860), .o(n_27696) );
oa22f80 g542713 ( .a(n_27039), .b(FE_OFN4_n_28682), .c(n_1764), .d(FE_OFN335_n_4860), .o(n_27695) );
oa22f80 g542714 ( .a(n_24501), .b(FE_OFN3_n_28682), .c(n_860), .d(FE_OFN358_n_4860), .o(n_25522) );
oa22f80 g542715 ( .a(n_26243), .b(n_29496), .c(n_1869), .d(FE_OFN142_n_27449), .o(n_27152) );
oa22f80 g542716 ( .a(n_26542), .b(FE_OFN212_n_29661), .c(n_507), .d(FE_OFN133_n_27449), .o(n_27349) );
oa22f80 g542717 ( .a(n_24500), .b(FE_OFN212_n_29661), .c(n_52), .d(FE_OFN138_n_27449), .o(n_25520) );
oa22f80 g542718 ( .a(n_26541), .b(FE_OFN240_n_4162), .c(n_1106), .d(FE_OFN141_n_27449), .o(n_27348) );
oa22f80 g542719 ( .a(FE_OFN488_n_27256), .b(n_29691), .c(n_409), .d(FE_OFN101_n_27449), .o(n_27859) );
oa22f80 g542720 ( .a(n_25438), .b(n_4162), .c(n_1797), .d(FE_OFN116_n_27449), .o(n_25797) );
oa22f80 g542721 ( .a(n_26242), .b(FE_OFN249_n_4162), .c(n_1842), .d(FE_OFN64_n_27012), .o(n_27150) );
oa22f80 g542722 ( .a(n_26241), .b(FE_OFN244_n_4162), .c(n_979), .d(FE_OFN77_n_27012), .o(n_27149) );
oa22f80 g542723 ( .a(n_27038), .b(FE_OFN259_n_4280), .c(n_540), .d(FE_OFN350_n_4860), .o(n_27691) );
oa22f80 g542724 ( .a(n_27037), .b(n_4162), .c(n_328), .d(FE_OFN115_n_27449), .o(n_27690) );
oa22f80 g542725 ( .a(n_24826), .b(FE_OFN180_n_27681), .c(n_859), .d(FE_OFN134_n_27449), .o(n_25796) );
oa22f80 g542726 ( .a(n_24859), .b(FE_OFN181_n_27681), .c(n_1604), .d(FE_OFN141_n_27449), .o(n_25233) );
oa22f80 g542727 ( .a(n_27032), .b(FE_OFN308_n_3069), .c(n_1963), .d(FE_OFN90_n_27449), .o(n_27686) );
oa22f80 g542728 ( .a(n_27034), .b(FE_OFN297_n_3069), .c(n_1118), .d(FE_OFN141_n_27449), .o(n_27685) );
oa22f80 g542729 ( .a(n_25975), .b(FE_OFN308_n_3069), .c(n_746), .d(FE_OFN90_n_27449), .o(n_26924) );
oa22f80 g542730 ( .a(n_24498), .b(FE_OFN235_n_4162), .c(n_1602), .d(n_27449), .o(n_25518) );
oa22f80 g542731 ( .a(n_27031), .b(n_29687), .c(n_1579), .d(FE_OFN1109_rst), .o(n_27684) );
oa22f80 g542732 ( .a(n_24825), .b(FE_OFN234_n_4162), .c(n_619), .d(FE_OFN100_n_27449), .o(n_25795) );
oa22f80 g542733 ( .a(n_27030), .b(n_27681), .c(n_1610), .d(FE_OFN105_n_27449), .o(n_27682) );
oa22f80 g542734 ( .a(n_24824), .b(FE_OFN180_n_27681), .c(n_849), .d(FE_OFN128_n_27449), .o(n_25794) );
oa22f80 g542735 ( .a(n_27253), .b(FE_OFN247_n_4162), .c(n_1763), .d(FE_OFN134_n_27449), .o(n_27858) );
oa22f80 g542736 ( .a(n_24823), .b(FE_OFN239_n_4162), .c(n_78), .d(FE_OFN135_n_27449), .o(n_25793) );
oa22f80 g542737 ( .a(n_25974), .b(FE_OFN259_n_4280), .c(n_298), .d(FE_OFN74_n_27012), .o(n_26923) );
oa22f80 g542738 ( .a(n_26815), .b(FE_OFN267_n_4280), .c(n_753), .d(FE_OFN91_n_27449), .o(n_27546) );
oa22f80 g542739 ( .a(n_26240), .b(FE_OFN4_n_28682), .c(n_270), .d(FE_OFN134_n_27449), .o(n_27147) );
oa22f80 g542740 ( .a(n_26239), .b(n_28682), .c(n_1217), .d(FE_OFN124_n_27449), .o(n_27146) );
oa22f80 g542741 ( .a(n_25404), .b(FE_OFN416_n_28303), .c(n_229), .d(FE_OFN134_n_27449), .o(n_26306) );
ao22s80 g542742 ( .a(n_25516), .b(n_24531), .c(x_out_33_30), .d(n_16028), .o(n_25517) );
ao22s80 g542743 ( .a(n_24182), .b(n_5398), .c(n_11854), .d(n_11853), .o(n_25228) );
na02f80 g542827 ( .a(n_25513), .b(n_25089), .o(n_25514) );
no02f80 g542828 ( .a(n_25408), .b(n_25407), .o(n_26618) );
in01f80 g542829 ( .a(n_26921), .o(n_26922) );
no02f80 g542830 ( .a(n_26602), .b(x_in_56_13), .o(n_26921) );
na02f80 g542831 ( .a(n_26602), .b(x_in_56_13), .o(n_27364) );
in01f80 g542832 ( .a(n_26919), .o(n_26920) );
no02f80 g542833 ( .a(n_26602), .b(x_in_56_14), .o(n_26919) );
na02f80 g542834 ( .a(n_26602), .b(x_in_56_14), .o(n_27363) );
na02f80 g542835 ( .a(n_26602), .b(x_in_56_15), .o(n_26601) );
no02f80 g542836 ( .a(n_24561), .b(n_12665), .o(n_24562) );
in01f80 g542837 ( .a(n_25511), .o(n_25512) );
no02f80 g542838 ( .a(n_25187), .b(x_in_58_12), .o(n_25511) );
no02f80 g542839 ( .a(n_27543), .b(n_27542), .o(n_27544) );
na02f80 g542840 ( .a(n_25792), .b(x_in_60_11), .o(n_26616) );
no02f80 g542841 ( .a(n_24966), .b(n_24559), .o(n_24560) );
no02f80 g542842 ( .a(n_27540), .b(n_27539), .o(n_27541) );
in01f80 g542843 ( .a(n_26010), .o(n_26011) );
no02f80 g542844 ( .a(n_25792), .b(x_in_60_11), .o(n_26010) );
no02f80 g542845 ( .a(n_27537), .b(n_27536), .o(n_27538) );
na02f80 g542846 ( .a(n_25510), .b(x_in_2_11), .o(n_26326) );
in01f80 g542847 ( .a(n_25790), .o(n_25791) );
no02f80 g542848 ( .a(n_25510), .b(x_in_2_11), .o(n_25790) );
na02f80 g542849 ( .a(n_24561), .b(n_24557), .o(n_24558) );
no02f80 g542850 ( .a(n_27534), .b(n_27533), .o(n_27535) );
na02f80 g542851 ( .a(n_25789), .b(x_in_34_11), .o(n_26615) );
in01f80 g542852 ( .a(n_26008), .o(n_26009) );
no02f80 g542853 ( .a(n_25789), .b(x_in_34_11), .o(n_26008) );
in01f80 g542854 ( .a(n_27531), .o(n_27532) );
na02f80 g542855 ( .a(n_27340), .b(n_26842), .o(n_27531) );
no02f80 g542856 ( .a(n_27529), .b(n_27528), .o(n_27530) );
na02f80 g542857 ( .a(n_25227), .b(x_in_18_11), .o(n_26049) );
in01f80 g542858 ( .a(n_25508), .o(n_25509) );
no02f80 g542859 ( .a(n_25227), .b(x_in_18_11), .o(n_25508) );
na02f80 g542860 ( .a(FE_OFN606_n_25225), .b(n_24846), .o(n_25226) );
no02f80 g542861 ( .a(n_27526), .b(n_27525), .o(n_27527) );
na02f80 g542862 ( .a(n_25224), .b(x_in_50_11), .o(n_26048) );
in01f80 g542863 ( .a(n_25506), .o(n_25507) );
no02f80 g542864 ( .a(n_25224), .b(x_in_50_11), .o(n_25506) );
no02f80 g542865 ( .a(n_27144), .b(n_27143), .o(n_27145) );
na02f80 g542866 ( .a(n_25504), .b(x_in_6_11), .o(n_26325) );
no02f80 g542867 ( .a(n_27338), .b(n_27337), .o(n_27339) );
na02f80 g542868 ( .a(n_25505), .b(x_in_10_11), .o(n_26324) );
in01f80 g542869 ( .a(n_25787), .o(n_25788) );
no02f80 g542870 ( .a(n_25505), .b(x_in_10_11), .o(n_25787) );
in01f80 g542871 ( .a(n_25785), .o(n_25786) );
no02f80 g542872 ( .a(n_25504), .b(x_in_6_11), .o(n_25785) );
no02f80 g542873 ( .a(n_25268), .b(n_24898), .o(n_24899) );
no02f80 g542874 ( .a(n_27335), .b(n_27334), .o(n_27336) );
na02f80 g542875 ( .a(n_25503), .b(x_in_42_11), .o(n_26323) );
in01f80 g542876 ( .a(n_25783), .o(n_25784) );
no02f80 g542877 ( .a(n_25503), .b(x_in_42_11), .o(n_25783) );
no02f80 g542878 ( .a(n_27332), .b(n_27331), .o(n_27333) );
na02f80 g542879 ( .a(n_25502), .b(x_in_26_11), .o(n_26322) );
in01f80 g542880 ( .a(n_25781), .o(n_25782) );
no02f80 g542881 ( .a(n_25502), .b(x_in_26_11), .o(n_25781) );
no02f80 g542882 ( .a(n_25269), .b(n_24896), .o(n_24897) );
no02f80 g542883 ( .a(n_27329), .b(n_27328), .o(n_27330) );
na02f80 g542884 ( .a(n_25223), .b(x_in_58_11), .o(n_26047) );
in01f80 g542885 ( .a(n_25500), .o(n_25501) );
no02f80 g542886 ( .a(n_25223), .b(x_in_58_11), .o(n_25500) );
na02f80 g542887 ( .a(n_25780), .b(x_in_6_10), .o(n_26614) );
in01f80 g542888 ( .a(n_26006), .o(n_26007) );
no02f80 g542889 ( .a(n_25780), .b(x_in_6_10), .o(n_26006) );
in01f80 g542890 ( .a(n_25778), .o(n_25779) );
na02f80 g542891 ( .a(n_25499), .b(n_24845), .o(n_25778) );
no02f80 g542892 ( .a(n_26917), .b(n_26916), .o(n_26918) );
in01f80 g542893 ( .a(n_26004), .o(n_26005) );
na02f80 g542894 ( .a(n_25777), .b(n_25129), .o(n_26004) );
no02f80 g542895 ( .a(n_27326), .b(n_27325), .o(n_27327) );
na02f80 g542896 ( .a(n_25498), .b(x_in_22_11), .o(n_26321) );
in01f80 g542897 ( .a(n_25775), .o(n_25776) );
no02f80 g542898 ( .a(n_25498), .b(x_in_22_11), .o(n_25775) );
no02f80 g542899 ( .a(n_27323), .b(n_27322), .o(n_27324) );
na02f80 g542900 ( .a(n_25222), .b(x_in_54_11), .o(n_26044) );
in01f80 g542901 ( .a(n_25496), .o(n_25497) );
no02f80 g542902 ( .a(n_25222), .b(x_in_54_11), .o(n_25496) );
no02f80 g542903 ( .a(n_27523), .b(n_27522), .o(n_27524) );
na02f80 g542904 ( .a(n_25495), .b(x_in_40_11), .o(n_26320) );
in01f80 g542905 ( .a(n_25773), .o(n_25774) );
no02f80 g542906 ( .a(n_25495), .b(x_in_40_11), .o(n_25773) );
no02f80 g542907 ( .a(n_27520), .b(n_27519), .o(n_27521) );
no02f80 g542908 ( .a(n_27517), .b(n_27516), .o(n_27518) );
na02f80 g542909 ( .a(n_25221), .b(x_in_22_12), .o(n_26042) );
na02f80 g542910 ( .a(n_25220), .b(x_in_2_12), .o(n_26043) );
no02f80 g542911 ( .a(n_26914), .b(n_26913), .o(n_26915) );
in01f80 g542912 ( .a(n_25493), .o(n_25494) );
no02f80 g542913 ( .a(n_25221), .b(x_in_22_12), .o(n_25493) );
in01f80 g542914 ( .a(n_25491), .o(n_25492) );
no02f80 g542915 ( .a(n_25220), .b(x_in_2_12), .o(n_25491) );
no02f80 g542916 ( .a(n_25266), .b(n_24894), .o(n_24895) );
na02f80 g542917 ( .a(n_24893), .b(x_in_52_11), .o(n_25829) );
no02f80 g542918 ( .a(n_26911), .b(n_26910), .o(n_26912) );
na02f80 g542919 ( .a(n_25219), .b(x_in_14_11), .o(n_26041) );
in01f80 g542920 ( .a(n_25489), .o(n_25490) );
no02f80 g542921 ( .a(n_25219), .b(x_in_14_11), .o(n_25489) );
in01f80 g542922 ( .a(n_25217), .o(n_25218) );
no02f80 g542923 ( .a(n_24893), .b(x_in_52_11), .o(n_25217) );
no02f80 g542924 ( .a(n_27320), .b(n_27319), .o(n_27321) );
na02f80 g542925 ( .a(n_25216), .b(x_in_46_11), .o(n_26040) );
in01f80 g542926 ( .a(n_25487), .o(n_25488) );
no02f80 g542927 ( .a(n_25216), .b(x_in_46_11), .o(n_25487) );
na02f80 g542928 ( .a(n_24640), .b(n_24201), .o(n_24202) );
no02f80 g542929 ( .a(n_27317), .b(n_27316), .o(n_27318) );
na02f80 g542930 ( .a(n_25215), .b(x_in_30_11), .o(n_26030) );
in01f80 g542931 ( .a(n_25485), .o(n_25486) );
no02f80 g542932 ( .a(n_25215), .b(x_in_30_11), .o(n_25485) );
no02f80 g542933 ( .a(n_27314), .b(n_27313), .o(n_27315) );
na02f80 g542934 ( .a(n_25214), .b(x_in_62_11), .o(n_26039) );
in01f80 g542935 ( .a(n_25483), .o(n_25484) );
no02f80 g542936 ( .a(n_25214), .b(x_in_62_11), .o(n_25483) );
no02f80 g542937 ( .a(n_27514), .b(n_27513), .o(n_27515) );
na02f80 g542938 ( .a(n_24892), .b(x_in_54_12), .o(n_25828) );
in01f80 g542939 ( .a(n_25212), .o(n_25213) );
no02f80 g542940 ( .a(n_24892), .b(x_in_54_12), .o(n_25212) );
no02f80 g542941 ( .a(n_24962), .b(n_24697), .o(n_24698) );
no02f80 g542942 ( .a(n_27616), .b(n_27739), .o(n_27617) );
no02f80 g542943 ( .a(n_27311), .b(n_27310), .o(n_27312) );
in01f80 g542944 ( .a(n_26303), .o(n_26304) );
no02f80 g542945 ( .a(n_26003), .b(x_in_36_11), .o(n_26303) );
no02f80 g542946 ( .a(n_27141), .b(n_27140), .o(n_27142) );
na02f80 g542947 ( .a(n_24891), .b(x_in_14_12), .o(n_25827) );
in01f80 g542948 ( .a(n_25210), .o(n_25211) );
no02f80 g542949 ( .a(n_24891), .b(x_in_14_12), .o(n_25210) );
no02f80 g542950 ( .a(n_24960), .b(n_24648), .o(n_24649) );
no02f80 g542951 ( .a(n_27855), .b(n_27854), .o(n_27856) );
na02f80 g542952 ( .a(n_25440), .b(x_in_34_12), .o(n_26318) );
in01f80 g542953 ( .a(n_25771), .o(n_25772) );
no02f80 g542954 ( .a(n_25440), .b(x_in_34_12), .o(n_25771) );
no02f80 g542955 ( .a(n_27511), .b(n_27510), .o(n_27512) );
na02f80 g542956 ( .a(n_24890), .b(x_in_46_12), .o(n_25826) );
in01f80 g542957 ( .a(n_25208), .o(n_25209) );
no02f80 g542958 ( .a(n_24890), .b(x_in_46_12), .o(n_25208) );
no02f80 g542959 ( .a(n_24958), .b(n_24563), .o(n_24564) );
no02f80 g542960 ( .a(n_27308), .b(n_27307), .o(n_27309) );
na02f80 g542961 ( .a(n_25207), .b(x_in_16_12), .o(n_26038) );
in01f80 g542962 ( .a(n_25481), .o(n_25482) );
no02f80 g542963 ( .a(n_25207), .b(x_in_16_12), .o(n_25481) );
no02f80 g542964 ( .a(n_24956), .b(n_24505), .o(n_24506) );
no02f80 g542965 ( .a(n_27508), .b(n_27507), .o(n_27509) );
na02f80 g542966 ( .a(n_24889), .b(x_in_30_12), .o(n_25825) );
in01f80 g542967 ( .a(n_25205), .o(n_25206) );
no02f80 g542968 ( .a(n_24889), .b(x_in_30_12), .o(n_25205) );
no02f80 g542969 ( .a(n_24954), .b(n_24554), .o(n_24555) );
no02f80 g542970 ( .a(n_27305), .b(n_27304), .o(n_27306) );
na02f80 g542971 ( .a(n_25204), .b(x_in_18_12), .o(n_26037) );
in01f80 g542972 ( .a(n_25479), .o(n_25480) );
no02f80 g542973 ( .a(n_25204), .b(x_in_18_12), .o(n_25479) );
no02f80 g542974 ( .a(n_27505), .b(n_27504), .o(n_27506) );
na02f80 g542975 ( .a(n_24888), .b(x_in_62_12), .o(n_25824) );
in01f80 g542976 ( .a(n_25202), .o(n_25203) );
no02f80 g542977 ( .a(n_24888), .b(x_in_62_12), .o(n_25202) );
no02f80 g542978 ( .a(n_24952), .b(n_24552), .o(n_24553) );
no02f80 g542979 ( .a(n_27138), .b(n_27137), .o(n_27139) );
na02f80 g542980 ( .a(n_25201), .b(x_in_12_12), .o(n_26036) );
in01f80 g542981 ( .a(n_25477), .o(n_25478) );
no02f80 g542982 ( .a(n_25201), .b(x_in_12_12), .o(n_25477) );
na02f80 g542983 ( .a(n_25476), .b(x_in_32_10), .o(n_26317) );
in01f80 g542984 ( .a(n_25769), .o(n_25770) );
no02f80 g542985 ( .a(n_25476), .b(x_in_32_10), .o(n_25769) );
no02f80 g542986 ( .a(n_26592), .b(n_26591), .o(n_26593) );
no02f80 g542987 ( .a(n_27135), .b(n_27134), .o(n_27136) );
na02f80 g542988 ( .a(n_25200), .b(x_in_16_11), .o(n_26035) );
in01f80 g542989 ( .a(n_25474), .o(n_25475) );
no02f80 g542990 ( .a(n_25200), .b(x_in_16_11), .o(n_25474) );
na02f80 g542991 ( .a(n_26003), .b(x_in_36_11), .o(n_26940) );
no02f80 g542992 ( .a(n_27501), .b(n_27500), .o(n_27502) );
na02f80 g542993 ( .a(n_25199), .b(x_in_50_12), .o(n_26034) );
in01f80 g542994 ( .a(n_25472), .o(n_25473) );
no02f80 g542995 ( .a(n_25199), .b(x_in_50_12), .o(n_25472) );
na02f80 g542996 ( .a(n_25768), .b(x_in_48_10), .o(n_26613) );
in01f80 g542997 ( .a(n_26001), .o(n_26002) );
no02f80 g542998 ( .a(n_25768), .b(x_in_48_10), .o(n_26001) );
in01f80 g542999 ( .a(n_27679), .o(n_27680) );
na02f80 g543000 ( .a(n_27499), .b(n_27068), .o(n_27679) );
na02f80 g543001 ( .a(n_25471), .b(x_in_40_10), .o(n_26316) );
in01f80 g543002 ( .a(n_25766), .o(n_25767) );
no02f80 g543003 ( .a(n_25471), .b(x_in_40_10), .o(n_25766) );
no02f80 g543004 ( .a(n_26903), .b(n_26902), .o(n_26904) );
na02f80 g543005 ( .a(n_25198), .b(x_in_32_11), .o(n_26033) );
in01f80 g543006 ( .a(n_25469), .o(n_25470) );
no02f80 g543007 ( .a(n_25198), .b(x_in_32_11), .o(n_25469) );
no02f80 g543008 ( .a(n_26899), .b(n_26898), .o(n_26900) );
na02f80 g543009 ( .a(n_26897), .b(x_in_56_12), .o(n_27578) );
in01f80 g543010 ( .a(n_27130), .o(n_27131) );
no02f80 g543011 ( .a(n_26897), .b(x_in_56_12), .o(n_27130) );
no02f80 g543012 ( .a(n_27497), .b(n_27496), .o(n_27498) );
na02f80 g543013 ( .a(n_25197), .b(x_in_10_12), .o(n_26032) );
in01f80 g543014 ( .a(n_25467), .o(n_25468) );
no02f80 g543015 ( .a(n_25197), .b(x_in_10_12), .o(n_25467) );
no02f80 g543016 ( .a(n_24947), .b(n_24550), .o(n_24551) );
in01f80 g543017 ( .a(n_25999), .o(n_26000) );
no02f80 g543018 ( .a(n_25765), .b(x_in_48_11), .o(n_25999) );
na02f80 g543019 ( .a(n_25765), .b(x_in_48_11), .o(n_26612) );
no02f80 g543020 ( .a(n_27677), .b(n_27676), .o(n_27678) );
na02f80 g543021 ( .a(n_25996), .b(x_in_20_11), .o(n_26935) );
in01f80 g543022 ( .a(n_25997), .o(n_25998) );
na02f80 g543023 ( .a(n_25764), .b(n_25111), .o(n_25997) );
in01f80 g543024 ( .a(n_26291), .o(n_26292) );
no02f80 g543025 ( .a(n_25996), .b(x_in_20_11), .o(n_26291) );
no02f80 g543026 ( .a(n_27492), .b(n_27491), .o(n_27493) );
na02f80 g543027 ( .a(n_25196), .b(x_in_42_12), .o(n_26031) );
in01f80 g543028 ( .a(n_25465), .o(n_25466) );
no02f80 g543029 ( .a(n_25196), .b(x_in_42_12), .o(n_25465) );
na02f80 g543030 ( .a(n_25463), .b(n_25462), .o(n_25464) );
na02f80 g543031 ( .a(n_25995), .b(x_in_36_10), .o(n_26934) );
in01f80 g543032 ( .a(n_26289), .o(n_26290) );
no02f80 g543033 ( .a(n_25995), .b(x_in_36_10), .o(n_26289) );
na02f80 g543034 ( .a(n_25460), .b(n_25459), .o(n_25461) );
no02f80 g543035 ( .a(n_25194), .b(n_25193), .o(n_25195) );
na02f80 g543036 ( .a(n_24887), .b(n_25193), .o(n_26113) );
no02f80 g543037 ( .a(n_27299), .b(n_27298), .o(n_27300) );
in01f80 g543038 ( .a(n_26287), .o(n_26288) );
no02f80 g543039 ( .a(n_25994), .b(x_in_20_10), .o(n_26287) );
na02f80 g543040 ( .a(n_25994), .b(x_in_20_10), .o(n_26933) );
no02f80 g543041 ( .a(n_25191), .b(n_25190), .o(n_25192) );
na02f80 g543042 ( .a(n_24886), .b(n_25190), .o(n_26110) );
no02f80 g543043 ( .a(n_27673), .b(n_27672), .o(n_27674) );
no02f80 g543044 ( .a(n_27489), .b(n_27488), .o(n_27490) );
na02f80 g543045 ( .a(n_25188), .b(x_in_26_12), .o(n_26029) );
na02f80 g543046 ( .a(n_25189), .b(x_in_52_10), .o(n_26028) );
in01f80 g543047 ( .a(n_25457), .o(n_25458) );
no02f80 g543048 ( .a(n_25189), .b(x_in_52_10), .o(n_25457) );
in01f80 g543049 ( .a(n_25455), .o(n_25456) );
no02f80 g543050 ( .a(n_25188), .b(x_in_26_12), .o(n_25455) );
no02f80 g543051 ( .a(n_26285), .b(n_26284), .o(n_26286) );
no02f80 g543052 ( .a(n_26893), .b(n_26892), .o(n_26894) );
na02f80 g543053 ( .a(n_25454), .b(x_in_12_11), .o(n_26315) );
in01f80 g543054 ( .a(n_25762), .o(n_25763) );
no02f80 g543055 ( .a(n_25454), .b(x_in_12_11), .o(n_25762) );
na02f80 g543056 ( .a(n_26588), .b(x_in_44_13), .o(n_27362) );
in01f80 g543057 ( .a(n_26890), .o(n_26891) );
no02f80 g543058 ( .a(n_26588), .b(x_in_44_13), .o(n_26890) );
in01f80 g543059 ( .a(n_25992), .o(n_25993) );
na02f80 g543060 ( .a(n_25761), .b(n_25107), .o(n_25992) );
no02f80 g543061 ( .a(n_27292), .b(n_27291), .o(n_27293) );
na02f80 g543062 ( .a(n_25187), .b(x_in_58_12), .o(n_26025) );
na02f80 g543063 ( .a(n_25991), .b(x_in_60_10), .o(n_26932) );
in01f80 g543064 ( .a(n_26282), .o(n_26283) );
no02f80 g543065 ( .a(n_25991), .b(x_in_60_10), .o(n_26282) );
na02f80 g543066 ( .a(n_24884), .b(n_24883), .o(n_24885) );
no02f80 g543067 ( .a(n_24943), .b(n_24548), .o(n_24549) );
no02f80 g543068 ( .a(n_25535), .b(n_25185), .o(n_25186) );
na02f80 g543069 ( .a(n_25184), .b(n_14479), .o(n_25820) );
na02f80 g543070 ( .a(n_25734), .b(FE_OFN290_n_27194), .o(n_26929) );
no02f80 g543071 ( .a(n_25263), .b(n_24881), .o(n_24882) );
no02f80 g543072 ( .a(n_24942), .b(n_24546), .o(n_24547) );
no02f80 g543073 ( .a(n_25806), .b(n_25452), .o(n_25453) );
no02f80 g543074 ( .a(n_24941), .b(n_24544), .o(n_24545) );
no02f80 g543075 ( .a(n_25262), .b(n_24879), .o(n_24880) );
no02f80 g543076 ( .a(n_24627), .b(n_24198), .o(n_24199) );
na02f80 g543077 ( .a(FE_OFN40_n_25450), .b(n_24742), .o(n_25451) );
in01f80 g543078 ( .a(n_25449), .o(n_26248) );
na02f80 g543079 ( .a(n_24508), .b(n_25183), .o(n_25449) );
na02f80 g543080 ( .a(n_25221), .b(n_25448), .o(n_25182) );
in01f80 g543081 ( .a(n_25760), .o(n_26543) );
na02f80 g543082 ( .a(n_24829), .b(n_25448), .o(n_25760) );
na02f80 g543083 ( .a(n_24892), .b(n_25181), .o(n_24878) );
in01f80 g543084 ( .a(n_25447), .o(n_26252) );
na02f80 g543085 ( .a(n_24510), .b(n_25181), .o(n_25447) );
na02f80 g543086 ( .a(n_24891), .b(n_25180), .o(n_24877) );
in01f80 g543087 ( .a(n_25446), .o(n_26250) );
na02f80 g543088 ( .a(n_24509), .b(n_25180), .o(n_25446) );
na02f80 g543089 ( .a(n_24890), .b(n_25183), .o(n_24876) );
in01f80 g543090 ( .a(n_25445), .o(n_26246) );
na02f80 g543091 ( .a(n_24504), .b(n_25179), .o(n_25445) );
na02f80 g543092 ( .a(n_24888), .b(n_25178), .o(n_24875) );
in01f80 g543093 ( .a(n_25444), .o(n_26244) );
na02f80 g543094 ( .a(n_24503), .b(n_25178), .o(n_25444) );
na02f80 g543095 ( .a(n_24889), .b(n_25179), .o(n_24874) );
na02f80 g543096 ( .a(n_25201), .b(n_25443), .o(n_25177) );
in01f80 g543097 ( .a(n_25759), .o(n_26693) );
na02f80 g543098 ( .a(n_24828), .b(n_25443), .o(n_25759) );
no02f80 g543099 ( .a(n_25533), .b(n_25175), .o(n_25176) );
no02f80 g543100 ( .a(n_24938), .b(n_24542), .o(n_24543) );
no02f80 g543101 ( .a(n_24937), .b(n_24540), .o(n_24541) );
no02f80 g543102 ( .a(n_25989), .b(n_25988), .o(n_25990) );
in01f80 g543103 ( .a(n_25987), .o(n_26610) );
na02f80 g543104 ( .a(n_25758), .b(n_25988), .o(n_25987) );
na02f80 g543105 ( .a(n_24936), .b(n_24538), .o(n_24539) );
no02f80 g543106 ( .a(n_24935), .b(n_24536), .o(n_24537) );
no02f80 g543107 ( .a(n_24934), .b(n_24534), .o(n_24535) );
na02f80 g543108 ( .a(n_24931), .b(n_24532), .o(n_24533) );
no02f80 g543109 ( .a(n_25184), .b(n_25173), .o(n_25174) );
no02f80 g543110 ( .a(n_25253), .b(n_24872), .o(n_24873) );
no02f80 g543111 ( .a(n_24181), .b(n_24872), .o(n_25867) );
no02f80 g543112 ( .a(n_27282), .b(FE_OFN492_n_28765), .o(n_27283) );
na02f80 g543113 ( .a(n_24196), .b(n_24195), .o(n_24197) );
na02f80 g543114 ( .a(n_24827), .b(FE_OFN1123_rst), .o(n_26021) );
in01f80 g543115 ( .a(n_24871), .o(n_25536) );
no02f80 g543116 ( .a(n_24531), .b(FE_OFN368_n_26312), .o(n_24871) );
in01f80 g543117 ( .a(n_25757), .o(n_26309) );
no02f80 g543118 ( .a(n_25442), .b(FE_OFN318_n_27400), .o(n_25757) );
no02f80 g543119 ( .a(n_25171), .b(n_25170), .o(n_25172) );
no02f80 g543120 ( .a(n_25171), .b(n_24735), .o(n_26365) );
na02f80 g543121 ( .a(n_24869), .b(n_25169), .o(n_24870) );
in01f80 g543122 ( .a(n_25441), .o(n_26091) );
no02f80 g543123 ( .a(n_25220), .b(n_25169), .o(n_25441) );
na02f80 g543124 ( .a(n_25167), .b(n_25439), .o(n_25168) );
in01f80 g543125 ( .a(n_25756), .o(n_26362) );
no02f80 g543126 ( .a(n_25440), .b(n_25439), .o(n_25756) );
na02f80 g543127 ( .a(n_25165), .b(n_25164), .o(n_25166) );
na02f80 g543128 ( .a(n_25165), .b(n_24731), .o(n_26090) );
na02f80 g543129 ( .a(n_25162), .b(n_25161), .o(n_25163) );
na02f80 g543130 ( .a(n_25162), .b(n_24730), .o(n_26089) );
no02f80 g543131 ( .a(n_25754), .b(n_25753), .o(n_25755) );
in01f80 g543132 ( .a(n_25752), .o(n_26313) );
na02f80 g543133 ( .a(n_25438), .b(n_25753), .o(n_25752) );
na02f80 g543134 ( .a(n_24867), .b(n_25160), .o(n_24868) );
in01f80 g543135 ( .a(n_25437), .o(n_26086) );
no02f80 g543136 ( .a(n_25197), .b(n_25160), .o(n_25437) );
na02f80 g543137 ( .a(n_24865), .b(n_25159), .o(n_24866) );
in01f80 g543138 ( .a(n_25436), .o(n_26083) );
no02f80 g543139 ( .a(n_25196), .b(n_25159), .o(n_25436) );
na02f80 g543140 ( .a(n_24863), .b(n_25158), .o(n_24864) );
in01f80 g543141 ( .a(n_25435), .o(n_26080) );
no02f80 g543142 ( .a(n_25188), .b(n_25158), .o(n_25435) );
na02f80 g543143 ( .a(n_25156), .b(n_25155), .o(n_25157) );
na02f80 g543144 ( .a(n_25156), .b(n_24729), .o(n_26079) );
na02f80 g543145 ( .a(n_25153), .b(n_25434), .o(n_25154) );
no02f80 g543146 ( .a(n_25504), .b(n_25434), .o(n_26355) );
in01f80 g543147 ( .a(n_26024), .o(n_26319) );
oa12f80 g543148 ( .a(n_24516), .b(n_24718), .c(n_6736), .o(n_26024) );
na02f80 g543149 ( .a(n_24861), .b(n_25152), .o(n_24862) );
in01f80 g543150 ( .a(n_25856), .o(n_25433) );
no02f80 g543151 ( .a(n_25198), .b(n_25152), .o(n_25856) );
na02f80 g543152 ( .a(n_25150), .b(n_25149), .o(n_25151) );
na02f80 g543153 ( .a(n_25150), .b(n_24725), .o(n_26077) );
na02f80 g543154 ( .a(n_25750), .b(n_25749), .o(n_25751) );
na02f80 g543155 ( .a(n_25750), .b(n_25377), .o(n_26632) );
no02f80 g543156 ( .a(n_25147), .b(n_25146), .o(n_25148) );
na02f80 g543157 ( .a(n_24859), .b(n_25146), .o(n_24860) );
na02f80 g543158 ( .a(n_25431), .b(n_25430), .o(n_25432) );
na02f80 g543159 ( .a(n_25431), .b(n_25047), .o(n_26350) );
no02f80 g543160 ( .a(n_24857), .b(n_24856), .o(n_24858) );
no02f80 g543161 ( .a(n_24857), .b(n_24409), .o(n_26072) );
na02f80 g543162 ( .a(n_25747), .b(n_25985), .o(n_25748) );
no02f80 g543163 ( .a(n_26003), .b(n_25985), .o(n_25986) );
na02f80 g543164 ( .a(n_25983), .b(n_25982), .o(n_25984) );
na02f80 g543165 ( .a(n_25983), .b(n_25708), .o(n_27211) );
na02f80 g543166 ( .a(n_24529), .b(n_24855), .o(n_24530) );
in01f80 g543167 ( .a(n_25569), .o(n_25145) );
no02f80 g543168 ( .a(n_24893), .b(n_24855), .o(n_25569) );
no02f80 g543169 ( .a(n_24853), .b(n_24852), .o(n_24854) );
no02f80 g543170 ( .a(n_24853), .b(n_24405), .o(n_26068) );
na02f80 g543171 ( .a(n_25428), .b(n_25746), .o(n_25429) );
no02f80 g543172 ( .a(n_25792), .b(n_25746), .o(n_26627) );
in01f80 g543173 ( .a(n_28080), .o(n_27850) );
oa12f80 g543174 ( .a(n_25105), .b(n_27210), .c(n_24745), .o(n_28080) );
in01f80 g543175 ( .a(n_28203), .o(n_27983) );
oa12f80 g543176 ( .a(n_25735), .b(n_25382), .c(n_27405), .o(n_28203) );
in01f80 g543177 ( .a(n_28200), .o(n_27982) );
oa12f80 g543178 ( .a(n_25134), .b(n_24812), .c(n_27428), .o(n_28200) );
in01f80 g543179 ( .a(n_28195), .o(n_27981) );
oa12f80 g543180 ( .a(n_25421), .b(n_25087), .c(n_27427), .o(n_28195) );
in01f80 g543181 ( .a(n_28192), .o(n_27980) );
oa12f80 g543182 ( .a(n_25420), .b(n_25085), .c(n_27425), .o(n_28192) );
in01f80 g543183 ( .a(n_28189), .o(n_27979) );
oa12f80 g543184 ( .a(n_25419), .b(n_25083), .c(n_27424), .o(n_28189) );
in01f80 g543185 ( .a(n_27923), .o(n_27671) );
oa12f80 g543186 ( .a(n_25418), .b(n_25081), .c(n_26992), .o(n_27923) );
in01f80 g543187 ( .a(n_28076), .o(n_27849) );
oa12f80 g543188 ( .a(n_25132), .b(n_27228), .c(n_24803), .o(n_28076) );
in01f80 g543189 ( .a(n_28073), .o(n_27848) );
oa12f80 g543190 ( .a(n_25131), .b(n_27227), .c(n_24801), .o(n_28073) );
in01f80 g543191 ( .a(n_28070), .o(n_27847) );
oa12f80 g543192 ( .a(n_25130), .b(n_27226), .c(n_24799), .o(n_28070) );
in01f80 g543193 ( .a(n_28067), .o(n_27846) );
oa12f80 g543194 ( .a(n_25417), .b(n_27225), .c(n_25079), .o(n_28067) );
in01f80 g543195 ( .a(n_27785), .o(n_27484) );
oa12f80 g543196 ( .a(n_25416), .b(n_25077), .c(n_26704), .o(n_27785) );
in01f80 g543197 ( .a(n_27845), .o(n_28271) );
ao12f80 g543198 ( .a(n_23161), .b(n_23789), .c(n_27656), .o(n_27845) );
in01f80 g543199 ( .a(n_27670), .o(n_28136) );
oa12f80 g543200 ( .a(n_24070), .b(n_23443), .c(n_27471), .o(n_27670) );
in01f80 g543201 ( .a(n_28064), .o(n_27844) );
oa12f80 g543202 ( .a(n_25415), .b(n_25064), .c(n_27223), .o(n_28064) );
in01f80 g543203 ( .a(n_28061), .o(n_27843) );
oa12f80 g543204 ( .a(n_25127), .b(n_24795), .c(n_27222), .o(n_28061) );
in01f80 g543205 ( .a(n_28186), .o(n_27978) );
oa12f80 g543206 ( .a(n_25413), .b(n_25073), .c(n_27420), .o(n_28186) );
in01f80 g543207 ( .a(n_28183), .o(n_27977) );
oa12f80 g543208 ( .a(n_25414), .b(n_25071), .c(n_27409), .o(n_28183) );
in01f80 g543209 ( .a(n_27777), .o(n_27481) );
oa12f80 g543210 ( .a(n_24848), .b(n_26703), .c(n_24485), .o(n_27777) );
in01f80 g543211 ( .a(n_28178), .o(n_27976) );
oa12f80 g543212 ( .a(n_25126), .b(n_24792), .c(n_27421), .o(n_28178) );
in01f80 g543213 ( .a(n_27780), .o(n_27480) );
oa12f80 g543214 ( .a(n_25125), .b(n_24789), .c(n_26701), .o(n_27780) );
in01f80 g543215 ( .a(n_28057), .o(n_27841) );
oa12f80 g543216 ( .a(n_25114), .b(n_24787), .c(n_27221), .o(n_28057) );
in01f80 g543217 ( .a(n_28054), .o(n_27840) );
oa12f80 g543218 ( .a(n_25124), .b(n_24785), .c(n_27220), .o(n_28054) );
in01f80 g543219 ( .a(n_28051), .o(n_27839) );
oa12f80 g543220 ( .a(n_25123), .b(n_24768), .c(n_27219), .o(n_28051) );
in01f80 g543221 ( .a(n_28174), .o(n_27975) );
oa12f80 g543222 ( .a(n_25133), .b(n_24783), .c(n_27417), .o(n_28174) );
in01f80 g543223 ( .a(n_27669), .o(n_28134) );
ao12f80 g543224 ( .a(n_22103), .b(n_27469), .c(n_22697), .o(n_27669) );
in01f80 g543225 ( .a(n_28048), .o(n_27838) );
oa12f80 g543226 ( .a(n_25738), .b(n_25393), .c(n_27218), .o(n_28048) );
in01f80 g543227 ( .a(n_27920), .o(n_27668) );
oa12f80 g543228 ( .a(n_25122), .b(n_24781), .c(n_26989), .o(n_27920) );
in01f80 g543229 ( .a(n_28386), .o(n_28239) );
oa12f80 g543230 ( .a(n_25412), .b(n_25068), .c(n_27799), .o(n_28386) );
in01f80 g543231 ( .a(n_28170), .o(n_27974) );
oa12f80 g543232 ( .a(n_25121), .b(n_24778), .c(n_27414), .o(n_28170) );
in01f80 g543233 ( .a(n_28043), .o(n_27837) );
oa12f80 g543234 ( .a(n_25120), .b(n_24776), .c(n_27217), .o(n_28043) );
in01f80 g543235 ( .a(n_28165), .o(n_27973) );
oa12f80 g543236 ( .a(n_25119), .b(n_24774), .c(n_27413), .o(n_28165) );
in01f80 g543237 ( .a(n_28040), .o(n_27836) );
oa12f80 g543238 ( .a(n_25118), .b(n_24772), .c(n_27216), .o(n_28040) );
in01f80 g543239 ( .a(n_28162), .o(n_27972) );
oa12f80 g543240 ( .a(n_25117), .b(n_24770), .c(n_27412), .o(n_28162) );
in01f80 g543241 ( .a(n_27917), .o(n_27666) );
oa12f80 g543242 ( .a(n_25411), .b(n_25066), .c(n_26988), .o(n_27917) );
in01f80 g543243 ( .a(n_27605), .o(n_27276) );
oa12f80 g543244 ( .a(n_25116), .b(n_24764), .c(n_26465), .o(n_27605) );
in01f80 g543245 ( .a(n_27914), .o(n_27665) );
oa12f80 g543246 ( .a(n_25410), .b(n_25062), .c(n_26987), .o(n_27914) );
in01f80 g543247 ( .a(n_28159), .o(n_27971) );
oa12f80 g543248 ( .a(n_25115), .b(n_24761), .c(n_27411), .o(n_28159) );
in01f80 g543249 ( .a(n_27773), .o(n_27478) );
oa12f80 g543250 ( .a(n_25737), .b(n_25390), .c(n_26700), .o(n_27773) );
in01f80 g543251 ( .a(n_27770), .o(n_27477) );
oa12f80 g543252 ( .a(n_25113), .b(n_24759), .c(n_26699), .o(n_27770) );
in01f80 g543253 ( .a(n_27833), .o(n_28269) );
oa12f80 g543254 ( .a(n_24978), .b(n_27654), .c(n_24236), .o(n_27833) );
in01f80 g543255 ( .a(n_27275), .o(n_27898) );
oa12f80 g543256 ( .a(n_23678), .b(n_27079), .c(n_23066), .o(n_27275) );
oa12f80 g543257 ( .a(n_14281), .b(n_24851), .c(n_13123), .o(n_25839) );
in01f80 g543258 ( .a(n_28154), .o(n_27967) );
oa12f80 g543259 ( .a(n_25112), .b(n_27410), .c(n_24757), .o(n_28154) );
in01f80 g543260 ( .a(n_27662), .o(n_28132) );
oa12f80 g543261 ( .a(n_24059), .b(n_23426), .c(n_27467), .o(n_27662) );
in01f80 g543262 ( .a(n_28285), .o(n_28100) );
oa12f80 g543263 ( .a(n_25980), .b(n_25720), .c(n_27626), .o(n_28285) );
in01f80 g543264 ( .a(n_28026), .o(n_27832) );
oa12f80 g543265 ( .a(n_25977), .b(n_25718), .c(n_27229), .o(n_28026) );
in01f80 g543266 ( .a(n_28151), .o(n_27966) );
oa12f80 g543267 ( .a(n_25109), .b(n_27408), .c(n_24752), .o(n_28151) );
in01f80 g543268 ( .a(n_28282), .o(n_28099) );
oa12f80 g543269 ( .a(n_26263), .b(n_25948), .c(n_27625), .o(n_28282) );
in01f80 g543270 ( .a(n_27389), .o(n_27085) );
oa12f80 g543271 ( .a(n_24841), .b(n_26192), .c(n_24458), .o(n_27389) );
in01f80 g543272 ( .a(n_28148), .o(n_27965) );
oa12f80 g543273 ( .a(n_25108), .b(n_27407), .c(n_24748), .o(n_28148) );
in01f80 g543274 ( .a(n_27767), .o(n_27476) );
oa12f80 g543275 ( .a(n_25409), .b(n_25056), .c(n_26696), .o(n_27767) );
in01f80 g543276 ( .a(n_27661), .o(n_28130) );
oa12f80 g543277 ( .a(n_25300), .b(n_27465), .c(n_24654), .o(n_27661) );
in01f80 g543278 ( .a(n_27660), .o(n_28128) );
oa12f80 g543279 ( .a(n_24056), .b(n_23422), .c(n_27463), .o(n_27660) );
in01f80 g543280 ( .a(n_28145), .o(n_27964) );
oa12f80 g543281 ( .a(n_25739), .b(n_25380), .c(n_27404), .o(n_28145) );
oa12f80 g543282 ( .a(n_25143), .b(n_815), .c(FE_OFN92_n_27449), .o(n_25144) );
ao22s80 g543283 ( .a(n_24191), .b(n_24438), .c(x_out_55_30), .d(FE_OFN318_n_27400), .o(n_25142) );
oa12f80 g543284 ( .a(n_25104), .b(n_402), .c(FE_OFN1181_rst), .o(n_25745) );
oa12f80 g543285 ( .a(n_25513), .b(n_343), .c(FE_OFN1109_rst), .o(n_25427) );
oa12f80 g543286 ( .a(n_26219), .b(n_25715), .c(n_25029), .o(n_26580) );
oa12f80 g543287 ( .a(n_25139), .b(n_1949), .c(FE_OFN1174_n_4860), .o(n_25141) );
oa12f80 g543288 ( .a(n_25139), .b(n_1629), .c(FE_OFN1174_n_4860), .o(n_25140) );
na02f80 g543289 ( .a(n_25733), .b(n_25716), .o(n_26606) );
oa22f80 g543290 ( .a(n_24167), .b(n_24108), .c(n_1295), .d(FE_OFN89_n_27449), .o(n_24850) );
ao22s80 g543291 ( .a(n_25424), .b(FE_OFN454_n_24837), .c(x_out_48_31), .d(FE_OFN1179_n_17184), .o(n_25425) );
na03f80 g543292 ( .a(n_4409), .b(n_24192), .c(FE_OFN60_n_27012), .o(n_25810) );
ao22s80 g543293 ( .a(n_24072), .b(n_27656), .c(n_24071), .d(n_27224), .o(n_27657) );
oa12f80 g543294 ( .a(n_24526), .b(n_24525), .c(x_in_38_15), .o(n_28863) );
ao22s80 g543295 ( .a(n_24358), .b(n_27471), .c(n_24357), .d(n_26991), .o(n_27472) );
oa12f80 g543296 ( .a(n_24520), .b(n_24527), .c(n_24838), .o(n_25830) );
ao22s80 g543297 ( .a(n_27469), .b(n_23019), .c(n_26990), .d(n_23018), .o(n_27470) );
in01f80 g543298 ( .a(n_25137), .o(n_25138) );
oa22f80 g543299 ( .a(n_24126), .b(n_9113), .c(n_8331), .d(n_5983), .o(n_25137) );
ao12f80 g543300 ( .a(n_26840), .b(n_26839), .c(n_26838), .o(n_27268) );
ao12f80 g543301 ( .a(n_26554), .b(n_26553), .c(n_26552), .o(n_27081) );
oa12f80 g543302 ( .a(n_26550), .b(n_26555), .c(n_26831), .o(n_27579) );
ao22s80 g543303 ( .a(n_27654), .b(n_25275), .c(n_27212), .d(n_25274), .o(n_27655) );
ao22s80 g543304 ( .a(n_27079), .b(n_23974), .c(n_26461), .d(n_23973), .o(n_27080) );
ao12f80 g543305 ( .a(n_25103), .b(n_25102), .c(n_25101), .o(n_25744) );
in01f80 g543306 ( .a(n_25814), .o(n_25423) );
oa12f80 g543307 ( .a(n_24524), .b(n_24851), .c(n_24523), .o(n_25814) );
ao22s80 g543308 ( .a(n_24349), .b(n_27467), .c(n_24348), .d(n_26986), .o(n_27468) );
oa22f80 g543309 ( .a(n_24849), .b(n_463), .c(n_24518), .d(x_in_28_15), .o(n_28798) );
ao22s80 g543310 ( .a(n_27465), .b(n_25574), .c(n_26985), .d(n_25573), .o(n_27466) );
ao22s80 g543311 ( .a(n_24344), .b(n_27463), .c(n_24343), .d(n_26984), .o(n_27464) );
oa12f80 g543312 ( .a(n_24522), .b(n_24839), .c(n_24521), .o(n_25822) );
oa22f80 g543313 ( .a(n_25040), .b(FE_OFN265_n_4280), .c(n_1716), .d(FE_OFN1181_rst), .o(n_25743) );
oa22f80 g543314 ( .a(n_24404), .b(FE_OFN405_n_28303), .c(n_1462), .d(FE_OFN1110_rst), .o(n_25136) );
oa22f80 g543315 ( .a(n_26983), .b(FE_OFN266_n_4280), .c(n_630), .d(n_29104), .o(n_27462) );
oa22f80 g543316 ( .a(n_26692), .b(FE_OFN266_n_4280), .c(n_1408), .d(FE_OFN56_n_27012), .o(n_27267) );
oa22f80 g543317 ( .a(n_26690), .b(FE_OFN251_n_4162), .c(n_1508), .d(FE_OFN93_n_27449), .o(n_27265) );
oa22f80 g543318 ( .a(n_24835), .b(FE_OFN409_n_28303), .c(n_695), .d(FE_OFN125_n_27449), .o(n_25135) );
oa22f80 g543319 ( .a(n_26190), .b(FE_OFN266_n_4280), .c(n_1400), .d(n_29261), .o(n_26850) );
oa22f80 g543320 ( .a(FE_OFN430_n_26458), .b(n_4280), .c(n_993), .d(n_29261), .o(n_27076) );
oa22f80 g543321 ( .a(n_25039), .b(FE_OFN212_n_29661), .c(n_1084), .d(FE_OFN352_n_4860), .o(n_25741) );
ao22s80 g543322 ( .a(n_24717), .b(n_25090), .c(x_out_34_31), .d(FE_OFN195_n_5003), .o(n_25740) );
oa22f80 g543323 ( .a(n_26189), .b(FE_OFN211_n_29661), .c(n_451), .d(FE_OFN360_n_4860), .o(n_26847) );
oa22f80 g543324 ( .a(n_26981), .b(FE_OFN412_n_28303), .c(n_715), .d(FE_OFN113_n_27449), .o(n_27461) );
oa22f80 g543325 ( .a(n_26187), .b(FE_OFN409_n_28303), .c(n_344), .d(rst), .o(n_26843) );
oa22f80 g543326 ( .a(n_24715), .b(FE_OFN409_n_28303), .c(n_1180), .d(FE_OFN125_n_27449), .o(n_25422) );
oa22f80 g543327 ( .a(n_26687), .b(FE_OFN244_n_4162), .c(n_530), .d(FE_OFN108_n_27449), .o(n_27264) );
oa22f80 g543328 ( .a(n_26683), .b(FE_OFN244_n_4162), .c(n_1846), .d(FE_OFN11_n_29204), .o(n_27261) );
oa22f80 g543329 ( .a(n_26685), .b(FE_OFN249_n_4162), .c(n_1964), .d(FE_OFN12_n_29204), .o(n_27260) );
na02f80 g543355 ( .a(n_25739), .b(n_25381), .o(n_27540) );
na02f80 g543356 ( .a(n_25134), .b(n_24813), .o(n_27537) );
na02f80 g543357 ( .a(n_25421), .b(n_25088), .o(n_27534) );
na02f80 g543358 ( .a(n_26555), .b(x_in_8_14), .o(n_27340) );
in01f80 g543359 ( .a(n_26841), .o(n_26842) );
no02f80 g543360 ( .a(n_26555), .b(x_in_8_14), .o(n_26841) );
na02f80 g543361 ( .a(n_25420), .b(n_25086), .o(n_27529) );
na02f80 g543362 ( .a(n_24848), .b(n_24486), .o(n_26914) );
no02f80 g543363 ( .a(n_24846), .b(FE_OFN23_n_26609), .o(n_24847) );
na02f80 g543364 ( .a(n_25419), .b(n_25084), .o(n_27526) );
na02f80 g543365 ( .a(n_25133), .b(n_24784), .o(n_27514) );
na02f80 g543366 ( .a(n_25418), .b(n_25082), .o(n_27144) );
na02f80 g543367 ( .a(n_25132), .b(n_24804), .o(n_27338) );
na02f80 g543368 ( .a(n_25131), .b(n_24802), .o(n_27335) );
na02f80 g543369 ( .a(n_25130), .b(n_24800), .o(n_27332) );
na02f80 g543370 ( .a(n_25417), .b(n_25080), .o(n_27329) );
na02f80 g543371 ( .a(n_24527), .b(x_in_38_14), .o(n_25499) );
in01f80 g543372 ( .a(n_24844), .o(n_24845) );
no02f80 g543373 ( .a(n_24527), .b(x_in_38_14), .o(n_24844) );
na02f80 g543374 ( .a(n_24525), .b(x_in_38_15), .o(n_24526) );
na02f80 g543375 ( .a(n_25416), .b(n_25078), .o(n_26917) );
na02f80 g543376 ( .a(n_24843), .b(x_in_38_13), .o(n_25777) );
in01f80 g543377 ( .a(n_25128), .o(n_25129) );
no02f80 g543378 ( .a(n_24843), .b(x_in_38_13), .o(n_25128) );
na02f80 g543379 ( .a(n_25415), .b(n_25065), .o(n_27326) );
na02f80 g543380 ( .a(n_25127), .b(n_24796), .o(n_27323) );
na02f80 g543381 ( .a(n_25126), .b(n_24793), .o(n_27520) );
na02f80 g543382 ( .a(n_25414), .b(n_25072), .o(n_27517) );
na02f80 g543383 ( .a(n_25413), .b(n_25074), .o(n_27523) );
na02f80 g543384 ( .a(n_25125), .b(n_24790), .o(n_26911) );
na02f80 g543385 ( .a(n_25124), .b(n_24786), .o(n_27317) );
na02f80 g543386 ( .a(n_25123), .b(n_24769), .o(n_27314) );
na02f80 g543387 ( .a(n_25738), .b(n_25394), .o(n_27311) );
na02f80 g543388 ( .a(n_25122), .b(n_24782), .o(n_27141) );
na02f80 g543389 ( .a(n_25412), .b(n_25069), .o(n_27855) );
na02f80 g543390 ( .a(n_25121), .b(n_24779), .o(n_27511) );
na02f80 g543391 ( .a(n_25120), .b(n_24777), .o(n_27308) );
na02f80 g543392 ( .a(n_25119), .b(n_24775), .o(n_27508) );
na02f80 g543393 ( .a(n_25118), .b(n_24773), .o(n_27305) );
na02f80 g543394 ( .a(n_25117), .b(n_24771), .o(n_27505) );
na02f80 g543395 ( .a(n_25411), .b(n_25067), .o(n_27138) );
no02f80 g543396 ( .a(n_26839), .b(n_26838), .o(n_26840) );
na02f80 g543397 ( .a(n_25116), .b(n_24765), .o(n_26592) );
na02f80 g543398 ( .a(n_25410), .b(n_25063), .o(n_27135) );
na02f80 g543399 ( .a(n_25115), .b(n_24762), .o(n_27501) );
no02f80 g543400 ( .a(n_26553), .b(n_26552), .o(n_26554) );
in01f80 g543401 ( .a(n_26264), .o(n_26265) );
na02f80 g543402 ( .a(n_25981), .b(n_25723), .o(n_26264) );
na02f80 g543403 ( .a(n_25114), .b(n_24788), .o(n_27320) );
in01f80 g543404 ( .a(n_27069), .o(n_27070) );
na02f80 g543405 ( .a(n_26837), .b(n_26479), .o(n_27069) );
na02f80 g543406 ( .a(n_26836), .b(x_in_8_13), .o(n_27499) );
in01f80 g543407 ( .a(n_27067), .o(n_27068) );
no02f80 g543408 ( .a(n_26836), .b(x_in_8_13), .o(n_27067) );
na02f80 g543409 ( .a(n_25113), .b(n_24760), .o(n_26903) );
na02f80 g543410 ( .a(n_25980), .b(n_25721), .o(n_27677) );
na02f80 g543411 ( .a(n_25737), .b(n_25391), .o(n_26899) );
in01f80 g543412 ( .a(n_26834), .o(n_26835) );
na02f80 g543413 ( .a(n_26551), .b(n_26197), .o(n_26834) );
na02f80 g543414 ( .a(n_24851), .b(n_24523), .o(n_24524) );
in01f80 g543415 ( .a(n_27065), .o(n_27066) );
na02f80 g543416 ( .a(n_26833), .b(n_26477), .o(n_27065) );
na02f80 g543417 ( .a(n_25112), .b(n_24758), .o(n_27497) );
in01f80 g543418 ( .a(n_25978), .o(n_25979) );
na02f80 g543419 ( .a(n_25736), .b(n_25389), .o(n_25978) );
na02f80 g543420 ( .a(n_24842), .b(x_in_28_14), .o(n_25764) );
in01f80 g543421 ( .a(n_25110), .o(n_25111) );
no02f80 g543422 ( .a(n_24842), .b(x_in_28_14), .o(n_25110) );
na02f80 g543423 ( .a(n_25109), .b(n_24753), .o(n_27492) );
na02f80 g543424 ( .a(n_25977), .b(n_25719), .o(n_27299) );
na02f80 g543425 ( .a(n_25735), .b(n_25383), .o(n_27543) );
na02f80 g543426 ( .a(n_25108), .b(n_24749), .o(n_27489) );
na02f80 g543427 ( .a(n_26263), .b(n_25949), .o(n_27673) );
na02f80 g543428 ( .a(n_24841), .b(n_24459), .o(n_26285) );
na02f80 g543429 ( .a(n_25409), .b(n_25057), .o(n_26893) );
in01f80 g543430 ( .a(n_27063), .o(n_27064) );
na02f80 g543431 ( .a(n_26832), .b(n_26472), .o(n_27063) );
na02f80 g543432 ( .a(n_24840), .b(x_in_28_13), .o(n_25761) );
in01f80 g543433 ( .a(n_25106), .o(n_25107) );
no02f80 g543434 ( .a(n_24840), .b(x_in_28_13), .o(n_25106) );
na02f80 g543435 ( .a(n_25105), .b(n_24746), .o(n_27292) );
in01f80 g543436 ( .a(n_25733), .o(n_25734) );
oa12f80 g543437 ( .a(n_25034), .b(n_24695), .c(n_8958), .o(n_25733) );
na02f80 g543438 ( .a(n_26262), .b(n_26213), .o(n_27616) );
na02f80 g543439 ( .a(n_24839), .b(n_24521), .o(n_24522) );
na02f80 g543440 ( .a(n_24839), .b(n_24369), .o(n_25541) );
no02f80 g543441 ( .a(n_25049), .b(FE_OFN402_n_28303), .o(n_26016) );
na02f80 g543442 ( .a(n_26555), .b(n_26831), .o(n_26550) );
na02f80 g543443 ( .a(n_26456), .b(n_26831), .o(n_27282) );
na02f80 g543444 ( .a(n_24527), .b(n_24838), .o(n_24520) );
na02f80 g543445 ( .a(n_24403), .b(n_24838), .o(n_25817) );
na02f80 g543446 ( .a(n_24123), .b(FE_OFN1110_rst), .o(n_25143) );
in01f80 g543447 ( .a(FE_OFN40_n_25450), .o(n_25104) );
no02f80 g543448 ( .a(FE_OFN454_n_24837), .b(FE_OFN369_n_26312), .o(n_25450) );
na02f80 g543449 ( .a(n_24716), .b(n_15183), .o(n_25513) );
no02f80 g543450 ( .a(n_24138), .b(n_27400), .o(n_25516) );
na02f80 g543451 ( .a(n_24518), .b(n_27194), .o(n_25139) );
na02f80 g543452 ( .a(n_24191), .b(n_24190), .o(n_24192) );
no02f80 g543453 ( .a(n_25102), .b(n_25101), .o(n_25103) );
in01f80 g543454 ( .a(n_25100), .o(n_25813) );
na02f80 g543455 ( .a(n_24835), .b(n_25101), .o(n_25100) );
oa12f80 g543456 ( .a(n_13716), .b(n_23902), .c(n_14832), .o(n_24947) );
oa12f80 g543457 ( .a(n_15082), .b(n_23901), .c(n_15759), .o(n_24966) );
oa12f80 g543458 ( .a(n_13980), .b(n_24189), .c(n_14917), .o(n_25269) );
in01f80 g543459 ( .a(n_27653), .o(n_28122) );
ao12f80 g543460 ( .a(n_25342), .b(n_25932), .c(n_27454), .o(n_27653) );
oa12f80 g543461 ( .a(n_16108), .b(n_24188), .c(n_16689), .o(n_25268) );
ao12f80 g543462 ( .a(n_14960), .b(n_24187), .c(n_15549), .o(n_25266) );
ao12f80 g543463 ( .a(n_15481), .b(n_23583), .c(n_16260), .o(n_24640) );
ao12f80 g543464 ( .a(n_14957), .b(n_23900), .c(n_15545), .o(n_24962) );
oa12f80 g543465 ( .a(n_26179), .b(n_25617), .c(n_27046), .o(n_27739) );
ao12f80 g543466 ( .a(n_14955), .b(n_23899), .c(n_15544), .o(n_24960) );
ao12f80 g543467 ( .a(n_14950), .b(n_23898), .c(n_15543), .o(n_24958) );
oa12f80 g543468 ( .a(n_13643), .b(n_23897), .c(n_14729), .o(n_24956) );
ao12f80 g543469 ( .a(n_14948), .b(n_23896), .c(n_15541), .o(n_24954) );
ao12f80 g543470 ( .a(n_14940), .b(n_23895), .c(n_15537), .o(n_24952) );
in01f80 g543471 ( .a(n_26830), .o(n_27563) );
oa12f80 g543472 ( .a(n_25031), .b(n_24354), .c(n_26540), .o(n_26830) );
in01f80 g543473 ( .a(n_27459), .o(n_28003) );
oa12f80 g543474 ( .a(n_25930), .b(n_25306), .c(n_27255), .o(n_27459) );
in01f80 g543475 ( .a(n_27259), .o(n_27875) );
oa12f80 g543476 ( .a(n_25928), .b(n_25301), .c(n_27036), .o(n_27259) );
in01f80 g543477 ( .a(n_27258), .o(n_27872) );
oa12f80 g543478 ( .a(n_25030), .b(n_24350), .c(n_27033), .o(n_27258) );
ao12f80 g543479 ( .a(n_15782), .b(n_24834), .c(n_16488), .o(n_25463) );
ao12f80 g543480 ( .a(n_15495), .b(n_24833), .c(n_16248), .o(n_25460) );
oa12f80 g543481 ( .a(n_10618), .b(n_24183), .c(n_11819), .o(n_24561) );
oa12f80 g543482 ( .a(n_13639), .b(n_24186), .c(n_14675), .o(n_24884) );
oa12f80 g543483 ( .a(n_24719), .b(n_24720), .c(n_24107), .o(n_25099) );
oa12f80 g543484 ( .a(n_15128), .b(n_23894), .c(n_15824), .o(n_24943) );
oa12f80 g543485 ( .a(n_16130), .b(n_24517), .c(n_16693), .o(n_25535) );
oa12f80 g543486 ( .a(n_14297), .b(n_24185), .c(n_15109), .o(n_25263) );
oa12f80 g543487 ( .a(n_24515), .b(n_24514), .c(n_24513), .o(n_24516) );
ao12f80 g543488 ( .a(n_13195), .b(n_23893), .c(n_14387), .o(n_24942) );
oa12f80 g543489 ( .a(n_13193), .b(n_24832), .c(n_14361), .o(n_25806) );
oa22f80 g543490 ( .a(n_25406), .b(n_25405), .c(n_3668), .d(x_in_45_14), .o(n_25408) );
ao12f80 g543491 ( .a(n_15166), .b(n_23892), .c(n_15844), .o(n_24941) );
ao12f80 g543492 ( .a(n_15149), .b(n_24184), .c(n_15832), .o(n_25262) );
ao12f80 g543493 ( .a(n_13613), .b(n_23582), .c(n_14645), .o(n_24627) );
ao12f80 g543494 ( .a(n_13701), .b(n_24502), .c(n_14814), .o(n_25531) );
ao12f80 g543495 ( .a(x_in_57_15), .b(n_25724), .c(n_25976), .o(n_26602) );
oa12f80 g543496 ( .a(n_13948), .b(n_24512), .c(n_14929), .o(n_25533) );
oa12f80 g543497 ( .a(n_15097), .b(n_23891), .c(n_15785), .o(n_24938) );
oa12f80 g543498 ( .a(n_15091), .b(n_23890), .c(n_15778), .o(n_24937) );
oa12f80 g543499 ( .a(n_15512), .b(n_23889), .c(n_16254), .o(n_24936) );
oa12f80 g543500 ( .a(n_15088), .b(n_23888), .c(n_15772), .o(n_24935) );
ao12f80 g543501 ( .a(n_15119), .b(n_23887), .c(n_15809), .o(n_24934) );
oa12f80 g543502 ( .a(n_10639), .b(n_23886), .c(n_11780), .o(n_24931) );
oa12f80 g543503 ( .a(n_15023), .b(n_24511), .c(n_14086), .o(n_25184) );
ao12f80 g543504 ( .a(n_14094), .b(n_23581), .c(n_14806), .o(n_24196) );
ao12f80 g543505 ( .a(n_11413), .b(n_25406), .c(n_25405), .o(n_25407) );
in01f80 g543506 ( .a(n_25428), .o(n_25792) );
ao12f80 g543507 ( .a(n_24456), .b(n_24517), .c(n_24455), .o(n_25428) );
ao12f80 g543508 ( .a(n_24738), .b(n_24737), .c(n_24736), .o(n_25098) );
ao12f80 g543509 ( .a(n_26758), .b(n_26757), .c(n_26756), .o(n_27062) );
oa12f80 g543510 ( .a(n_24436), .b(n_24435), .c(n_24434), .o(n_25510) );
in01f80 g543511 ( .a(n_24886), .o(n_25191) );
ao12f80 g543512 ( .a(n_23883), .b(n_24183), .c(n_23882), .o(n_24886) );
ao12f80 g543513 ( .a(n_26755), .b(n_26754), .c(n_26753), .o(n_27061) );
oa12f80 g543514 ( .a(n_24734), .b(n_24733), .c(n_24732), .o(n_25789) );
ao12f80 g543515 ( .a(n_25379), .b(n_25402), .c(n_25378), .o(n_25732) );
ao12f80 g543516 ( .a(n_26752), .b(n_26751), .c(n_26750), .o(n_27060) );
ao12f80 g543517 ( .a(n_27005), .b(n_27004), .c(n_27003), .o(n_27257) );
ao22s80 g543518 ( .a(n_26182), .b(n_27454), .c(n_26181), .d(n_26979), .o(n_27455) );
oa12f80 g543519 ( .a(n_24147), .b(n_24146), .c(n_24433), .o(n_25227) );
ao12f80 g543520 ( .a(n_24809), .b(n_24820), .c(n_24808), .o(n_25097) );
ao12f80 g543521 ( .a(n_26749), .b(n_26748), .c(n_26747), .o(n_27059) );
oa12f80 g543522 ( .a(n_24145), .b(n_24144), .c(n_24432), .o(n_25224) );
ao12f80 g543523 ( .a(n_24431), .b(FE_OFN923_n_24430), .c(n_24429), .o(n_24831) );
ao12f80 g543524 ( .a(n_26746), .b(n_26745), .c(n_26744), .o(n_27058) );
in01f80 g543525 ( .a(n_25153), .o(n_25504) );
ao12f80 g543526 ( .a(n_24177), .b(n_24188), .c(n_24176), .o(n_25153) );
oa12f80 g543527 ( .a(n_24428), .b(n_24427), .c(n_24426), .o(n_25505) );
ao12f80 g543528 ( .a(n_26514), .b(n_26513), .c(n_26512), .o(n_26829) );
oa12f80 g543529 ( .a(n_24425), .b(n_24424), .c(n_24423), .o(n_25503) );
ao12f80 g543530 ( .a(n_26511), .b(n_26510), .c(n_26509), .o(n_26828) );
oa12f80 g543531 ( .a(n_24422), .b(n_24421), .c(n_24420), .o(n_25502) );
in01f80 g543532 ( .a(n_25171), .o(n_24830) );
oa12f80 g543533 ( .a(n_24174), .b(n_24189), .c(n_24173), .o(n_25171) );
ao12f80 g543534 ( .a(n_26212), .b(n_26211), .c(n_26210), .o(n_26548) );
ao12f80 g543535 ( .a(n_26507), .b(n_26506), .c(n_26505), .o(n_26827) );
ao12f80 g543536 ( .a(n_26742), .b(n_26741), .c(n_26740), .o(n_27057) );
oa12f80 g543537 ( .a(n_24143), .b(n_24142), .c(n_24419), .o(n_25223) );
ao12f80 g543538 ( .a(n_26736), .b(n_26735), .c(n_26734), .o(n_27056) );
ao12f80 g543539 ( .a(n_26504), .b(n_26503), .c(n_26502), .o(n_26826) );
oa12f80 g543540 ( .a(n_24728), .b(n_24727), .c(n_24726), .o(n_25780) );
ao12f80 g543541 ( .a(n_26209), .b(n_26208), .c(n_26466), .o(n_26547) );
ao12f80 g543542 ( .a(n_26739), .b(n_26738), .c(n_26737), .o(n_27055) );
oa12f80 g543543 ( .a(n_24453), .b(n_24452), .c(n_24740), .o(n_25498) );
ao12f80 g543544 ( .a(n_26500), .b(n_26499), .c(n_26498), .o(n_26825) );
ao12f80 g543545 ( .a(n_26497), .b(n_26496), .c(n_26495), .o(n_26824) );
in01f80 g543546 ( .a(n_24869), .o(n_25220) );
ao12f80 g543547 ( .a(n_23860), .b(n_23892), .c(n_23859), .o(n_24869) );
in01f80 g543548 ( .a(n_25221), .o(n_24829) );
oa12f80 g543549 ( .a(n_24172), .b(n_24187), .c(n_24171), .o(n_25221) );
in01f80 g543550 ( .a(n_24529), .o(n_24893) );
ao12f80 g543551 ( .a(n_23578), .b(n_23583), .c(n_23577), .o(n_24529) );
oa12f80 g543552 ( .a(n_24158), .b(n_24157), .c(n_24448), .o(n_25219) );
ao12f80 g543553 ( .a(n_25962), .b(n_25961), .c(n_25960), .o(n_26259) );
ao12f80 g543554 ( .a(n_26730), .b(n_26729), .c(n_26728), .o(n_27053) );
oa12f80 g543555 ( .a(n_24156), .b(n_24155), .c(n_24449), .o(n_25216) );
ao12f80 g543556 ( .a(n_26494), .b(n_26493), .c(n_26492), .o(n_26823) );
oa12f80 g543557 ( .a(n_24154), .b(n_24153), .c(n_24450), .o(n_25215) );
ao12f80 g543558 ( .a(n_26488), .b(n_26487), .c(n_26486), .o(n_26822) );
in01f80 g543559 ( .a(n_24892), .o(n_24510) );
oa12f80 g543560 ( .a(n_23881), .b(n_23900), .c(n_23880), .o(n_24892) );
ao12f80 g543561 ( .a(n_26491), .b(n_26490), .c(n_26489), .o(n_26821) );
ao22s80 g543562 ( .a(n_26446), .b(n_27046), .c(n_26445), .d(n_26440), .o(n_27047) );
ao12f80 g543563 ( .a(n_26207), .b(n_26206), .c(n_26205), .o(n_26546) );
ao12f80 g543564 ( .a(n_27235), .b(n_27234), .c(n_27233), .o(n_27446) );
oa12f80 g543565 ( .a(n_24152), .b(n_24151), .c(n_24454), .o(n_25214) );
ao12f80 g543566 ( .a(n_26475), .b(n_26474), .c(n_26473), .o(n_26820) );
in01f80 g543567 ( .a(n_24891), .o(n_24509) );
oa12f80 g543568 ( .a(n_23879), .b(n_23899), .c(n_23878), .o(n_24891) );
ao12f80 g543569 ( .a(n_26727), .b(n_26726), .c(n_26725), .o(n_27043) );
in01f80 g543570 ( .a(n_25167), .o(n_25440) );
ao12f80 g543571 ( .a(n_24162), .b(n_24184), .c(n_24161), .o(n_25167) );
in01f80 g543572 ( .a(n_24890), .o(n_24508) );
oa12f80 g543573 ( .a(n_23877), .b(n_23898), .c(n_23876), .o(n_24890) );
in01f80 g543574 ( .a(n_24853), .o(n_24507) );
oa12f80 g543575 ( .a(n_23862), .b(n_23893), .c(n_23861), .o(n_24853) );
ao12f80 g543576 ( .a(n_26485), .b(n_26484), .c(n_26483), .o(n_26819) );
in01f80 g543577 ( .a(n_25150), .o(n_25207) );
ao12f80 g543578 ( .a(n_23875), .b(n_23897), .c(n_23874), .o(n_25150) );
ao12f80 g543579 ( .a(n_25959), .b(n_25958), .c(n_25957), .o(n_26254) );
in01f80 g543580 ( .a(n_25758), .o(n_25989) );
ao12f80 g543581 ( .a(n_24744), .b(n_24832), .c(n_24743), .o(n_25758) );
ao12f80 g543582 ( .a(n_26204), .b(n_26203), .c(n_26202), .o(n_26545) );
ao12f80 g543583 ( .a(n_26482), .b(n_26481), .c(n_26480), .o(n_26818) );
ao12f80 g543584 ( .a(n_26724), .b(n_26723), .c(n_26722), .o(n_27042) );
oa12f80 g543585 ( .a(n_24160), .b(n_24159), .c(n_24451), .o(n_25222) );
in01f80 g543586 ( .a(n_24889), .o(n_24504) );
oa12f80 g543587 ( .a(n_23873), .b(n_23896), .c(n_23872), .o(n_24889) );
in01f80 g543588 ( .a(n_25165), .o(n_25204) );
ao12f80 g543589 ( .a(n_23864), .b(n_23894), .c(n_23863), .o(n_25165) );
ao12f80 g543590 ( .a(n_26721), .b(n_26720), .c(n_26719), .o(n_27041) );
in01f80 g543591 ( .a(n_24888), .o(n_24503) );
oa12f80 g543592 ( .a(n_23871), .b(n_23895), .c(n_23870), .o(n_24888) );
in01f80 g543593 ( .a(n_25201), .o(n_24828) );
oa12f80 g543594 ( .a(n_24169), .b(n_24186), .c(n_24168), .o(n_25201) );
in01f80 g543595 ( .a(FE_OFN606_n_25225), .o(n_24827) );
ao22s80 g543596 ( .a(n_23824), .b(n_15033), .c(n_24502), .d(n_15032), .o(n_25225) );
oa12f80 g543597 ( .a(n_24418), .b(n_24417), .c(n_24416), .o(n_25476) );
ao12f80 g543598 ( .a(n_26733), .b(n_26732), .c(n_26731), .o(n_27040) );
ao12f80 g543599 ( .a(n_26718), .b(n_26717), .c(n_26716), .o(n_27039) );
ao12f80 g543600 ( .a(n_24141), .b(n_24140), .c(n_24139), .o(n_24501) );
ao12f80 g543601 ( .a(n_25941), .b(n_25940), .c(n_26193), .o(n_26243) );
oa12f80 g543602 ( .a(n_24136), .b(n_24135), .c(n_24415), .o(n_25200) );
ao12f80 g543603 ( .a(n_26201), .b(n_26200), .c(n_26199), .o(n_26542) );
in01f80 g543604 ( .a(n_25162), .o(n_25199) );
ao12f80 g543605 ( .a(n_23850), .b(n_23887), .c(n_23849), .o(n_25162) );
oa12f80 g543606 ( .a(n_24724), .b(n_24723), .c(n_25048), .o(n_25768) );
in01f80 g543607 ( .a(n_25750), .o(n_25765) );
ao12f80 g543608 ( .a(n_24445), .b(n_24512), .c(n_24444), .o(n_25750) );
ao12f80 g543609 ( .a(n_24134), .b(n_24133), .c(n_24132), .o(n_24500) );
in01f80 g543610 ( .a(n_24859), .o(n_25147) );
ao12f80 g543611 ( .a(n_23869), .b(n_23868), .c(n_23867), .o(n_24859) );
oa12f80 g543612 ( .a(n_11855), .b(n_23560), .c(n_11466), .o(n_24182) );
ao22s80 g543613 ( .a(n_25369), .b(n_26540), .c(n_25368), .d(n_25925), .o(n_26541) );
ao22s80 g543614 ( .a(n_26177), .b(n_27255), .c(n_26176), .d(n_26678), .o(n_27256) );
in01f80 g543615 ( .a(n_25438), .o(n_25754) );
ao12f80 g543616 ( .a(n_24443), .b(n_24511), .c(n_24442), .o(n_25438) );
oa12f80 g543617 ( .a(n_24414), .b(n_24413), .c(n_24722), .o(n_25471) );
in01f80 g543618 ( .a(n_25431), .o(n_25495) );
ao12f80 g543619 ( .a(n_24164), .b(n_24185), .c(n_24163), .o(n_25431) );
in01f80 g543620 ( .a(n_24861), .o(n_25198) );
ao12f80 g543621 ( .a(n_23854), .b(n_23889), .c(n_23853), .o(n_24861) );
ao12f80 g543622 ( .a(n_25956), .b(n_25955), .c(n_25954), .o(n_26242) );
ao12f80 g543623 ( .a(n_23573), .b(n_23581), .c(n_23572), .o(n_24531) );
ao12f80 g543624 ( .a(n_25952), .b(n_25951), .c(n_25950), .o(n_26241) );
ao12f80 g543625 ( .a(n_26715), .b(n_26714), .c(n_26713), .o(n_27038) );
ao22s80 g543626 ( .a(n_26173), .b(n_27036), .c(n_26172), .d(n_26439), .o(n_27037) );
oa12f80 g543627 ( .a(n_25942), .b(n_25976), .c(n_25967), .o(n_26897) );
in01f80 g543628 ( .a(n_24867), .o(n_25197) );
ao12f80 g543629 ( .a(n_23858), .b(n_23891), .c(n_23857), .o(n_24867) );
ao12f80 g543630 ( .a(n_24412), .b(n_24411), .c(n_24410), .o(n_24826) );
in01f80 g543631 ( .a(n_24857), .o(n_24499) );
oa12f80 g543632 ( .a(n_23846), .b(n_23902), .c(n_23845), .o(n_24857) );
ao22s80 g543633 ( .a(n_25367), .b(n_27033), .c(n_25366), .d(n_26438), .o(n_27034) );
ao12f80 g543634 ( .a(n_26712), .b(n_26711), .c(n_26710), .o(n_27032) );
ao12f80 g543635 ( .a(n_25713), .b(n_25712), .c(n_25711), .o(n_25975) );
in01f80 g543636 ( .a(n_25983), .o(n_25996) );
ao12f80 g543637 ( .a(n_24755), .b(n_24834), .c(n_24754), .o(n_25983) );
ao12f80 g543638 ( .a(n_24150), .b(n_24149), .c(n_24148), .o(n_24498) );
in01f80 g543639 ( .a(n_24181), .o(n_25253) );
oa12f80 g543640 ( .a(n_23575), .b(n_23582), .c(n_23574), .o(n_24181) );
in01f80 g543641 ( .a(n_24865), .o(n_25196) );
ao12f80 g543642 ( .a(n_23856), .b(n_23890), .c(n_23855), .o(n_24865) );
oa12f80 g543643 ( .a(n_25046), .b(n_25070), .c(n_25376), .o(n_25995) );
in01f80 g543644 ( .a(n_25747), .o(n_26003) );
ao12f80 g543645 ( .a(n_24751), .b(n_24833), .c(n_24750), .o(n_25747) );
ao12f80 g543646 ( .a(n_26707), .b(n_26706), .c(n_26705), .o(n_27031) );
ao12f80 g543647 ( .a(n_24441), .b(n_24440), .c(n_24439), .o(n_25442) );
ao12f80 g543648 ( .a(n_24464), .b(n_24493), .c(n_24463), .o(n_24825) );
in01f80 g543649 ( .a(n_24887), .o(n_25194) );
ao12f80 g543650 ( .a(n_23848), .b(n_23886), .c(n_23847), .o(n_24887) );
ao12f80 g543651 ( .a(n_26709), .b(n_26708), .c(n_26993), .o(n_27030) );
oa12f80 g543652 ( .a(n_25045), .b(n_25044), .c(n_25375), .o(n_25994) );
ao12f80 g543653 ( .a(n_24462), .b(n_24496), .c(n_24461), .o(n_24824) );
ao12f80 g543654 ( .a(n_26996), .b(n_26995), .c(n_26994), .o(n_27253) );
in01f80 g543655 ( .a(n_24863), .o(n_25188) );
ao12f80 g543656 ( .a(n_23852), .b(n_23888), .c(n_23851), .o(n_24863) );
oa12f80 g543657 ( .a(n_24130), .b(n_24129), .c(n_24128), .o(n_25189) );
ao12f80 g543658 ( .a(n_24408), .b(FE_OFN942_n_24127), .c(n_24406), .o(n_24823) );
ao12f80 g543659 ( .a(n_25710), .b(n_25709), .c(n_25939), .o(n_25974) );
oa12f80 g543660 ( .a(n_24447), .b(n_24446), .c(n_24739), .o(n_25454) );
ao12f80 g543661 ( .a(n_26470), .b(n_26469), .c(n_26468), .o(n_26815) );
ao12f80 g543662 ( .a(n_25947), .b(n_25946), .c(n_25945), .o(n_26240) );
in01f80 g543663 ( .a(n_26588), .o(n_26239) );
oa12f80 g543664 ( .a(n_25714), .b(n_25725), .c(n_25943), .o(n_26588) );
ao12f80 g543665 ( .a(n_25052), .b(n_25092), .c(n_25051), .o(n_25404) );
in01f80 g543666 ( .a(n_25156), .o(n_25187) );
ao12f80 g543667 ( .a(n_23866), .b(n_23901), .c(n_23865), .o(n_25156) );
oa12f80 g543668 ( .a(n_25043), .b(n_25042), .c(n_25041), .o(n_25991) );
oa22f80 g543669 ( .a(n_24097), .b(FE_OFN251_n_4162), .c(n_1157), .d(FE_OFN119_n_27449), .o(n_24822) );
oa22f80 g543670 ( .a(FE_OFN1037_n_26168), .b(n_29683), .c(n_189), .d(FE_OFN94_n_27449), .o(n_26814) );
oa22f80 g543671 ( .a(n_24496), .b(FE_OFN247_n_4162), .c(n_1632), .d(FE_OFN128_n_27449), .o(n_24497) );
oa22f80 g543672 ( .a(FE_OFN436_n_26167), .b(n_29046), .c(n_1893), .d(n_27449), .o(n_26812) );
oa22f80 g543673 ( .a(n_25027), .b(FE_OFN244_n_4162), .c(n_87), .d(FE_OFN131_n_27449), .o(n_25731) );
oa22f80 g543674 ( .a(n_26165), .b(FE_OFN254_n_4280), .c(n_781), .d(FE_OFN1124_rst), .o(n_26811) );
oa22f80 g543675 ( .a(n_26435), .b(FE_OFN256_n_4280), .c(n_134), .d(FE_OFN1174_n_4860), .o(n_27028) );
oa22f80 g543676 ( .a(n_25924), .b(FE_OFN412_n_28303), .c(n_1259), .d(FE_OFN113_n_27449), .o(n_26539) );
oa22f80 g543677 ( .a(n_26674), .b(FE_OFN410_n_28303), .c(n_924), .d(FE_OFN127_n_27449), .o(n_27252) );
oa22f80 g543678 ( .a(n_24368), .b(FE_OFN244_n_4162), .c(n_1957), .d(FE_OFN1174_n_4860), .o(n_25096) );
oa22f80 g543679 ( .a(n_26164), .b(FE_OFN244_n_4162), .c(n_267), .d(FE_OFN80_n_27012), .o(n_26810) );
oa22f80 g543680 ( .a(n_24367), .b(FE_OFN269_n_4280), .c(n_1054), .d(FE_OFN1113_rst), .o(n_25095) );
oa22f80 g543681 ( .a(n_26163), .b(FE_OFN208_n_29661), .c(n_1268), .d(FE_OFN335_n_4860), .o(n_26809) );
oa22f80 g543682 ( .a(n_25923), .b(FE_OFN211_n_29661), .c(n_826), .d(FE_OFN350_n_4860), .o(n_26538) );
oa22f80 g543683 ( .a(n_25922), .b(FE_OFN308_n_3069), .c(n_1142), .d(FE_OFN326_n_4860), .o(n_26537) );
oa22f80 g543684 ( .a(n_24437), .b(FE_OFN171_n_22948), .c(n_1130), .d(FE_OFN65_n_27012), .o(n_24495) );
oa22f80 g543685 ( .a(n_25921), .b(FE_OFN292_n_3069), .c(n_819), .d(FE_OFN336_n_4860), .o(n_26536) );
oa22f80 g543686 ( .a(n_25920), .b(n_4280), .c(n_1208), .d(FE_OFN68_n_27012), .o(n_26535) );
oa22f80 g543687 ( .a(FE_OFN1045_n_26162), .b(n_29683), .c(n_1222), .d(FE_OFN64_n_27012), .o(n_26808) );
oa22f80 g543688 ( .a(n_25919), .b(FE_OFN248_n_4162), .c(n_665), .d(FE_OFN113_n_27449), .o(n_26534) );
oa22f80 g543689 ( .a(n_25918), .b(n_29683), .c(n_1606), .d(n_27449), .o(n_26533) );
oa22f80 g543690 ( .a(n_25911), .b(FE_OFN181_n_27681), .c(n_1482), .d(FE_OFN1119_rst), .o(n_26532) );
oa22f80 g543691 ( .a(n_25917), .b(n_27681), .c(n_1701), .d(FE_OFN1117_rst), .o(n_26530) );
oa22f80 g543692 ( .a(n_26152), .b(FE_OFN264_n_4280), .c(n_1275), .d(FE_OFN98_n_27449), .o(n_26806) );
oa22f80 g543693 ( .a(n_25698), .b(FE_OFN260_n_4280), .c(n_599), .d(FE_OFN125_n_27449), .o(n_26238) );
oa22f80 g543694 ( .a(n_26166), .b(FE_OFN253_n_4280), .c(n_1859), .d(FE_OFN350_n_4860), .o(n_26803) );
oa22f80 g543695 ( .a(n_25916), .b(n_29683), .c(n_1918), .d(FE_OFN94_n_27449), .o(n_26528) );
oa22f80 g543696 ( .a(n_25915), .b(FE_OFN1151_n_3069), .c(n_512), .d(FE_OFN60_n_27012), .o(n_26526) );
oa22f80 g543697 ( .a(n_25914), .b(n_29683), .c(n_258), .d(n_27449), .o(n_26524) );
oa22f80 g543698 ( .a(n_26161), .b(FE_OFN180_n_27681), .c(n_70), .d(FE_OFN134_n_27449), .o(n_26800) );
oa22f80 g543699 ( .a(n_26159), .b(n_27681), .c(n_782), .d(FE_OFN101_n_27449), .o(n_26799) );
oa22f80 g543700 ( .a(n_24131), .b(FE_OFN199_n_29637), .c(n_179), .d(FE_OFN115_n_27449), .o(n_24180) );
oa22f80 g543701 ( .a(n_26158), .b(FE_OFN402_n_28303), .c(n_113), .d(FE_OFN69_n_27012), .o(n_26796) );
oa22f80 g543702 ( .a(n_23844), .b(FE_OFN400_n_28303), .c(n_1547), .d(FE_OFN56_n_27012), .o(n_23885) );
oa22f80 g543703 ( .a(n_24493), .b(FE_OFN410_n_28303), .c(n_1145), .d(FE_OFN76_n_27012), .o(n_24494) );
oa22f80 g543704 ( .a(n_26157), .b(FE_OFN209_n_29661), .c(n_1345), .d(FE_OFN105_n_27449), .o(n_26794) );
oa22f80 g543705 ( .a(n_25697), .b(FE_OFN409_n_28303), .c(n_1832), .d(FE_OFN125_n_27449), .o(n_26237) );
oa22f80 g543706 ( .a(FE_OFN943_n_24127), .b(FE_OFN404_n_28303), .c(n_647), .d(n_28362), .o(n_24179) );
oa22f80 g543707 ( .a(n_26156), .b(FE_OFN264_n_4280), .c(n_589), .d(FE_OFN1106_rst), .o(n_26790) );
oa22f80 g543708 ( .a(n_25402), .b(FE_OFN3_n_28682), .c(n_1689), .d(FE_OFN131_n_27449), .o(n_25403) );
oa22f80 g543709 ( .a(n_25696), .b(n_28682), .c(n_395), .d(FE_OFN1120_rst), .o(n_26234) );
oa22f80 g543710 ( .a(n_26671), .b(FE_OFN313_n_3069), .c(n_1647), .d(FE_OFN139_n_27449), .o(n_27248) );
oa22f80 g543711 ( .a(n_25913), .b(FE_OFN294_n_3069), .c(n_1486), .d(FE_OFN133_n_27449), .o(n_26523) );
oa22f80 g543712 ( .a(n_26155), .b(FE_OFN411_n_28303), .c(n_430), .d(FE_OFN1114_rst), .o(n_26785) );
oa22f80 g543713 ( .a(n_26154), .b(FE_OFN405_n_28303), .c(n_639), .d(FE_OFN1106_rst), .o(n_26783) );
oa22f80 g543714 ( .a(n_24820), .b(FE_OFN416_n_28303), .c(n_1425), .d(FE_OFN1123_rst), .o(n_24821) );
oa22f80 g543715 ( .a(n_25912), .b(FE_OFN417_n_28303), .c(n_1664), .d(FE_OFN1124_rst), .o(n_26522) );
oa22f80 g543716 ( .a(n_23552), .b(FE_OFN214_n_29687), .c(n_1237), .d(FE_OFN104_n_27449), .o(n_24178) );
oa22f80 g543717 ( .a(n_25695), .b(FE_OFN417_n_28303), .c(n_1227), .d(FE_OFN142_n_27449), .o(n_26233) );
oa22f80 g543718 ( .a(n_25694), .b(FE_OFN404_n_28303), .c(n_1453), .d(FE_OFN78_n_27012), .o(n_26231) );
oa22f80 g543719 ( .a(n_25693), .b(FE_OFN414_n_28303), .c(n_1353), .d(FE_OFN1143_n_27012), .o(n_26229) );
oa22f80 g543720 ( .a(n_24095), .b(FE_OFN253_n_4280), .c(n_1723), .d(FE_OFN1121_rst), .o(n_24819) );
oa22f80 g543721 ( .a(n_25692), .b(FE_OFN413_n_28303), .c(n_1876), .d(FE_OFN1121_rst), .o(n_26228) );
oa22f80 g543722 ( .a(n_26433), .b(FE_OFN406_n_28303), .c(n_1131), .d(FE_OFN127_n_27449), .o(n_27014) );
oa22f80 g543723 ( .a(n_24094), .b(FE_OFN414_n_28303), .c(n_319), .d(FE_OFN116_n_27449), .o(n_24817) );
oa22f80 g543724 ( .a(n_26153), .b(FE_OFN248_n_4162), .c(n_634), .d(n_29617), .o(n_26774) );
oa22f80 g543725 ( .a(n_25026), .b(FE_OFN406_n_28303), .c(n_795), .d(FE_OFN17_n_29617), .o(n_25727) );
oa22f80 g543726 ( .a(n_25362), .b(FE_OFN405_n_28303), .c(n_632), .d(FE_OFN98_n_27449), .o(n_25971) );
oa22f80 g543727 ( .a(n_23843), .b(FE_OFN413_n_28303), .c(n_773), .d(FE_OFN77_n_27012), .o(n_23884) );
oa22f80 g543728 ( .a(n_25725), .b(FE_OFN268_n_4280), .c(n_1104), .d(FE_OFN1111_rst), .o(n_25726) );
oa22f80 g543729 ( .a(n_25690), .b(FE_OFN417_n_28303), .c(n_36), .d(FE_OFN1124_rst), .o(n_26223) );
oa22f80 g543730 ( .a(n_23818), .b(FE_OFN414_n_28303), .c(n_734), .d(FE_OFN1113_rst), .o(n_24492) );
oa22f80 g543731 ( .a(n_26151), .b(FE_OFN414_n_28303), .c(n_1932), .d(FE_OFN1113_rst), .o(n_26771) );
oa22f80 g543732 ( .a(n_23820), .b(FE_OFN253_n_4280), .c(n_684), .d(FE_OFN78_n_27012), .o(n_24491) );
oa22f80 g543733 ( .a(n_26149), .b(FE_OFN239_n_4162), .c(n_1940), .d(FE_OFN135_n_27449), .o(n_26767) );
oa22f80 g543734 ( .a(n_26148), .b(FE_OFN258_n_4280), .c(n_1824), .d(FE_OFN1121_rst), .o(n_26766) );
oa22f80 g543735 ( .a(n_25360), .b(FE_OFN269_n_4280), .c(n_1095), .d(FE_OFN1114_rst), .o(n_25970) );
oa22f80 g543736 ( .a(n_25361), .b(n_26184), .c(n_1826), .d(FE_OFN90_n_27449), .o(n_25969) );
oa22f80 g543737 ( .a(n_23817), .b(FE_OFN235_n_4162), .c(n_661), .d(n_27449), .o(n_24490) );
oa22f80 g543738 ( .a(n_26145), .b(FE_OFN248_n_4162), .c(n_1092), .d(FE_OFN90_n_27449), .o(n_26765) );
oa22f80 g543739 ( .a(n_25092), .b(FE_OFN244_n_4162), .c(n_1088), .d(FE_OFN108_n_27449), .o(n_25093) );
oa22f80 g543740 ( .a(n_24093), .b(n_4280), .c(n_549), .d(FE_OFN100_n_27449), .o(n_24816) );
oa22f80 g543741 ( .a(n_26427), .b(FE_OFN234_n_4162), .c(n_544), .d(FE_OFN105_n_27449), .o(n_27243) );
oa22f80 g543742 ( .a(n_24092), .b(FE_OFN247_n_4162), .c(n_585), .d(FE_OFN364_n_4860), .o(n_25091) );
oa22f80 g543743 ( .a(n_26425), .b(FE_OFN402_n_28303), .c(n_175), .d(n_28362), .o(n_27242) );
oa22f80 g543744 ( .a(FE_OFN941_n_23815), .b(n_29698), .c(n_1537), .d(FE_OFN1109_rst), .o(n_24815) );
oa22f80 g543745 ( .a(n_25359), .b(FE_OFN410_n_28303), .c(n_1203), .d(FE_OFN76_n_27012), .o(n_26220) );
oa22f80 g543746 ( .a(n_26143), .b(n_28303), .c(n_1583), .d(n_29104), .o(n_27011) );
oa22f80 g543747 ( .a(FE_OFN522_n_25685), .b(FE_OFN411_n_28303), .c(n_1017), .d(n_29104), .o(n_26516) );
oa22f80 g543748 ( .a(n_25909), .b(FE_OFN268_n_4280), .c(n_1052), .d(FE_OFN1111_rst), .o(n_26760) );
oa22f80 g543749 ( .a(n_24365), .b(FE_OFN256_n_4280), .c(n_32), .d(FE_OFN1123_rst), .o(n_25400) );
oa22f80 g543750 ( .a(FE_OFN1230_n_24166), .b(FE_OFN264_n_4280), .c(n_1836), .d(FE_OFN324_n_4860), .o(n_24489) );
ao22s80 g543751 ( .a(n_25363), .b(n_24336), .c(x_out_36_31), .d(n_27400), .o(n_26219) );
in01f80 g543832 ( .a(n_25089), .o(n_25090) );
na02f80 g543833 ( .a(n_24814), .b(n_15183), .o(n_25089) );
no02f80 g543834 ( .a(n_26757), .b(n_26756), .o(n_26758) );
na02f80 g543835 ( .a(n_24488), .b(x_in_2_10), .o(n_25134) );
in01f80 g543836 ( .a(n_24812), .o(n_24813) );
no02f80 g543837 ( .a(n_24488), .b(x_in_2_10), .o(n_24812) );
no02f80 g543838 ( .a(n_24183), .b(n_23882), .o(n_23883) );
no02f80 g543839 ( .a(n_26754), .b(n_26753), .o(n_26755) );
na02f80 g543840 ( .a(n_24811), .b(x_in_34_10), .o(n_25421) );
in01f80 g543841 ( .a(n_25087), .o(n_25088) );
no02f80 g543842 ( .a(n_24811), .b(x_in_34_10), .o(n_25087) );
no02f80 g543843 ( .a(n_26751), .b(n_26750), .o(n_26752) );
no02f80 g543844 ( .a(n_27004), .b(n_27003), .o(n_27005) );
in01f80 g543845 ( .a(n_27238), .o(n_27239) );
na02f80 g543846 ( .a(n_27002), .b(n_26448), .o(n_27238) );
na02f80 g543847 ( .a(n_24810), .b(x_in_18_10), .o(n_25420) );
in01f80 g543848 ( .a(n_25085), .o(n_25086) );
no02f80 g543849 ( .a(n_24810), .b(x_in_18_10), .o(n_25085) );
na02f80 g543850 ( .a(n_24175), .b(x_in_52_10), .o(n_24848) );
no02f80 g543851 ( .a(n_24820), .b(n_24808), .o(n_24809) );
in01f80 g543852 ( .a(n_24846), .o(n_24807) );
no02f80 g543853 ( .a(n_24096), .b(n_24808), .o(n_24846) );
no02f80 g543854 ( .a(n_26748), .b(n_26747), .o(n_26749) );
na02f80 g543855 ( .a(n_24806), .b(x_in_50_10), .o(n_25419) );
in01f80 g543856 ( .a(n_25083), .o(n_25084) );
no02f80 g543857 ( .a(n_24806), .b(x_in_50_10), .o(n_25083) );
na02f80 g543858 ( .a(n_24805), .b(x_in_6_10), .o(n_25418) );
no02f80 g543859 ( .a(n_26745), .b(n_26744), .o(n_26746) );
na02f80 g543860 ( .a(n_24477), .b(x_in_54_11), .o(n_25133) );
in01f80 g543861 ( .a(n_25081), .o(n_25082) );
no02f80 g543862 ( .a(n_24805), .b(x_in_6_10), .o(n_25081) );
na02f80 g543863 ( .a(n_24487), .b(x_in_10_10), .o(n_25132) );
in01f80 g543864 ( .a(n_24803), .o(n_24804) );
no02f80 g543865 ( .a(n_24487), .b(x_in_10_10), .o(n_24803) );
no02f80 g543866 ( .a(n_24188), .b(n_24176), .o(n_24177) );
no02f80 g543867 ( .a(n_26513), .b(n_26512), .o(n_26514) );
in01f80 g543868 ( .a(n_24485), .o(n_24486) );
no02f80 g543869 ( .a(n_24175), .b(x_in_52_10), .o(n_24485) );
na02f80 g543870 ( .a(n_24484), .b(x_in_42_10), .o(n_25131) );
in01f80 g543871 ( .a(n_24801), .o(n_24802) );
no02f80 g543872 ( .a(n_24484), .b(x_in_42_10), .o(n_24801) );
in01f80 g543873 ( .a(n_26213), .o(n_26214) );
na02f80 g543874 ( .a(n_25967), .b(x_in_56_12), .o(n_26213) );
no02f80 g543875 ( .a(n_26510), .b(n_26509), .o(n_26511) );
na02f80 g543876 ( .a(n_24483), .b(x_in_26_10), .o(n_25130) );
in01f80 g543877 ( .a(n_24799), .o(n_24800) );
no02f80 g543878 ( .a(n_24483), .b(x_in_26_10), .o(n_24799) );
na02f80 g543879 ( .a(n_24189), .b(n_24173), .o(n_24174) );
no02f80 g543880 ( .a(n_26211), .b(n_26210), .o(n_26212) );
no02f80 g543881 ( .a(n_26506), .b(n_26505), .o(n_26507) );
na02f80 g543882 ( .a(n_24798), .b(x_in_58_10), .o(n_25417) );
in01f80 g543883 ( .a(n_25079), .o(n_25080) );
no02f80 g543884 ( .a(n_24798), .b(x_in_58_10), .o(n_25079) );
no02f80 g543885 ( .a(n_26741), .b(n_26740), .o(n_26742) );
no02f80 g543886 ( .a(n_26208), .b(n_26466), .o(n_26209) );
no02f80 g543887 ( .a(n_26503), .b(n_26502), .o(n_26504) );
na02f80 g543888 ( .a(n_24797), .b(x_in_6_9), .o(n_25416) );
in01f80 g543889 ( .a(n_25077), .o(n_25078) );
no02f80 g543890 ( .a(n_24797), .b(x_in_6_9), .o(n_25077) );
in01f80 g543891 ( .a(n_25397), .o(n_25398) );
na02f80 g543892 ( .a(n_25076), .b(n_24393), .o(n_25397) );
in01f80 g543893 ( .a(n_25395), .o(n_25396) );
na02f80 g543894 ( .a(n_25075), .b(n_24391), .o(n_25395) );
no02f80 g543895 ( .a(n_26738), .b(n_26737), .o(n_26739) );
na02f80 g543896 ( .a(n_24766), .b(x_in_22_10), .o(n_25415) );
no02f80 g543897 ( .a(n_26499), .b(n_26498), .o(n_26500) );
na02f80 g543898 ( .a(n_24482), .b(x_in_54_10), .o(n_25127) );
in01f80 g543899 ( .a(n_24795), .o(n_24796) );
no02f80 g543900 ( .a(n_24482), .b(x_in_54_10), .o(n_24795) );
no02f80 g543901 ( .a(n_26735), .b(n_26734), .o(n_26736) );
na02f80 g543902 ( .a(n_24481), .b(x_in_2_11), .o(n_25126) );
na02f80 g543903 ( .a(n_24791), .b(x_in_22_11), .o(n_25414) );
no02f80 g543904 ( .a(n_26496), .b(n_26495), .o(n_26497) );
na02f80 g543905 ( .a(n_24794), .b(x_in_40_10), .o(n_25413) );
in01f80 g543906 ( .a(n_25073), .o(n_25074) );
no02f80 g543907 ( .a(n_24794), .b(x_in_40_10), .o(n_25073) );
in01f80 g543908 ( .a(n_24792), .o(n_24793) );
no02f80 g543909 ( .a(n_24481), .b(x_in_2_11), .o(n_24792) );
in01f80 g543910 ( .a(n_25071), .o(n_25072) );
no02f80 g543911 ( .a(n_24791), .b(x_in_22_11), .o(n_25071) );
na02f80 g543912 ( .a(n_24187), .b(n_24171), .o(n_24172) );
no02f80 g543913 ( .a(n_26732), .b(n_26731), .o(n_26733) );
no02f80 g543914 ( .a(n_23583), .b(n_23577), .o(n_23578) );
na02f80 g543915 ( .a(n_24480), .b(x_in_14_10), .o(n_25125) );
in01f80 g543916 ( .a(n_24789), .o(n_24790) );
no02f80 g543917 ( .a(n_24480), .b(x_in_14_10), .o(n_24789) );
no02f80 g543918 ( .a(n_25961), .b(n_25960), .o(n_25962) );
na02f80 g543919 ( .a(n_24479), .b(x_in_46_10), .o(n_25114) );
in01f80 g543920 ( .a(n_24787), .o(n_24788) );
no02f80 g543921 ( .a(n_24479), .b(x_in_46_10), .o(n_24787) );
no02f80 g543922 ( .a(n_26493), .b(n_26492), .o(n_26494) );
na02f80 g543923 ( .a(n_24478), .b(x_in_30_10), .o(n_25124) );
in01f80 g543924 ( .a(n_24785), .o(n_24786) );
no02f80 g543925 ( .a(n_24478), .b(x_in_30_10), .o(n_24785) );
no02f80 g543926 ( .a(n_26490), .b(n_26489), .o(n_26491) );
no02f80 g543927 ( .a(n_26487), .b(n_26486), .o(n_26488) );
na02f80 g543928 ( .a(n_24470), .b(x_in_62_10), .o(n_25123) );
no02f80 g543929 ( .a(n_26729), .b(n_26728), .o(n_26730) );
in01f80 g543930 ( .a(n_24783), .o(n_24784) );
no02f80 g543931 ( .a(n_24477), .b(x_in_54_11), .o(n_24783) );
na02f80 g543932 ( .a(n_23900), .b(n_23880), .o(n_23881) );
na02f80 g543933 ( .a(n_25724), .b(n_246), .o(n_26262) );
na02f80 g543934 ( .a(n_25070), .b(x_in_36_10), .o(n_25738) );
in01f80 g543935 ( .a(n_25393), .o(n_25394) );
no02f80 g543936 ( .a(n_25070), .b(x_in_36_10), .o(n_25393) );
no02f80 g543937 ( .a(n_26206), .b(n_26205), .o(n_26207) );
na02f80 g543938 ( .a(n_24476), .b(x_in_14_11), .o(n_25122) );
in01f80 g543939 ( .a(n_24781), .o(n_24782) );
no02f80 g543940 ( .a(n_24476), .b(x_in_14_11), .o(n_24781) );
na02f80 g543941 ( .a(n_23899), .b(n_23878), .o(n_23879) );
no02f80 g543942 ( .a(n_27234), .b(n_27233), .o(n_27235) );
na02f80 g543943 ( .a(n_24780), .b(x_in_34_11), .o(n_25412) );
in01f80 g543944 ( .a(n_25068), .o(n_25069) );
no02f80 g543945 ( .a(n_24780), .b(x_in_34_11), .o(n_25068) );
no02f80 g543946 ( .a(n_26726), .b(n_26725), .o(n_26727) );
na02f80 g543947 ( .a(n_24475), .b(x_in_46_11), .o(n_25121) );
in01f80 g543948 ( .a(n_24778), .o(n_24779) );
no02f80 g543949 ( .a(n_24475), .b(x_in_46_11), .o(n_24778) );
na02f80 g543950 ( .a(n_23898), .b(n_23876), .o(n_23877) );
no02f80 g543951 ( .a(n_26484), .b(n_26483), .o(n_26485) );
na02f80 g543952 ( .a(n_24474), .b(x_in_16_11), .o(n_25120) );
in01f80 g543953 ( .a(n_24776), .o(n_24777) );
no02f80 g543954 ( .a(n_24474), .b(x_in_16_11), .o(n_24776) );
no02f80 g543955 ( .a(n_23897), .b(n_23874), .o(n_23875) );
no02f80 g543956 ( .a(n_25958), .b(n_25957), .o(n_25959) );
no02f80 g543957 ( .a(n_26723), .b(n_26722), .o(n_26724) );
na02f80 g543958 ( .a(n_24473), .b(x_in_30_11), .o(n_25119) );
in01f80 g543959 ( .a(n_24774), .o(n_24775) );
no02f80 g543960 ( .a(n_24473), .b(x_in_30_11), .o(n_24774) );
na02f80 g543961 ( .a(n_23896), .b(n_23872), .o(n_23873) );
no02f80 g543962 ( .a(n_26481), .b(n_26480), .o(n_26482) );
in01f80 g543963 ( .a(n_24772), .o(n_24773) );
no02f80 g543964 ( .a(n_24472), .b(x_in_18_11), .o(n_24772) );
na02f80 g543965 ( .a(n_24472), .b(x_in_18_11), .o(n_25118) );
no02f80 g543966 ( .a(n_26720), .b(n_26719), .o(n_26721) );
na02f80 g543967 ( .a(n_24471), .b(x_in_62_11), .o(n_25117) );
in01f80 g543968 ( .a(n_24770), .o(n_24771) );
no02f80 g543969 ( .a(n_24471), .b(x_in_62_11), .o(n_24770) );
na02f80 g543970 ( .a(n_23895), .b(n_23870), .o(n_23871) );
no02f80 g543971 ( .a(n_26203), .b(n_26202), .o(n_26204) );
na02f80 g543972 ( .a(n_24767), .b(x_in_12_11), .o(n_25411) );
in01f80 g543973 ( .a(n_24768), .o(n_24769) );
no02f80 g543974 ( .a(n_24470), .b(x_in_62_10), .o(n_24768) );
in01f80 g543975 ( .a(n_25066), .o(n_25067) );
no02f80 g543976 ( .a(n_24767), .b(x_in_12_11), .o(n_25066) );
in01f80 g543977 ( .a(n_25064), .o(n_25065) );
no02f80 g543978 ( .a(n_24766), .b(x_in_22_10), .o(n_25064) );
na02f80 g543979 ( .a(n_24469), .b(x_in_32_9), .o(n_25116) );
in01f80 g543980 ( .a(n_24764), .o(n_24765) );
no02f80 g543981 ( .a(n_24469), .b(x_in_32_9), .o(n_24764) );
na02f80 g543982 ( .a(n_24763), .b(x_in_16_10), .o(n_25410) );
in01f80 g543983 ( .a(n_25062), .o(n_25063) );
no02f80 g543984 ( .a(n_24763), .b(x_in_16_10), .o(n_25062) );
no02f80 g543985 ( .a(n_26200), .b(n_26199), .o(n_26201) );
in01f80 g543986 ( .a(n_25722), .o(n_25723) );
no02f80 g543987 ( .a(n_25392), .b(x_in_48_9), .o(n_25722) );
no02f80 g543988 ( .a(n_26717), .b(n_26716), .o(n_26718) );
na02f80 g543989 ( .a(n_24468), .b(x_in_50_11), .o(n_25115) );
in01f80 g543990 ( .a(n_24761), .o(n_24762) );
no02f80 g543991 ( .a(n_24468), .b(x_in_50_11), .o(n_24761) );
na02f80 g543992 ( .a(n_25392), .b(x_in_48_9), .o(n_25981) );
no02f80 g543993 ( .a(n_23868), .b(n_23867), .o(n_23869) );
na02f80 g543994 ( .a(n_26198), .b(x_in_8_12), .o(n_26837) );
in01f80 g543995 ( .a(n_26478), .o(n_26479) );
no02f80 g543996 ( .a(n_26198), .b(x_in_8_12), .o(n_26478) );
na02f80 g543997 ( .a(n_24467), .b(x_in_32_10), .o(n_25113) );
na02f80 g543998 ( .a(n_25387), .b(x_in_20_10), .o(n_25980) );
na02f80 g543999 ( .a(n_25061), .b(x_in_40_9), .o(n_25737) );
in01f80 g544000 ( .a(n_25390), .o(n_25391) );
no02f80 g544001 ( .a(n_25061), .b(x_in_40_9), .o(n_25390) );
in01f80 g544002 ( .a(n_24759), .o(n_24760) );
no02f80 g544003 ( .a(n_24467), .b(x_in_32_10), .o(n_24759) );
no02f80 g544004 ( .a(n_25955), .b(n_25954), .o(n_25956) );
na02f80 g544005 ( .a(n_25953), .b(x_in_44_13), .o(n_26551) );
in01f80 g544006 ( .a(n_26196), .o(n_26197) );
no02f80 g544007 ( .a(n_25953), .b(x_in_44_13), .o(n_26196) );
no02f80 g544008 ( .a(n_25951), .b(n_25950), .o(n_25952) );
na02f80 g544009 ( .a(n_26195), .b(x_in_56_11), .o(n_26833) );
in01f80 g544010 ( .a(n_26476), .o(n_26477) );
no02f80 g544011 ( .a(n_26195), .b(x_in_56_11), .o(n_26476) );
no02f80 g544012 ( .a(n_26714), .b(n_26713), .o(n_26715) );
na02f80 g544013 ( .a(n_24466), .b(x_in_10_11), .o(n_25112) );
in01f80 g544014 ( .a(n_24757), .o(n_24758) );
no02f80 g544015 ( .a(n_24466), .b(x_in_10_11), .o(n_24757) );
na02f80 g544016 ( .a(n_25060), .b(x_in_48_10), .o(n_25736) );
in01f80 g544017 ( .a(n_25388), .o(n_25389) );
no02f80 g544018 ( .a(n_25060), .b(x_in_48_10), .o(n_25388) );
in01f80 g544019 ( .a(n_25058), .o(n_25059) );
na02f80 g544020 ( .a(n_24756), .b(n_24112), .o(n_25058) );
in01f80 g544021 ( .a(n_25720), .o(n_25721) );
no02f80 g544022 ( .a(n_25387), .b(x_in_20_10), .o(n_25720) );
no02f80 g544023 ( .a(n_24834), .b(n_24754), .o(n_24755) );
no02f80 g544024 ( .a(n_26711), .b(n_26710), .o(n_26712) );
na02f80 g544025 ( .a(n_24465), .b(x_in_42_11), .o(n_25109) );
in01f80 g544026 ( .a(n_25718), .o(n_25719) );
no02f80 g544027 ( .a(n_25386), .b(x_in_36_9), .o(n_25718) );
in01f80 g544028 ( .a(n_24752), .o(n_24753) );
no02f80 g544029 ( .a(n_24465), .b(x_in_42_11), .o(n_24752) );
na02f80 g544030 ( .a(n_25386), .b(x_in_36_9), .o(n_25977) );
no02f80 g544031 ( .a(n_24833), .b(n_24750), .o(n_24751) );
no02f80 g544032 ( .a(n_24493), .b(n_24463), .o(n_24464) );
no02f80 g544033 ( .a(n_23816), .b(n_24463), .o(n_25193) );
no02f80 g544034 ( .a(n_26708), .b(n_26993), .o(n_26709) );
in01f80 g544035 ( .a(n_25948), .o(n_25949) );
no02f80 g544036 ( .a(n_25717), .b(x_in_20_9), .o(n_25948) );
na02f80 g544037 ( .a(n_25717), .b(x_in_20_9), .o(n_26263) );
na02f80 g544038 ( .a(n_25054), .b(x_in_60_10), .o(n_25735) );
no02f80 g544039 ( .a(n_26706), .b(n_26705), .o(n_26707) );
no02f80 g544040 ( .a(n_24496), .b(n_24461), .o(n_24462) );
no02f80 g544041 ( .a(n_23821), .b(n_24461), .o(n_25190) );
na02f80 g544042 ( .a(n_24460), .b(x_in_26_11), .o(n_25108) );
no02f80 g544043 ( .a(n_26995), .b(n_26994), .o(n_26996) );
in01f80 g544044 ( .a(n_24748), .o(n_24749) );
no02f80 g544045 ( .a(n_24460), .b(x_in_26_11), .o(n_24748) );
in01f80 g544046 ( .a(n_24458), .o(n_24459) );
no02f80 g544047 ( .a(n_24170), .b(x_in_52_9), .o(n_24458) );
na02f80 g544048 ( .a(n_24170), .b(x_in_52_9), .o(n_24841) );
no02f80 g544049 ( .a(n_26474), .b(n_26473), .o(n_26475) );
na02f80 g544050 ( .a(n_24747), .b(x_in_12_10), .o(n_25409) );
in01f80 g544051 ( .a(n_25056), .o(n_25057) );
no02f80 g544052 ( .a(n_24747), .b(x_in_12_10), .o(n_25056) );
no02f80 g544053 ( .a(n_25946), .b(n_25945), .o(n_25947) );
na02f80 g544054 ( .a(n_26194), .b(x_in_44_12), .o(n_26832) );
in01f80 g544055 ( .a(n_26471), .o(n_26472) );
no02f80 g544056 ( .a(n_26194), .b(x_in_44_12), .o(n_26471) );
in01f80 g544057 ( .a(n_25384), .o(n_25385) );
na02f80 g544058 ( .a(n_25055), .b(n_24373), .o(n_25384) );
in01f80 g544059 ( .a(n_25382), .o(n_25383) );
no02f80 g544060 ( .a(n_25054), .b(x_in_60_10), .o(n_25382) );
no02f80 g544061 ( .a(n_26469), .b(n_26468), .o(n_26470) );
na02f80 g544062 ( .a(n_24457), .b(x_in_58_11), .o(n_25105) );
na02f80 g544063 ( .a(n_25053), .b(x_in_60_9), .o(n_25739) );
in01f80 g544064 ( .a(n_24745), .o(n_24746) );
no02f80 g544065 ( .a(n_24457), .b(x_in_58_11), .o(n_24745) );
no02f80 g544066 ( .a(n_23901), .b(n_23865), .o(n_23866) );
in01f80 g544067 ( .a(n_25380), .o(n_25381) );
no02f80 g544068 ( .a(n_25053), .b(x_in_60_9), .o(n_25380) );
na02f80 g544069 ( .a(n_24186), .b(n_24168), .o(n_24169) );
no02f80 g544070 ( .a(n_23894), .b(n_23863), .o(n_23864) );
na02f80 g544071 ( .a(FE_OFN1230_n_24166), .b(FE_OFN1106_rst), .o(n_24167) );
no02f80 g544072 ( .a(n_24517), .b(n_24455), .o(n_24456) );
na02f80 g544073 ( .a(n_25706), .b(n_25715), .o(n_25716) );
no02f80 g544074 ( .a(n_24185), .b(n_24163), .o(n_24164) );
na02f80 g544075 ( .a(n_23893), .b(n_23861), .o(n_23862) );
no02f80 g544076 ( .a(n_24832), .b(n_24743), .o(n_24744) );
no02f80 g544077 ( .a(n_23892), .b(n_23859), .o(n_23860) );
no02f80 g544078 ( .a(n_24184), .b(n_24161), .o(n_24162) );
na02f80 g544079 ( .a(n_23582), .b(n_23574), .o(n_23575) );
no02f80 g544080 ( .a(n_24742), .b(FE_OFN411_n_28303), .o(n_25424) );
no02f80 g544081 ( .a(n_24471), .b(n_24454), .o(n_25178) );
na02f80 g544082 ( .a(n_24452), .b(n_24740), .o(n_24453) );
no02f80 g544083 ( .a(n_24791), .b(n_24740), .o(n_25448) );
na02f80 g544084 ( .a(n_24159), .b(n_24451), .o(n_24160) );
no02f80 g544085 ( .a(n_24477), .b(n_24451), .o(n_25181) );
na02f80 g544086 ( .a(n_24157), .b(n_24448), .o(n_24158) );
na02f80 g544087 ( .a(n_24155), .b(n_24449), .o(n_24156) );
na02f80 g544088 ( .a(n_24153), .b(n_24450), .o(n_24154) );
no02f80 g544089 ( .a(n_24473), .b(n_24450), .o(n_25179) );
na02f80 g544090 ( .a(n_24151), .b(n_24454), .o(n_24152) );
no02f80 g544091 ( .a(n_24475), .b(n_24449), .o(n_25183) );
no02f80 g544092 ( .a(n_24476), .b(n_24448), .o(n_25180) );
na02f80 g544093 ( .a(n_24446), .b(n_24739), .o(n_24447) );
no02f80 g544094 ( .a(n_24767), .b(n_24739), .o(n_25443) );
no02f80 g544095 ( .a(n_24512), .b(n_24444), .o(n_24445) );
no02f80 g544096 ( .a(n_23891), .b(n_23857), .o(n_23858) );
no02f80 g544097 ( .a(n_23890), .b(n_23855), .o(n_23856) );
no02f80 g544098 ( .a(n_25402), .b(n_25378), .o(n_25379) );
no02f80 g544099 ( .a(n_24691), .b(n_25378), .o(n_25988) );
na02f80 g544100 ( .a(n_25725), .b(n_25943), .o(n_25714) );
no02f80 g544101 ( .a(n_25953), .b(n_25943), .o(n_25944) );
no02f80 g544102 ( .a(n_23889), .b(n_23853), .o(n_23854) );
no02f80 g544103 ( .a(n_23888), .b(n_23851), .o(n_23852) );
no02f80 g544104 ( .a(n_23887), .b(n_23849), .o(n_23850) );
no02f80 g544105 ( .a(n_23886), .b(n_23847), .o(n_23848) );
no02f80 g544106 ( .a(n_25092), .b(n_25051), .o(n_25052) );
in01f80 g544107 ( .a(n_25049), .o(n_25050) );
no02f80 g544108 ( .a(n_24366), .b(n_25051), .o(n_25049) );
na02f80 g544109 ( .a(n_23902), .b(n_23845), .o(n_23846) );
no02f80 g544110 ( .a(n_24511), .b(n_24442), .o(n_24443) );
na02f80 g544111 ( .a(n_25976), .b(n_25967), .o(n_25942) );
no02f80 g544112 ( .a(n_24149), .b(n_24148), .o(n_24150) );
na02f80 g544113 ( .a(n_23844), .b(n_24148), .o(n_24872) );
no02f80 g544114 ( .a(n_25712), .b(n_25711), .o(n_25713) );
no02f80 g544115 ( .a(n_24440), .b(n_24439), .o(n_24441) );
no02f80 g544116 ( .a(n_25940), .b(n_26193), .o(n_25941) );
no02f80 g544117 ( .a(n_25709), .b(n_25939), .o(n_25710) );
no02f80 g544118 ( .a(n_23581), .b(n_23572), .o(n_23573) );
no02f80 g544119 ( .a(n_24190), .b(n_26312), .o(n_24438) );
no02f80 g544120 ( .a(n_24737), .b(n_24736), .o(n_24738) );
in01f80 g544121 ( .a(n_24735), .o(n_25170) );
na02f80 g544122 ( .a(n_24437), .b(n_24736), .o(n_24735) );
na02f80 g544123 ( .a(n_24435), .b(n_24434), .o(n_24436) );
na02f80 g544124 ( .a(n_24435), .b(n_23735), .o(n_25169) );
na02f80 g544125 ( .a(n_24733), .b(n_24732), .o(n_24734) );
na02f80 g544126 ( .a(n_24733), .b(n_24052), .o(n_25439) );
na02f80 g544127 ( .a(n_24146), .b(n_24433), .o(n_24147) );
in01f80 g544128 ( .a(n_24731), .o(n_25164) );
no02f80 g544129 ( .a(n_24472), .b(n_24433), .o(n_24731) );
na02f80 g544130 ( .a(n_24144), .b(n_24432), .o(n_24145) );
in01f80 g544131 ( .a(n_24730), .o(n_25161) );
no02f80 g544132 ( .a(n_24468), .b(n_24432), .o(n_24730) );
no02f80 g544133 ( .a(FE_OFN923_n_24430), .b(n_24429), .o(n_24431) );
no02f80 g544134 ( .a(FE_OFN923_n_24430), .b(n_23730), .o(n_25753) );
na02f80 g544135 ( .a(n_24427), .b(n_24426), .o(n_24428) );
na02f80 g544136 ( .a(n_24427), .b(n_23729), .o(n_25160) );
na02f80 g544137 ( .a(n_24424), .b(n_24423), .o(n_24425) );
na02f80 g544138 ( .a(n_24424), .b(n_23728), .o(n_25159) );
na02f80 g544139 ( .a(n_24421), .b(n_24420), .o(n_24422) );
na02f80 g544140 ( .a(n_24421), .b(n_23727), .o(n_25158) );
na02f80 g544141 ( .a(n_24142), .b(n_24419), .o(n_24143) );
in01f80 g544142 ( .a(n_24729), .o(n_25155) );
no02f80 g544143 ( .a(n_24457), .b(n_24419), .o(n_24729) );
in01f80 g544144 ( .a(n_26916), .o(n_26704) );
oa12f80 g544145 ( .a(n_24073), .b(n_26466), .c(n_24704), .o(n_26916) );
na02f80 g544146 ( .a(n_24727), .b(n_24726), .o(n_24728) );
na02f80 g544147 ( .a(n_24727), .b(n_24051), .o(n_25434) );
na02f80 g544148 ( .a(n_24417), .b(n_24416), .o(n_24418) );
in01f80 g544149 ( .a(n_26591), .o(n_26465) );
oa12f80 g544150 ( .a(n_23764), .b(n_24383), .c(n_26193), .o(n_26591) );
na02f80 g544151 ( .a(n_24417), .b(n_23725), .o(n_25152) );
no02f80 g544152 ( .a(n_24140), .b(n_24139), .o(n_24141) );
in01f80 g544153 ( .a(n_24137), .o(n_24138) );
na02f80 g544154 ( .a(n_23843), .b(n_24139), .o(n_24137) );
na02f80 g544155 ( .a(n_24135), .b(n_24415), .o(n_24136) );
in01f80 g544156 ( .a(n_24725), .o(n_25149) );
no02f80 g544157 ( .a(n_24474), .b(n_24415), .o(n_24725) );
na02f80 g544158 ( .a(n_24723), .b(n_25048), .o(n_24724) );
in01f80 g544159 ( .a(n_25377), .o(n_25749) );
no02f80 g544160 ( .a(n_25060), .b(n_25048), .o(n_25377) );
no02f80 g544161 ( .a(n_24133), .b(n_24132), .o(n_24134) );
no02f80 g544162 ( .a(n_24133), .b(n_23460), .o(n_25146) );
na02f80 g544163 ( .a(n_24413), .b(n_24722), .o(n_24414) );
in01f80 g544164 ( .a(n_25047), .o(n_25430) );
no02f80 g544165 ( .a(n_24794), .b(n_24722), .o(n_25047) );
no02f80 g544166 ( .a(n_24411), .b(n_24410), .o(n_24412) );
in01f80 g544167 ( .a(n_24409), .o(n_24856) );
na02f80 g544168 ( .a(n_24131), .b(n_24410), .o(n_24409) );
in01f80 g544169 ( .a(n_27298), .o(n_27229) );
oa12f80 g544170 ( .a(n_24681), .b(n_26993), .c(n_25365), .o(n_27298) );
na02f80 g544171 ( .a(n_25070), .b(n_25376), .o(n_25046) );
na02f80 g544172 ( .a(n_24690), .b(n_25376), .o(n_25985) );
na02f80 g544173 ( .a(n_25044), .b(n_25375), .o(n_25045) );
in01f80 g544174 ( .a(n_25708), .o(n_25982) );
no02f80 g544175 ( .a(n_25387), .b(n_25375), .o(n_25708) );
in01f80 g544176 ( .a(n_26284), .o(n_26192) );
oa12f80 g544177 ( .a(n_23504), .b(n_25939), .c(n_24110), .o(n_26284) );
na02f80 g544178 ( .a(n_24129), .b(n_24128), .o(n_24130) );
na02f80 g544179 ( .a(n_24129), .b(n_23459), .o(n_24855) );
no02f80 g544180 ( .a(FE_OFN942_n_24127), .b(n_24406), .o(n_24408) );
in01f80 g544181 ( .a(n_24405), .o(n_24852) );
na02f80 g544182 ( .a(n_24127), .b(n_24406), .o(n_24405) );
na02f80 g544183 ( .a(n_25042), .b(n_25041), .o(n_25043) );
na02f80 g544184 ( .a(n_25042), .b(n_24327), .o(n_25746) );
in01f80 g544185 ( .a(n_27536), .o(n_27428) );
oa12f80 g544186 ( .a(n_24709), .b(n_24084), .c(n_26348), .o(n_27536) );
in01f80 g544187 ( .a(n_27533), .o(n_27427) );
oa12f80 g544188 ( .a(n_25033), .b(n_24359), .c(n_26347), .o(n_27533) );
in01f80 g544189 ( .a(n_27143), .o(n_26992) );
oa12f80 g544190 ( .a(n_24706), .b(n_24081), .c(n_25845), .o(n_27143) );
in01f80 g544191 ( .a(n_27528), .o(n_27425) );
oa12f80 g544192 ( .a(n_24399), .b(n_23802), .c(n_26346), .o(n_27528) );
in01f80 g544193 ( .a(n_27525), .o(n_27424) );
oa12f80 g544194 ( .a(n_24398), .b(n_23797), .c(n_26345), .o(n_27525) );
in01f80 g544195 ( .a(n_27337), .o(n_27228) );
oa12f80 g544196 ( .a(n_24708), .b(n_26065), .c(n_24079), .o(n_27337) );
in01f80 g544197 ( .a(n_27334), .o(n_27227) );
oa12f80 g544198 ( .a(n_24707), .b(n_26064), .c(n_24077), .o(n_27334) );
in01f80 g544199 ( .a(n_27331), .o(n_27226) );
oa12f80 g544200 ( .a(n_24705), .b(n_26063), .c(n_24075), .o(n_27331) );
in01f80 g544201 ( .a(n_27328), .o(n_27225) );
oa12f80 g544202 ( .a(n_24395), .b(n_26062), .c(n_23791), .o(n_27328) );
in01f80 g544203 ( .a(n_26913), .o(n_26703) );
oa12f80 g544204 ( .a(n_24117), .b(n_25564), .c(n_23518), .o(n_26913) );
in01f80 g544205 ( .a(n_27224), .o(n_27656) );
oa12f80 g544206 ( .a(n_23115), .b(n_22454), .c(n_26982), .o(n_27224) );
in01f80 g544207 ( .a(n_26991), .o(n_27471) );
oa12f80 g544208 ( .a(n_23114), .b(n_26691), .c(n_22462), .o(n_26991) );
in01f80 g544209 ( .a(n_27325), .o(n_27223) );
oa12f80 g544210 ( .a(n_24703), .b(n_24068), .c(n_26060), .o(n_27325) );
in01f80 g544211 ( .a(n_27322), .o(n_27222) );
oa12f80 g544212 ( .a(n_24400), .b(n_23782), .c(n_26059), .o(n_27322) );
in01f80 g544213 ( .a(n_27519), .o(n_27421) );
oa12f80 g544214 ( .a(n_24396), .b(n_23786), .c(n_26344), .o(n_27519) );
in01f80 g544215 ( .a(n_27522), .o(n_27420) );
oa12f80 g544216 ( .a(n_24701), .b(n_24064), .c(n_26343), .o(n_27522) );
in01f80 g544217 ( .a(n_26910), .o(n_26701) );
oa12f80 g544218 ( .a(n_24401), .b(n_23780), .c(n_25565), .o(n_26910) );
in01f80 g544219 ( .a(n_27319), .o(n_27221) );
oa12f80 g544220 ( .a(n_24397), .b(n_23778), .c(n_26058), .o(n_27319) );
in01f80 g544221 ( .a(n_27316), .o(n_27220) );
oa12f80 g544222 ( .a(n_24394), .b(n_23776), .c(n_26057), .o(n_27316) );
in01f80 g544223 ( .a(n_27313), .o(n_27219) );
oa12f80 g544224 ( .a(n_24388), .b(n_23774), .c(n_26056), .o(n_27313) );
in01f80 g544225 ( .a(n_27513), .o(n_27417) );
oa12f80 g544226 ( .a(n_24119), .b(n_23534), .c(n_26342), .o(n_27513) );
in01f80 g544227 ( .a(n_26990), .o(n_27469) );
oa12f80 g544228 ( .a(n_22698), .b(n_26689), .c(n_22101), .o(n_26990) );
in01f80 g544229 ( .a(n_27310), .o(n_27218) );
oa12f80 g544230 ( .a(n_25370), .b(n_24688), .c(n_26066), .o(n_27310) );
in01f80 g544231 ( .a(n_27140), .o(n_26989) );
oa12f80 g544232 ( .a(n_24113), .b(n_23530), .c(n_25842), .o(n_27140) );
in01f80 g544233 ( .a(n_27854), .o(n_27799) );
oa12f80 g544234 ( .a(n_24702), .b(n_24066), .c(n_26946), .o(n_27854) );
in01f80 g544235 ( .a(n_27510), .o(n_27414) );
oa12f80 g544236 ( .a(n_24118), .b(n_23528), .c(n_26341), .o(n_27510) );
in01f80 g544237 ( .a(n_27307), .o(n_27217) );
oa12f80 g544238 ( .a(n_24387), .b(n_23770), .c(n_26055), .o(n_27307) );
ao12f80 g544239 ( .a(n_13173), .b(n_24125), .c(n_14356), .o(n_24126) );
in01f80 g544240 ( .a(n_27507), .o(n_27413) );
oa12f80 g544241 ( .a(n_24116), .b(n_23524), .c(n_26340), .o(n_27507) );
in01f80 g544242 ( .a(n_27304), .o(n_27216) );
oa12f80 g544243 ( .a(n_24385), .b(n_23768), .c(n_26054), .o(n_27304) );
in01f80 g544244 ( .a(n_27504), .o(n_27412) );
oa12f80 g544245 ( .a(n_24115), .b(n_23521), .c(n_26339), .o(n_27504) );
in01f80 g544246 ( .a(n_27137), .o(n_26988) );
oa12f80 g544247 ( .a(n_24386), .b(n_23766), .c(n_25841), .o(n_27137) );
oa12f80 g544248 ( .a(n_18838), .b(n_26457), .c(n_18257), .o(n_26839) );
in01f80 g544249 ( .a(n_27134), .o(n_26987) );
oa12f80 g544250 ( .a(n_24379), .b(n_23762), .c(n_25840), .o(n_27134) );
in01f80 g544251 ( .a(n_27500), .o(n_27411) );
oa12f80 g544252 ( .a(n_24384), .b(n_23760), .c(n_26338), .o(n_27500) );
oa12f80 g544253 ( .a(n_2703), .b(n_26188), .c(n_2175), .o(n_26553) );
in01f80 g544254 ( .a(n_26898), .o(n_26700) );
oa12f80 g544255 ( .a(n_24700), .b(n_24061), .c(n_25560), .o(n_26898) );
in01f80 g544256 ( .a(n_26902), .o(n_26699) );
oa12f80 g544257 ( .a(n_24378), .b(n_23755), .c(n_25563), .o(n_26902) );
in01f80 g544258 ( .a(n_27212), .o(n_27654) );
oa12f80 g544259 ( .a(n_23976), .b(n_26980), .c(n_23357), .o(n_27212) );
in01f80 g544260 ( .a(n_26461), .o(n_27079) );
oa12f80 g544261 ( .a(n_22739), .b(n_26186), .c(n_22130), .o(n_26461) );
oa12f80 g544262 ( .a(n_13620), .b(n_24124), .c(n_14265), .o(n_24851) );
in01f80 g544263 ( .a(n_27496), .o(n_27410) );
oa12f80 g544264 ( .a(n_24377), .b(n_26336), .c(n_23753), .o(n_27496) );
in01f80 g544265 ( .a(n_26986), .o(n_27467) );
oa12f80 g544266 ( .a(n_22790), .b(n_22179), .c(n_26686), .o(n_26986) );
in01f80 g544267 ( .a(n_27676), .o(n_27626) );
oa12f80 g544268 ( .a(n_25371), .b(n_24683), .c(n_26623), .o(n_27676) );
in01f80 g544269 ( .a(n_27516), .o(n_27409) );
oa12f80 g544270 ( .a(n_24389), .b(n_23784), .c(n_26337), .o(n_27516) );
in01f80 g544271 ( .a(n_27491), .o(n_27408) );
oa12f80 g544272 ( .a(n_24376), .b(n_26335), .c(n_23751), .o(n_27491) );
in01f80 g544273 ( .a(n_27672), .o(n_27625) );
oa12f80 g544274 ( .a(n_25364), .b(n_24679), .c(n_26622), .o(n_27672) );
in01f80 g544275 ( .a(n_27488), .o(n_27407) );
oa12f80 g544276 ( .a(n_24375), .b(n_26334), .c(n_23747), .o(n_27488) );
in01f80 g544277 ( .a(n_26892), .o(n_26696) );
oa12f80 g544278 ( .a(n_24699), .b(n_24057), .c(n_25562), .o(n_26892) );
in01f80 g544279 ( .a(n_26985), .o(n_27465) );
oa12f80 g544280 ( .a(n_24226), .b(n_26684), .c(n_23641), .o(n_26985) );
in01f80 g544281 ( .a(n_26984), .o(n_27463) );
oa12f80 g544282 ( .a(n_23097), .b(n_26682), .c(n_22439), .o(n_26984) );
in01f80 g544283 ( .a(n_27542), .o(n_27405) );
oa12f80 g544284 ( .a(n_25032), .b(n_24341), .c(n_26333), .o(n_27542) );
in01f80 g544285 ( .a(n_27539), .o(n_27404) );
oa12f80 g544286 ( .a(n_25372), .b(n_24675), .c(n_26332), .o(n_27539) );
in01f80 g544287 ( .a(n_27291), .o(n_27210) );
oa12f80 g544288 ( .a(n_24374), .b(n_26052), .c(n_23744), .o(n_27291) );
oa12f80 g544289 ( .a(n_25706), .b(n_756), .c(FE_OFN99_n_27449), .o(n_25707) );
oa12f80 g544290 ( .a(n_24720), .b(n_800), .c(FE_OFN1106_rst), .o(n_24721) );
ao22s80 g544291 ( .a(n_23458), .b(n_23743), .c(x_out_37_32), .d(n_5003), .o(n_24719) );
no03m80 g544292 ( .a(n_24513), .b(n_24514), .c(n_24515), .o(n_24718) );
in01f80 g544293 ( .a(n_24849), .o(n_24518) );
oa12f80 g544294 ( .a(n_11544), .b(n_23842), .c(n_12267), .o(n_24849) );
oa22f80 g544295 ( .a(n_22579), .b(FE_OFN542_n_23570), .c(n_751), .d(FE_OFN1113_rst), .o(n_23571) );
ao12f80 g544296 ( .a(n_24371), .b(n_24712), .c(n_24370), .o(n_25040) );
in01f80 g544297 ( .a(n_24191), .o(n_24123) );
ao12f80 g544298 ( .a(n_23240), .b(n_23239), .c(n_23238), .o(n_24191) );
ao12f80 g544299 ( .a(n_23828), .b(n_23827), .c(n_23826), .o(n_24404) );
ao22s80 g544300 ( .a(n_23404), .b(n_26982), .c(n_23403), .d(n_26061), .o(n_26983) );
in01f80 g544301 ( .a(n_24527), .o(n_24403) );
oa12f80 g544302 ( .a(n_23564), .b(n_23563), .c(n_23562), .o(n_24527) );
ao12f80 g544303 ( .a(n_10997), .b(n_23167), .c(n_9195), .o(n_24525) );
ao22s80 g544304 ( .a(n_23402), .b(n_26691), .c(n_23401), .d(n_25838), .o(n_26692) );
oa12f80 g544305 ( .a(n_23831), .b(n_23830), .c(n_24105), .o(n_24843) );
ao22s80 g544306 ( .a(n_26689), .b(n_23021), .c(n_25843), .d(n_23020), .o(n_26690) );
ao12f80 g544307 ( .a(n_23834), .b(n_23835), .c(n_23833), .o(n_24837) );
ao12f80 g544308 ( .a(n_25704), .b(n_25703), .c(n_25702), .o(n_26190) );
in01f80 g544309 ( .a(n_24716), .o(n_24717) );
oa12f80 g544310 ( .a(n_23840), .b(n_24125), .c(n_23839), .o(n_24716) );
ao22s80 g544311 ( .a(n_26457), .b(n_19142), .c(n_25561), .d(n_19141), .o(n_26458) );
ao12f80 g544312 ( .a(n_24382), .b(n_24381), .c(n_24380), .o(n_25039) );
ao22s80 g544313 ( .a(n_26188), .b(n_3715), .c(n_25292), .d(n_3714), .o(n_26189) );
ao22s80 g544314 ( .a(n_26980), .b(n_24239), .c(n_26053), .d(n_24238), .o(n_26981) );
oa12f80 g544315 ( .a(n_25927), .b(n_25926), .c(n_26169), .o(n_26836) );
in01f80 g544316 ( .a(n_26555), .o(n_26456) );
oa12f80 g544317 ( .a(n_25701), .b(n_25700), .c(n_25699), .o(n_26555) );
ao22s80 g544318 ( .a(n_26186), .b(n_23069), .c(n_25291), .d(n_23068), .o(n_26187) );
ao12f80 g544319 ( .a(n_24103), .b(n_24102), .c(n_24101), .o(n_24715) );
in01f80 g544320 ( .a(n_24835), .o(n_25102) );
ao12f80 g544321 ( .a(n_23838), .b(n_24124), .c(n_23837), .o(n_24835) );
ao22s80 g544322 ( .a(n_23101), .b(n_26686), .c(n_23100), .d(n_25837), .o(n_26687) );
in01f80 g544323 ( .a(n_24839), .o(n_24842) );
ao12f80 g544324 ( .a(n_23566), .b(n_23842), .c(n_23565), .o(n_24839) );
ao22s80 g544325 ( .a(n_26684), .b(n_24582), .c(n_25836), .d(n_24581), .o(n_26685) );
ao22s80 g544326 ( .a(n_23387), .b(n_26682), .c(n_23386), .d(n_25835), .o(n_26683) );
oa12f80 g544327 ( .a(n_23832), .b(n_23836), .c(n_24106), .o(n_24840) );
oa22f80 g544328 ( .a(n_24043), .b(n_26184), .c(n_1722), .d(FE_OFN1181_rst), .o(n_25038) );
oa22f80 g544329 ( .a(n_23561), .b(FE_OFN1159_n_26184), .c(n_351), .d(FE_OFN1110_rst), .o(n_23841) );
oa22f80 g544330 ( .a(n_25834), .b(FE_OFN162_n_26454), .c(n_1794), .d(FE_OFN347_n_4860), .o(n_26681) );
oa22f80 g544331 ( .a(n_23165), .b(n_26454), .c(n_56), .d(FE_OFN326_n_4860), .o(n_24122) );
oa22f80 g544332 ( .a(n_25558), .b(FE_OFN162_n_26454), .c(n_1803), .d(n_29617), .o(n_26455) );
oa22f80 g544333 ( .a(n_25556), .b(FE_OFN306_n_3069), .c(n_1805), .d(FE_OFN330_n_4860), .o(n_26453) );
oa22f80 g544334 ( .a(n_23717), .b(FE_OFN306_n_3069), .c(n_1724), .d(rst), .o(n_24714) );
oa22f80 g544335 ( .a(n_24712), .b(FE_OFN309_n_3069), .c(n_1819), .d(FE_OFN1181_rst), .o(n_24713) );
oa22f80 g544336 ( .a(n_25289), .b(n_26184), .c(n_655), .d(FE_OFN90_n_27449), .o(n_26185) );
oa22f80 g544337 ( .a(n_24668), .b(FE_OFN208_n_29661), .c(n_1827), .d(FE_OFN114_n_27449), .o(n_25705) );
oa22f80 g544338 ( .a(n_24114), .b(FE_OFN175_n_26184), .c(n_668), .d(FE_OFN352_n_4860), .o(n_24402) );
oa22f80 g544339 ( .a(n_25288), .b(FE_OFN295_n_3069), .c(n_1814), .d(FE_OFN360_n_4860), .o(n_26183) );
oa22f80 g544340 ( .a(n_24042), .b(FE_OFN294_n_3069), .c(n_176), .d(FE_OFN78_n_27012), .o(n_25036) );
oa22f80 g544341 ( .a(n_24989), .b(FE_OFN234_n_4162), .c(n_1967), .d(FE_OFN76_n_27012), .o(n_25934) );
oa22f80 g544342 ( .a(n_24326), .b(FE_OFN307_n_3069), .c(n_1098), .d(FE_OFN1112_rst), .o(n_25374) );
oa22f80 g544343 ( .a(n_23718), .b(n_26454), .c(n_1050), .d(FE_OFN1106_rst), .o(n_24711) );
oa22f80 g544344 ( .a(n_24041), .b(n_26454), .c(n_560), .d(FE_OFN72_n_27012), .o(n_25035) );
oa22f80 g544345 ( .a(n_25832), .b(FE_OFN249_n_4162), .c(n_456), .d(FE_OFN65_n_27012), .o(n_26680) );
oa22f80 g544346 ( .a(n_24987), .b(FE_OFN251_n_4162), .c(n_417), .d(rst), .o(n_25933) );
oa22f80 g544347 ( .a(n_25554), .b(FE_OFN244_n_4162), .c(n_1962), .d(FE_OFN1174_n_4860), .o(n_26451) );
oa22f80 g544348 ( .a(n_25552), .b(FE_OFN249_n_4162), .c(n_752), .d(FE_OFN124_n_27449), .o(n_26450) );
oa22f80 g544349 ( .a(n_25550), .b(FE_OFN256_n_4280), .c(n_609), .d(FE_OFN134_n_27449), .o(n_26449) );
ao22s80 g544350 ( .a(n_24694), .b(n_24693), .c(n_2991), .d(n_6726), .o(n_25034) );
na02f80 g544379 ( .a(n_25372), .b(n_24676), .o(n_26757) );
na02f80 g544380 ( .a(n_24709), .b(n_24085), .o(n_26754) );
na02f80 g544381 ( .a(n_25033), .b(n_24360), .o(n_26751) );
na02f80 g544382 ( .a(n_25371), .b(n_24684), .o(n_27004) );
in01f80 g544383 ( .a(n_26181), .o(n_26182) );
na02f80 g544384 ( .a(n_25932), .b(n_25343), .o(n_26181) );
na02f80 g544385 ( .a(n_26180), .b(x_in_8_13), .o(n_27002) );
in01f80 g544386 ( .a(n_26447), .o(n_26448) );
no02f80 g544387 ( .a(n_26180), .b(x_in_8_13), .o(n_26447) );
na02f80 g544388 ( .a(n_24401), .b(n_23781), .o(n_25961) );
na02f80 g544389 ( .a(n_24400), .b(n_23783), .o(n_26496) );
na02f80 g544390 ( .a(n_24399), .b(n_23803), .o(n_26748) );
na02f80 g544391 ( .a(n_24398), .b(n_23798), .o(n_26745) );
na02f80 g544392 ( .a(n_24708), .b(n_24080), .o(n_26513) );
na02f80 g544393 ( .a(n_24397), .b(n_23779), .o(n_26493) );
na02f80 g544394 ( .a(n_24707), .b(n_24078), .o(n_26510) );
na02f80 g544395 ( .a(n_24706), .b(n_24082), .o(n_26211) );
na02f80 g544396 ( .a(n_24705), .b(n_24076), .o(n_26506) );
na02f80 g544397 ( .a(n_25032), .b(n_24342), .o(n_26741) );
na02f80 g544398 ( .a(n_24396), .b(n_23787), .o(n_26735) );
na02f80 g544399 ( .a(n_24395), .b(n_23792), .o(n_26503) );
na02f80 g544400 ( .a(n_24394), .b(n_23777), .o(n_26487) );
na02f80 g544401 ( .a(n_24121), .b(x_in_38_13), .o(n_25076) );
in01f80 g544402 ( .a(n_24392), .o(n_24393) );
no02f80 g544403 ( .a(n_24121), .b(x_in_38_13), .o(n_24392) );
no02f80 g544404 ( .a(n_24074), .b(n_24704), .o(n_26208) );
na02f80 g544405 ( .a(n_24120), .b(x_in_38_12), .o(n_25075) );
in01f80 g544406 ( .a(n_24390), .o(n_24391) );
no02f80 g544407 ( .a(n_24120), .b(x_in_38_12), .o(n_24390) );
na02f80 g544408 ( .a(n_24389), .b(n_23785), .o(n_26738) );
na02f80 g544409 ( .a(n_24703), .b(n_24069), .o(n_26499) );
na02f80 g544410 ( .a(n_24119), .b(n_23535), .o(n_26729) );
na02f80 g544411 ( .a(n_24388), .b(n_23775), .o(n_26490) );
in01f80 g544412 ( .a(n_26445), .o(n_26446) );
na02f80 g544413 ( .a(n_26179), .b(n_25618), .o(n_26445) );
na02f80 g544414 ( .a(n_24702), .b(n_24067), .o(n_27234) );
na02f80 g544415 ( .a(n_25370), .b(n_24689), .o(n_26474) );
na02f80 g544416 ( .a(n_24118), .b(n_23529), .o(n_26726) );
na02f80 g544417 ( .a(n_24387), .b(n_23771), .o(n_26484) );
na02f80 g544418 ( .a(n_24117), .b(n_23519), .o(n_25958) );
na02f80 g544419 ( .a(n_24386), .b(n_23767), .o(n_26203) );
na02f80 g544420 ( .a(n_24385), .b(n_23769), .o(n_26481) );
na02f80 g544421 ( .a(n_24125), .b(n_23839), .o(n_23840) );
na02f80 g544422 ( .a(n_24116), .b(n_23525), .o(n_26723) );
na02f80 g544423 ( .a(n_24115), .b(n_23522), .o(n_26720) );
na02f80 g544424 ( .a(n_24701), .b(n_24065), .o(n_26732) );
in01f80 g544425 ( .a(n_23568), .o(n_23569) );
na02f80 g544426 ( .a(n_23241), .b(n_22587), .o(n_23568) );
na02f80 g544427 ( .a(n_24384), .b(n_23761), .o(n_26717) );
no02f80 g544428 ( .a(n_23765), .b(n_24383), .o(n_25940) );
no02f80 g544429 ( .a(n_24381), .b(n_24380), .o(n_24382) );
na02f80 g544430 ( .a(n_24114), .b(n_24380), .o(n_24814) );
na02f80 g544431 ( .a(n_24379), .b(n_23763), .o(n_26200) );
in01f80 g544432 ( .a(n_25368), .o(n_25369) );
na02f80 g544433 ( .a(n_25031), .b(n_24355), .o(n_25368) );
in01f80 g544434 ( .a(n_26176), .o(n_26177) );
na02f80 g544435 ( .a(n_25930), .b(n_25307), .o(n_26176) );
na02f80 g544436 ( .a(n_24113), .b(n_23531), .o(n_26206) );
oa22f80 g544437 ( .a(n_22575), .b(n_8910), .c(n_2213), .d(x_in_41_14), .o(n_24166) );
na02f80 g544438 ( .a(n_24700), .b(n_24062), .o(n_25955) );
in01f80 g544439 ( .a(n_26174), .o(n_26175) );
na02f80 g544440 ( .a(n_25929), .b(n_25304), .o(n_26174) );
no02f80 g544441 ( .a(n_24124), .b(n_23837), .o(n_23838) );
na02f80 g544442 ( .a(n_24378), .b(n_23756), .o(n_25951) );
na02f80 g544443 ( .a(n_24377), .b(n_23754), .o(n_26714) );
in01f80 g544444 ( .a(n_26172), .o(n_26173) );
na02f80 g544445 ( .a(n_25928), .b(n_25302), .o(n_26172) );
in01f80 g544446 ( .a(n_25366), .o(n_25367) );
na02f80 g544447 ( .a(n_25030), .b(n_24351), .o(n_25366) );
na02f80 g544448 ( .a(n_24376), .b(n_23752), .o(n_26711) );
na02f80 g544449 ( .a(n_23836), .b(x_in_28_13), .o(n_24756) );
in01f80 g544450 ( .a(n_24111), .o(n_24112) );
no02f80 g544451 ( .a(n_23836), .b(x_in_28_13), .o(n_24111) );
no02f80 g544452 ( .a(n_23842), .b(n_23565), .o(n_23566) );
na02f80 g544453 ( .a(n_24375), .b(n_23748), .o(n_26706) );
no02f80 g544454 ( .a(n_24682), .b(n_25365), .o(n_26708) );
na02f80 g544455 ( .a(n_25364), .b(n_24680), .o(n_26995) );
no02f80 g544456 ( .a(n_23505), .b(n_24110), .o(n_25709) );
na02f80 g544457 ( .a(n_24374), .b(n_23745), .o(n_26469) );
na02f80 g544458 ( .a(n_24699), .b(n_24058), .o(n_25946) );
in01f80 g544459 ( .a(n_26441), .o(n_26442) );
na02f80 g544460 ( .a(n_26171), .b(n_25572), .o(n_26441) );
na02f80 g544461 ( .a(n_24109), .b(x_in_28_12), .o(n_25055) );
in01f80 g544462 ( .a(n_24372), .o(n_24373) );
no02f80 g544463 ( .a(n_24109), .b(x_in_28_12), .o(n_24372) );
na02f80 g544464 ( .a(n_23563), .b(n_23562), .o(n_23564) );
na02f80 g544465 ( .a(n_24335), .b(FE_OFN360_n_4860), .o(n_25715) );
no02f80 g544466 ( .a(n_24104), .b(n_24107), .o(n_24108) );
no02f80 g544467 ( .a(n_23239), .b(n_23238), .o(n_23240) );
no02f80 g544468 ( .a(n_25703), .b(n_25702), .o(n_25704) );
no02f80 g544469 ( .a(n_23835), .b(n_14291), .o(n_24514) );
no02f80 g544470 ( .a(n_23835), .b(n_23833), .o(n_23834) );
na02f80 g544471 ( .a(n_25700), .b(n_25699), .o(n_25701) );
no02f80 g544472 ( .a(n_24712), .b(n_24370), .o(n_24371) );
no02f80 g544473 ( .a(n_23719), .b(n_24370), .o(n_24742) );
no02f80 g544474 ( .a(n_24694), .b(n_24693), .o(n_24695) );
na02f80 g544475 ( .a(n_23836), .b(n_24106), .o(n_23832) );
in01f80 g544476 ( .a(n_24521), .o(n_24369) );
na02f80 g544477 ( .a(n_23457), .b(n_24106), .o(n_24521) );
na02f80 g544478 ( .a(n_25926), .b(n_26169), .o(n_25927) );
no02f80 g544479 ( .a(n_26180), .b(n_26169), .o(n_26831) );
na02f80 g544480 ( .a(n_23830), .b(n_24105), .o(n_23831) );
no02f80 g544481 ( .a(n_24121), .b(n_24105), .o(n_24838) );
in01f80 g544482 ( .a(n_25706), .o(n_25363) );
na02f80 g544483 ( .a(n_25029), .b(FE_OFN146_n_2667), .o(n_25706) );
na02f80 g544484 ( .a(n_24104), .b(FE_OFN1106_rst), .o(n_24720) );
in01f80 g544485 ( .a(n_23829), .o(n_24190) );
na02f80 g544486 ( .a(n_23561), .b(n_23826), .o(n_23829) );
no02f80 g544487 ( .a(n_23827), .b(n_23826), .o(n_23828) );
in01f80 g544488 ( .a(n_23868), .o(n_23560) );
oa12f80 g544489 ( .a(n_13736), .b(n_23237), .c(n_14836), .o(n_23868) );
no02f80 g544490 ( .a(n_24102), .b(n_24101), .o(n_24103) );
no02f80 g544491 ( .a(n_24102), .b(n_23414), .o(n_25101) );
ao12f80 g544492 ( .a(n_14321), .b(n_23236), .c(n_15089), .o(n_23901) );
ao12f80 g544493 ( .a(n_13671), .b(n_23559), .c(n_14791), .o(n_24189) );
in01f80 g544494 ( .a(n_26979), .o(n_27454) );
oa12f80 g544495 ( .a(n_24982), .b(n_24276), .c(n_26673), .o(n_26979) );
oa12f80 g544496 ( .a(n_16678), .b(n_23558), .c(n_16128), .o(n_24188) );
oa12f80 g544497 ( .a(n_15168), .b(n_23557), .c(n_15851), .o(n_24187) );
ao12f80 g544498 ( .a(n_16267), .b(n_22931), .c(n_15564), .o(n_23583) );
oa12f80 g544499 ( .a(n_15163), .b(n_23235), .c(n_15839), .o(n_23900) );
in01f80 g544500 ( .a(n_26440), .o(n_27046) );
oa12f80 g544501 ( .a(n_24981), .b(n_24258), .c(n_26160), .o(n_26440) );
oa12f80 g544502 ( .a(n_15159), .b(n_23234), .c(n_15836), .o(n_23899) );
oa12f80 g544503 ( .a(n_15147), .b(n_23233), .c(n_15829), .o(n_23898) );
ao12f80 g544504 ( .a(n_14731), .b(n_23232), .c(n_15390), .o(n_23897) );
oa12f80 g544505 ( .a(n_15135), .b(n_23231), .c(n_15826), .o(n_23896) );
oa12f80 g544506 ( .a(n_15126), .b(n_23230), .c(n_15823), .o(n_23895) );
in01f80 g544507 ( .a(n_25925), .o(n_26540) );
oa12f80 g544508 ( .a(n_24321), .b(n_23680), .c(n_25691), .o(n_25925) );
in01f80 g544509 ( .a(n_26678), .o(n_27255) );
oa12f80 g544510 ( .a(n_24660), .b(n_23977), .c(n_26432), .o(n_26678) );
ao12f80 g544511 ( .a(n_11829), .b(n_24692), .c(n_13134), .o(n_25406) );
in01f80 g544512 ( .a(n_26439), .o(n_27036) );
oa12f80 g544513 ( .a(n_24657), .b(n_23967), .c(n_26150), .o(n_26439) );
in01f80 g544514 ( .a(n_26438), .o(n_27033) );
oa12f80 g544515 ( .a(n_24028), .b(n_23391), .c(n_26147), .o(n_26438) );
oa12f80 g544516 ( .a(n_15794), .b(n_24100), .c(n_16478), .o(n_24834) );
oa12f80 g544517 ( .a(n_15496), .b(n_24099), .c(n_16249), .o(n_24833) );
ao12f80 g544518 ( .a(n_11438), .b(n_23229), .c(n_12480), .o(n_24183) );
oa12f80 g544519 ( .a(n_22273), .b(n_22881), .c(n_22578), .o(n_23228) );
ao12f80 g544520 ( .a(n_14677), .b(n_23556), .c(n_15360), .o(n_24186) );
ao12f80 g544521 ( .a(n_13969), .b(n_23227), .c(n_14945), .o(n_23894) );
in01f80 g544522 ( .a(n_25724), .o(n_25967) );
ao12f80 g544523 ( .a(n_3642), .b(n_24027), .c(n_8264), .o(n_25724) );
oa12f80 g544524 ( .a(n_16677), .b(n_23825), .c(n_16090), .o(n_24517) );
oa22f80 g544525 ( .a(n_25028), .b(n_23062), .c(n_23346), .d(n_16725), .o(n_25712) );
oa12f80 g544526 ( .a(n_15110), .b(n_23555), .c(n_14298), .o(n_24185) );
oa12f80 g544527 ( .a(n_13647), .b(n_23226), .c(n_14388), .o(n_23893) );
in01f80 g544528 ( .a(n_23824), .o(n_24502) );
ao12f80 g544529 ( .a(n_13680), .b(n_23554), .c(n_14805), .o(n_23824) );
ao12f80 g544530 ( .a(n_13191), .b(n_24098), .c(n_14363), .o(n_24832) );
ao12f80 g544531 ( .a(n_11571), .b(n_23225), .c(n_12509), .o(n_23886) );
oa12f80 g544532 ( .a(n_14490), .b(n_23819), .c(n_13275), .o(n_24511) );
oa12f80 g544533 ( .a(n_13988), .b(n_23224), .c(n_14921), .o(n_23892) );
oa12f80 g544534 ( .a(n_14395), .b(n_23553), .c(n_15150), .o(n_24184) );
oa12f80 g544535 ( .a(n_11444), .b(n_22930), .c(n_12439), .o(n_23582) );
oa12f80 g544536 ( .a(n_14101), .b(n_22929), .c(n_14810), .o(n_23581) );
ao12f80 g544537 ( .a(n_13635), .b(n_23823), .c(n_14669), .o(n_24512) );
ao12f80 g544538 ( .a(n_13917), .b(n_23223), .c(n_14914), .o(n_23891) );
ao12f80 g544539 ( .a(n_13893), .b(n_23222), .c(n_14909), .o(n_23890) );
oa12f80 g544540 ( .a(n_16479), .b(n_23221), .c(n_15801), .o(n_23889) );
ao12f80 g544541 ( .a(n_13873), .b(n_23220), .c(n_14905), .o(n_23888) );
oa12f80 g544542 ( .a(n_13953), .b(n_23219), .c(n_14930), .o(n_23887) );
ao12f80 g544543 ( .a(n_11448), .b(n_23218), .c(n_12441), .o(n_23902) );
ao12f80 g544544 ( .a(n_13678), .b(n_23822), .c(n_14801), .o(n_24440) );
ao12f80 g544545 ( .a(n_23488), .b(n_23487), .c(n_23486), .o(n_24097) );
ao12f80 g544546 ( .a(n_25653), .b(n_25652), .c(n_25651), .o(n_26168) );
oa12f80 g544547 ( .a(n_23187), .b(n_23186), .c(n_23485), .o(n_24488) );
in01f80 g544548 ( .a(n_23821), .o(n_24496) );
oa12f80 g544549 ( .a(n_22927), .b(n_23229), .c(n_22926), .o(n_23821) );
ao12f80 g544550 ( .a(n_25650), .b(n_25649), .c(n_25648), .o(n_26167) );
oa12f80 g544551 ( .a(n_23484), .b(n_23483), .c(n_23734), .o(n_24811) );
ao12f80 g544552 ( .a(n_24334), .b(n_24333), .c(n_24332), .o(n_25027) );
ao12f80 g544553 ( .a(n_25625), .b(n_25624), .c(n_25623), .o(n_26166) );
ao12f80 g544554 ( .a(n_25647), .b(n_25646), .c(n_25645), .o(n_26165) );
ao12f80 g544555 ( .a(n_25346), .b(n_25345), .c(n_25344), .o(n_25924) );
ao12f80 g544556 ( .a(n_25876), .b(n_25875), .c(n_25874), .o(n_26435) );
ao22s80 g544557 ( .a(n_25279), .b(n_26673), .c(n_25278), .d(n_25823), .o(n_26674) );
oa12f80 g544558 ( .a(n_23482), .b(n_23481), .c(n_23480), .o(n_24810) );
in01f80 g544559 ( .a(n_24129), .o(n_24175) );
ao12f80 g544560 ( .a(n_22585), .b(n_22931), .c(n_22584), .o(n_24129) );
ao12f80 g544561 ( .a(n_23801), .b(n_23800), .c(n_23799), .o(n_24368) );
ao12f80 g544562 ( .a(n_25644), .b(n_25643), .c(n_25642), .o(n_26164) );
oa12f80 g544563 ( .a(n_23479), .b(n_23478), .c(n_23477), .o(n_24806) );
ao12f80 g544564 ( .a(n_23733), .b(n_23732), .c(n_23731), .o(n_24367) );
in01f80 g544565 ( .a(n_24727), .o(n_24805) );
ao12f80 g544566 ( .a(n_23217), .b(n_23558), .c(n_23216), .o(n_24727) );
ao12f80 g544567 ( .a(n_25641), .b(n_25640), .c(n_25639), .o(n_26163) );
oa12f80 g544568 ( .a(n_23185), .b(n_23184), .c(n_23475), .o(n_24487) );
ao12f80 g544569 ( .a(n_25341), .b(n_25340), .c(n_25339), .o(n_25923) );
oa12f80 g544570 ( .a(n_23183), .b(n_23182), .c(n_23474), .o(n_24484) );
ao12f80 g544571 ( .a(n_25338), .b(n_25337), .c(n_25336), .o(n_25922) );
oa12f80 g544572 ( .a(n_23181), .b(n_23180), .c(n_23473), .o(n_24483) );
in01f80 g544573 ( .a(n_24437), .o(n_24737) );
ao12f80 g544574 ( .a(n_23215), .b(n_23559), .c(n_23214), .o(n_24437) );
ao12f80 g544575 ( .a(n_25335), .b(n_25334), .c(n_25566), .o(n_25921) );
ao12f80 g544576 ( .a(n_25333), .b(n_25332), .c(n_25331), .o(n_25920) );
oa12f80 g544577 ( .a(n_23472), .b(n_23471), .c(n_23470), .o(n_24798) );
ao12f80 g544578 ( .a(n_25638), .b(n_25637), .c(n_25636), .o(n_26162) );
ao12f80 g544579 ( .a(n_25020), .b(n_25019), .c(n_25297), .o(n_25698) );
ao12f80 g544580 ( .a(n_25349), .b(n_25348), .c(n_25347), .o(n_25919) );
oa12f80 g544581 ( .a(n_23469), .b(n_23468), .c(n_23726), .o(n_24797) );
ao12f80 g544582 ( .a(n_25330), .b(n_25329), .c(n_25559), .o(n_25918) );
oa12f80 g544583 ( .a(n_23500), .b(n_23540), .c(n_23740), .o(n_24766) );
oa12f80 g544584 ( .a(n_23195), .b(n_23211), .c(n_23499), .o(n_24482) );
in01f80 g544585 ( .a(n_24435), .o(n_24481) );
ao12f80 g544586 ( .a(n_22904), .b(n_23224), .c(n_22903), .o(n_24435) );
ao12f80 g544587 ( .a(n_25328), .b(n_25327), .c(n_25326), .o(n_25917) );
in01f80 g544588 ( .a(n_24452), .o(n_24791) );
ao12f80 g544589 ( .a(n_23213), .b(n_23557), .c(n_23212), .o(n_24452) );
oa12f80 g544590 ( .a(n_23194), .b(n_23210), .c(n_23498), .o(n_24480) );
oa12f80 g544591 ( .a(n_23192), .b(n_23209), .c(n_23497), .o(n_24479) );
ao12f80 g544592 ( .a(n_25319), .b(n_25318), .c(n_25317), .o(n_25916) );
oa12f80 g544593 ( .a(n_23196), .b(n_23208), .c(n_23495), .o(n_24478) );
ao12f80 g544594 ( .a(n_25316), .b(n_25315), .c(n_25314), .o(n_25915) );
oa12f80 g544595 ( .a(n_23193), .b(n_23207), .c(n_23496), .o(n_24470) );
in01f80 g544596 ( .a(n_24159), .o(n_24477) );
ao12f80 g544597 ( .a(n_22925), .b(n_23235), .c(n_22924), .o(n_24159) );
ao12f80 g544598 ( .a(n_25322), .b(n_25321), .c(n_25320), .o(n_25914) );
ao22s80 g544599 ( .a(n_25277), .b(n_26160), .c(n_25276), .d(n_25273), .o(n_26161) );
ao12f80 g544600 ( .a(n_25616), .b(n_25615), .c(n_25614), .o(n_26159) );
ao12f80 g544601 ( .a(n_25611), .b(n_25610), .c(n_25609), .o(n_26158) );
ao12f80 g544602 ( .a(n_25568), .b(n_25567), .c(n_25844), .o(n_26157) );
in01f80 g544603 ( .a(n_24157), .o(n_24476) );
ao12f80 g544604 ( .a(n_22923), .b(n_23234), .c(n_22922), .o(n_24157) );
ao12f80 g544605 ( .a(n_25018), .b(n_25017), .c(n_25016), .o(n_25697) );
in01f80 g544606 ( .a(n_24733), .o(n_24780) );
ao12f80 g544607 ( .a(n_23198), .b(n_23553), .c(n_23197), .o(n_24733) );
in01f80 g544608 ( .a(n_24155), .o(n_24475) );
ao12f80 g544609 ( .a(n_22921), .b(n_23233), .c(n_22920), .o(n_24155) );
ao12f80 g544611 ( .a(n_22906), .b(n_23226), .c(n_22905), .o(n_24127) );
ao12f80 g544612 ( .a(n_25599), .b(n_25598), .c(n_25597), .o(n_26156) );
in01f80 g544613 ( .a(n_24135), .o(n_24474) );
ao12f80 g544614 ( .a(n_22919), .b(n_23232), .c(n_22918), .o(n_24135) );
ao12f80 g544615 ( .a(n_25015), .b(n_25014), .c(FE_OFN1252_n_25296), .o(n_25696) );
in01f80 g544616 ( .a(n_24691), .o(n_25402) );
oa12f80 g544617 ( .a(n_23742), .b(n_24098), .c(n_23741), .o(n_24691) );
ao12f80 g544618 ( .a(n_26097), .b(n_26096), .c(n_26095), .o(n_26671) );
ao12f80 g544619 ( .a(n_25313), .b(n_25312), .c(n_25311), .o(n_25913) );
in01f80 g544620 ( .a(n_24153), .o(n_24473) );
ao12f80 g544621 ( .a(n_22917), .b(n_23231), .c(n_22916), .o(n_24153) );
in01f80 g544622 ( .a(n_24146), .o(n_24472) );
ao12f80 g544623 ( .a(n_22908), .b(n_23227), .c(n_22907), .o(n_24146) );
ao12f80 g544624 ( .a(n_25596), .b(n_25595), .c(n_25594), .o(n_26155) );
in01f80 g544625 ( .a(n_24151), .o(n_24471) );
ao12f80 g544626 ( .a(n_22915), .b(n_23230), .c(n_22914), .o(n_24151) );
in01f80 g544627 ( .a(n_24446), .o(n_24767) );
ao12f80 g544628 ( .a(n_23202), .b(n_23556), .c(n_23201), .o(n_24446) );
ao12f80 g544629 ( .a(n_25593), .b(n_25592), .c(n_25591), .o(n_26154) );
in01f80 g544630 ( .a(n_24096), .o(n_24820) );
oa12f80 g544631 ( .a(n_23191), .b(n_23554), .c(n_23190), .o(n_24096) );
oa12f80 g544632 ( .a(n_23179), .b(n_23178), .c(n_23467), .o(n_24469) );
ao12f80 g544633 ( .a(n_25310), .b(n_25309), .c(n_25308), .o(n_25912) );
ao12f80 g544634 ( .a(n_22888), .b(n_22887), .c(n_22886), .o(n_23552) );
ao12f80 g544635 ( .a(n_25013), .b(n_25012), .c(n_25290), .o(n_25695) );
oa12f80 g544636 ( .a(n_23466), .b(n_23465), .c(n_23464), .o(n_24763) );
oa12f80 g544637 ( .a(n_22274), .b(FE_OFN542_n_23570), .c(x_in_12_15), .o(n_29140) );
ao12f80 g544638 ( .a(n_25011), .b(n_25010), .c(n_25009), .o(n_25694) );
oa12f80 g544639 ( .a(n_24050), .b(n_24049), .c(n_24048), .o(n_25392) );
in01f80 g544640 ( .a(n_24144), .o(n_24468) );
ao12f80 g544641 ( .a(n_22894), .b(n_23219), .c(n_22893), .o(n_24144) );
oa22f80 g544642 ( .a(n_21979), .b(FE_OFN269_n_4280), .c(n_689), .d(FE_OFN116_n_27449), .o(n_22928) );
in01f80 g544643 ( .a(n_24723), .o(n_25060) );
ao12f80 g544644 ( .a(n_23493), .b(n_23823), .c(n_23492), .o(n_24723) );
ao12f80 g544645 ( .a(n_25008), .b(n_25007), .c(n_25006), .o(n_25693) );
ao12f80 g544646 ( .a(n_23463), .b(n_23462), .c(n_23461), .o(n_24095) );
in01f80 g544647 ( .a(n_24133), .o(n_23820) );
oa12f80 g544648 ( .a(n_22890), .b(n_23237), .c(n_22889), .o(n_24133) );
ao22s80 g544649 ( .a(n_24662), .b(n_25691), .c(n_24661), .d(n_24647), .o(n_25692) );
ao22s80 g544650 ( .a(n_24980), .b(n_26432), .c(n_24979), .d(n_25543), .o(n_26433) );
in01f80 g544651 ( .a(FE_OFN923_n_24430), .o(n_24094) );
oa22f80 g544652 ( .a(n_22868), .b(n_14818), .c(n_23819), .d(n_14819), .o(n_24430) );
oa12f80 g544653 ( .a(n_24995), .b(n_25021), .c(n_25298), .o(n_26198) );
ao12f80 g544654 ( .a(n_25587), .b(n_25586), .c(n_25585), .o(n_26153) );
in01f80 g544655 ( .a(n_24417), .o(n_24467) );
ao12f80 g544656 ( .a(n_22898), .b(n_23221), .c(n_22897), .o(n_24417) );
ao12f80 g544657 ( .a(n_24339), .b(n_24338), .c(n_24337), .o(n_25026) );
in01f80 g544658 ( .a(n_25044), .o(n_25387) );
ao12f80 g544659 ( .a(n_23759), .b(n_24100), .c(n_23758), .o(n_25044) );
oa12f80 g544660 ( .a(n_23724), .b(n_23723), .c(n_23722), .o(n_25061) );
in01f80 g544661 ( .a(n_24413), .o(n_24794) );
ao12f80 g544662 ( .a(n_23200), .b(n_23555), .c(n_23199), .o(n_24413) );
ao12f80 g544663 ( .a(n_24687), .b(n_24686), .c(n_24685), .o(n_25362) );
in01f80 g544664 ( .a(n_25725), .o(n_25953) );
ao12f80 g544665 ( .a(n_24353), .b(n_24692), .c(n_24352), .o(n_25725) );
ao12f80 g544666 ( .a(n_25325), .b(n_25324), .c(n_25323), .o(n_25911) );
in01f80 g544667 ( .a(n_23843), .o(n_24140) );
ao12f80 g544668 ( .a(n_22583), .b(n_22929), .c(n_22582), .o(n_23843) );
ao12f80 g544669 ( .a(n_25003), .b(n_25002), .c(n_25295), .o(n_25690) );
ao12f80 g544670 ( .a(n_25590), .b(n_25589), .c(n_25588), .o(n_26152) );
oa12f80 g544671 ( .a(n_24994), .b(n_24993), .c(n_25294), .o(n_26195) );
in01f80 g544672 ( .a(n_24427), .o(n_24466) );
ao12f80 g544673 ( .a(n_22902), .b(n_23223), .c(n_22901), .o(n_24427) );
ao12f80 g544674 ( .a(n_23176), .b(n_23175), .c(n_23174), .o(n_23818) );
in01f80 g544675 ( .a(n_24131), .o(n_24411) );
ao12f80 g544676 ( .a(n_22892), .b(n_23218), .c(n_22891), .o(n_24131) );
ao22s80 g544677 ( .a(n_24973), .b(n_26150), .c(n_24972), .d(n_25272), .o(n_26151) );
ao12f80 g544678 ( .a(n_25583), .b(n_25582), .c(n_25581), .o(n_26149) );
ao22s80 g544679 ( .a(n_24318), .b(n_26147), .c(n_24317), .d(n_25271), .o(n_26148) );
ao12f80 g544680 ( .a(n_24671), .b(n_24670), .c(n_24669), .o(n_25361) );
ao12f80 g544681 ( .a(n_24674), .b(n_25028), .c(n_24673), .o(n_25360) );
ao12f80 g544682 ( .a(n_23189), .b(n_23548), .c(n_23188), .o(n_23817) );
in01f80 g544683 ( .a(n_23844), .o(n_24149) );
ao12f80 g544684 ( .a(n_22581), .b(n_22930), .c(n_22580), .o(n_23844) );
in01f80 g544685 ( .a(n_24424), .o(n_24465) );
ao12f80 g544686 ( .a(n_22900), .b(n_23222), .c(n_22899), .o(n_24424) );
oa12f80 g544687 ( .a(n_24047), .b(n_24046), .c(n_24331), .o(n_25386) );
in01f80 g544688 ( .a(n_25070), .o(n_24690) );
oa12f80 g544689 ( .a(n_23750), .b(n_24099), .c(n_23749), .o(n_25070) );
ao12f80 g544690 ( .a(n_25580), .b(n_25579), .c(n_25578), .o(n_26145) );
in01f80 g544691 ( .a(n_24366), .o(n_25092) );
oa12f80 g544692 ( .a(n_23490), .b(n_23822), .c(n_23489), .o(n_24366) );
ao12f80 g544693 ( .a(n_23512), .b(n_23511), .c(n_23510), .o(n_24093) );
in01f80 g544694 ( .a(n_23816), .o(n_24493) );
oa12f80 g544695 ( .a(n_22912), .b(n_23225), .c(n_22911), .o(n_23816) );
ao12f80 g544696 ( .a(n_25853), .b(n_25852), .c(n_26050), .o(n_26427) );
oa12f80 g544697 ( .a(n_24330), .b(n_24329), .c(n_24328), .o(n_25717) );
in01f80 g544698 ( .a(n_25042), .o(n_25054) );
ao12f80 g544699 ( .a(n_23502), .b(n_23825), .c(n_23501), .o(n_25042) );
ao12f80 g544700 ( .a(n_23508), .b(n_23507), .c(n_23506), .o(n_24092) );
in01f80 g544701 ( .a(n_24421), .o(n_24460) );
ao12f80 g544702 ( .a(n_22896), .b(n_23220), .c(n_22895), .o(n_24421) );
ao12f80 g544703 ( .a(n_25851), .b(n_25850), .c(n_25849), .o(n_26425) );
oa12f80 g544704 ( .a(n_22884), .b(n_22883), .c(n_23173), .o(n_24170) );
ao12f80 g544705 ( .a(n_23172), .b(n_23171), .c(n_23170), .o(n_23815) );
ao12f80 g544706 ( .a(n_24678), .b(n_24677), .c(n_24991), .o(n_25359) );
oa12f80 g544707 ( .a(n_23494), .b(n_23526), .c(n_23739), .o(n_24747) );
ao12f80 g544708 ( .a(n_25577), .b(n_25576), .c(n_25575), .o(n_26143) );
ao12f80 g544709 ( .a(n_25000), .b(n_24999), .c(n_25293), .o(n_25685) );
in01f80 g544710 ( .a(n_26194), .o(n_25909) );
oa12f80 g544711 ( .a(n_24998), .b(n_24997), .c(n_25004), .o(n_26194) );
ao12f80 g544712 ( .a(n_23738), .b(n_23737), .c(n_23736), .o(n_24365) );
in01f80 g544713 ( .a(n_24142), .o(n_24457) );
ao12f80 g544714 ( .a(n_22910), .b(n_23236), .c(n_22909), .o(n_24142) );
oa12f80 g544715 ( .a(n_23721), .b(n_23720), .c(n_24045), .o(n_25053) );
oa22f80 g544716 ( .a(n_23413), .b(FE_OFN268_n_4280), .c(n_1464), .d(FE_OFN119_n_27449), .o(n_24364) );
oa22f80 g544717 ( .a(n_24971), .b(FE_OFN268_n_4280), .c(n_19), .d(FE_OFN72_n_27012), .o(n_25908) );
oa22f80 g544718 ( .a(n_23204), .b(FE_OFN402_n_28303), .c(n_255), .d(FE_OFN128_n_27449), .o(n_23551) );
oa22f80 g544719 ( .a(n_24970), .b(FE_OFN265_n_4280), .c(n_1838), .d(FE_OFN128_n_27449), .o(n_25907) );
oa22f80 g544720 ( .a(n_24951), .b(FE_OFN230_n_4162), .c(n_29), .d(n_29261), .o(n_25904) );
oa22f80 g544721 ( .a(FE_OFN742_n_24025), .b(FE_OFN257_n_4280), .c(n_358), .d(n_29261), .o(n_25025) );
oa22f80 g544722 ( .a(n_25270), .b(n_29691), .c(n_1694), .d(FE_OFN1108_rst), .o(n_26141) );
oa22f80 g544723 ( .a(n_24646), .b(FE_OFN267_n_4280), .c(n_671), .d(FE_OFN1110_rst), .o(n_25684) );
oa22f80 g544724 ( .a(n_24969), .b(FE_OFN1157_n_26184), .c(n_1861), .d(FE_OFN1124_rst), .o(n_25902) );
oa22f80 g544725 ( .a(n_25540), .b(FE_OFN175_n_26184), .c(n_983), .d(FE_OFN127_n_27449), .o(n_26415) );
oa22f80 g544726 ( .a(n_23412), .b(FE_OFN149_n_25677), .c(n_188), .d(FE_OFN1174_n_4860), .o(n_24363) );
oa22f80 g544727 ( .a(n_24968), .b(FE_OFN244_n_4162), .c(n_1516), .d(FE_OFN361_n_4860), .o(n_25900) );
oa22f80 g544728 ( .a(n_23144), .b(n_4162), .c(n_1198), .d(FE_OFN353_n_4860), .o(n_24091) );
oa22f80 g544729 ( .a(FE_OFN905_n_24967), .b(n_21988), .c(n_736), .d(FE_OFN56_n_27012), .o(n_25899) );
oa22f80 g544730 ( .a(n_24645), .b(FE_OFN295_n_3069), .c(n_505), .d(FE_OFN15_n_29068), .o(n_25682) );
oa22f80 g544731 ( .a(FE_OFN821_n_24644), .b(n_21988), .c(n_278), .d(n_25680), .o(n_25681) );
oa22f80 g544732 ( .a(n_23143), .b(FE_OFN268_n_4280), .c(n_161), .d(FE_OFN65_n_27012), .o(n_24090) );
oa22f80 g544733 ( .a(n_24965), .b(FE_OFN257_n_4280), .c(n_1047), .d(FE_OFN63_n_27012), .o(n_25898) );
oa22f80 g544734 ( .a(n_24964), .b(FE_OFN251_n_4162), .c(n_1669), .d(FE_OFN65_n_27012), .o(n_25897) );
oa22f80 g544735 ( .a(n_24643), .b(n_21988), .c(n_1532), .d(FE_OFN1172_n_4860), .o(n_25679) );
oa22f80 g544736 ( .a(n_24642), .b(FE_OFN148_n_25677), .c(n_39), .d(FE_OFN329_n_4860), .o(n_25678) );
oa22f80 g544737 ( .a(n_24641), .b(FE_OFN150_n_25677), .c(n_257), .d(n_27709), .o(n_25676) );
oa22f80 g544738 ( .a(n_24639), .b(FE_OFN253_n_4280), .c(n_1236), .d(FE_OFN1119_rst), .o(n_25675) );
oa22f80 g544739 ( .a(n_24638), .b(n_21988), .c(n_1739), .d(FE_OFN1117_rst), .o(n_25673) );
oa22f80 g544740 ( .a(FE_OFN809_n_24927), .b(n_21988), .c(n_208), .d(n_27449), .o(n_25896) );
oa22f80 g544741 ( .a(n_24957), .b(FE_OFN240_n_4162), .c(n_1645), .d(FE_OFN1119_rst), .o(n_25894) );
oa22f80 g544742 ( .a(n_24637), .b(FE_OFN148_n_25677), .c(n_1691), .d(FE_OFN125_n_27449), .o(n_25672) );
oa22f80 g544743 ( .a(n_24636), .b(FE_OFN148_n_25677), .c(n_1051), .d(FE_OFN98_n_27449), .o(n_25671) );
oa22f80 g544744 ( .a(n_24635), .b(FE_OFN150_n_25677), .c(n_1269), .d(FE_OFN129_n_27449), .o(n_25670) );
oa22f80 g544745 ( .a(n_24634), .b(n_21988), .c(n_1529), .d(FE_OFN75_n_27012), .o(n_25669) );
oa22f80 g544746 ( .a(n_22857), .b(n_23813), .c(n_1820), .d(FE_OFN335_n_4860), .o(n_23814) );
oa22f80 g544747 ( .a(FE_OFN1007_n_24950), .b(n_21988), .c(n_1270), .d(FE_OFN56_n_27012), .o(n_25893) );
oa22f80 g544748 ( .a(FE_OFN446_n_24948), .b(n_26184), .c(n_1286), .d(FE_OFN190_n_28362), .o(n_25892) );
oa22f80 g544749 ( .a(n_23548), .b(n_26184), .c(n_348), .d(FE_OFN190_n_28362), .o(n_23549) );
oa22f80 g544750 ( .a(n_23205), .b(FE_OFN160_n_28014), .c(n_603), .d(FE_OFN360_n_4860), .o(n_23547) );
oa22f80 g544751 ( .a(n_25265), .b(FE_OFN156_n_28014), .c(n_1192), .d(FE_OFN286_n_29266), .o(n_26134) );
oa22f80 g544752 ( .a(n_24633), .b(FE_OFN156_n_28014), .c(n_511), .d(FE_OFN288_n_29266), .o(n_25668) );
oa22f80 g544753 ( .a(n_22862), .b(FE_OFN160_n_28014), .c(n_1381), .d(FE_OFN1120_rst), .o(n_23812) );
oa22f80 g544754 ( .a(n_24946), .b(n_23813), .c(n_1531), .d(FE_OFN357_n_4860), .o(n_25889) );
oa22f80 g544755 ( .a(n_24632), .b(FE_OFN259_n_4280), .c(n_1886), .d(FE_OFN360_n_4860), .o(n_25667) );
oa22f80 g544756 ( .a(n_24053), .b(FE_OFN254_n_4280), .c(n_762), .d(FE_OFN131_n_27449), .o(n_24362) );
oa22f80 g544757 ( .a(n_25538), .b(FE_OFN313_n_3069), .c(n_1211), .d(FE_OFN1124_rst), .o(n_26397) );
oa22f80 g544758 ( .a(n_24631), .b(FE_OFN294_n_3069), .c(n_895), .d(FE_OFN133_n_27449), .o(n_25666) );
oa22f80 g544759 ( .a(n_24945), .b(FE_OFN157_n_28014), .c(n_1254), .d(FE_OFN114_n_27449), .o(n_25888) );
oa22f80 g544760 ( .a(n_24944), .b(FE_OFN156_n_28014), .c(n_755), .d(FE_OFN357_n_4860), .o(n_25887) );
oa22f80 g544761 ( .a(n_23543), .b(FE_OFN157_n_28014), .c(n_1752), .d(FE_OFN134_n_27449), .o(n_23811) );
oa22f80 g544762 ( .a(n_24630), .b(FE_OFN244_n_4162), .c(n_1894), .d(FE_OFN361_n_4860), .o(n_25664) );
oa22f80 g544763 ( .a(n_22859), .b(FE_OFN258_n_4280), .c(n_1882), .d(FE_OFN104_n_27449), .o(n_23810) );
oa22f80 g544764 ( .a(n_24315), .b(FE_OFN254_n_4280), .c(n_1840), .d(FE_OFN142_n_27449), .o(n_25355) );
oa22f80 g544765 ( .a(n_24314), .b(FE_OFN299_n_3069), .c(n_1493), .d(FE_OFN133_n_27449), .o(n_25353) );
oa22f80 g544766 ( .a(n_24629), .b(FE_OFN265_n_4280), .c(n_1112), .d(FE_OFN1143_n_27012), .o(n_25663) );
oa22f80 g544767 ( .a(n_22858), .b(FE_OFN297_n_3069), .c(n_1094), .d(FE_OFN138_n_27449), .o(n_23809) );
oa22f80 g544768 ( .a(n_24313), .b(FE_OFN413_n_28303), .c(n_747), .d(FE_OFN104_n_27449), .o(n_25351) );
oa22f80 g544769 ( .a(n_23476), .b(FE_OFN414_n_28303), .c(n_1014), .d(FE_OFN116_n_27449), .o(n_23808) );
oa22f80 g544770 ( .a(n_24940), .b(FE_OFN235_n_4162), .c(n_1685), .d(FE_OFN335_n_4860), .o(n_25886) );
oa22f80 g544771 ( .a(n_25261), .b(FE_OFN406_n_28303), .c(n_897), .d(FE_OFN360_n_4860), .o(n_26127) );
oa22f80 g544772 ( .a(n_24024), .b(FE_OFN249_n_4162), .c(n_45), .d(FE_OFN330_n_4860), .o(n_25024) );
oa22f80 g544773 ( .a(n_22556), .b(FE_OFN240_n_4162), .c(n_1324), .d(FE_OFN104_n_27449), .o(n_23546) );
oa22f80 g544774 ( .a(n_24672), .b(FE_OFN248_n_4162), .c(n_100), .d(FE_OFN113_n_27449), .o(n_25023) );
oa22f80 g544775 ( .a(n_24626), .b(FE_OFN254_n_4280), .c(n_878), .d(FE_OFN142_n_27449), .o(n_25658) );
oa22f80 g544776 ( .a(n_23140), .b(FE_OFN269_n_4280), .c(n_1504), .d(FE_OFN1143_n_27012), .o(n_24089) );
oa22f80 g544777 ( .a(n_24933), .b(n_4162), .c(n_41), .d(FE_OFN1143_n_27012), .o(n_25884) );
oa22f80 g544778 ( .a(n_23177), .b(FE_OFN297_n_3069), .c(n_1221), .d(FE_OFN78_n_27012), .o(n_23545) );
oa22f80 g544779 ( .a(n_24930), .b(FE_OFN239_n_4162), .c(n_166), .d(FE_OFN135_n_27449), .o(n_25883) );
oa22f80 g544780 ( .a(n_24929), .b(FE_OFN258_n_4280), .c(n_667), .d(FE_OFN77_n_27012), .o(n_25881) );
oa22f80 g544781 ( .a(n_22856), .b(FE_OFN266_n_4280), .c(n_1488), .d(FE_OFN60_n_27012), .o(n_23807) );
oa22f80 g544782 ( .a(n_23491), .b(FE_OFN416_n_28303), .c(n_126), .d(FE_OFN108_n_27449), .o(n_23806) );
oa22f80 g544783 ( .a(n_24926), .b(FE_OFN248_n_4162), .c(n_11), .d(FE_OFN90_n_27449), .o(n_25880) );
oa22f80 g544784 ( .a(n_23139), .b(FE_OFN406_n_28303), .c(n_786), .d(FE_OFN360_n_4860), .o(n_24088) );
oa22f80 g544785 ( .a(n_25259), .b(FE_OFN404_n_28303), .c(n_389), .d(FE_OFN357_n_4860), .o(n_26122) );
oa22f80 g544786 ( .a(n_23138), .b(FE_OFN309_n_3069), .c(n_1760), .d(FE_OFN69_n_27012), .o(n_24087) );
oa22f80 g544787 ( .a(n_25258), .b(FE_OFN247_n_4162), .c(n_33), .d(FE_OFN1174_n_4860), .o(n_26121) );
oa22f80 g544788 ( .a(n_23137), .b(FE_OFN239_n_4162), .c(n_1100), .d(FE_OFN135_n_27449), .o(n_24086) );
oa22f80 g544789 ( .a(n_24023), .b(FE_OFN259_n_4280), .c(n_733), .d(FE_OFN130_n_27449), .o(n_25022) );
oa22f80 g544790 ( .a(n_24925), .b(n_4280), .c(n_1822), .d(FE_OFN105_n_27449), .o(n_25879) );
oa22f80 g544791 ( .a(n_24625), .b(FE_OFN414_n_28303), .c(n_1927), .d(FE_OFN134_n_27449), .o(n_25656) );
oa22f80 g544792 ( .a(n_24924), .b(FE_OFN412_n_28303), .c(n_607), .d(FE_OFN113_n_27449), .o(n_25878) );
oa22f80 g544793 ( .a(n_23411), .b(FE_OFN416_n_28303), .c(n_158), .d(FE_OFN102_n_27449), .o(n_24361) );
in01f80 g544871 ( .a(n_22586), .o(n_22587) );
no02f80 g544872 ( .a(FE_OFN542_n_23570), .b(x_in_12_14), .o(n_22586) );
na02f80 g544873 ( .a(FE_OFN542_n_23570), .b(x_in_12_14), .o(n_23241) );
na02f80 g544874 ( .a(FE_OFN542_n_23570), .b(x_in_12_15), .o(n_22274) );
no02f80 g544875 ( .a(n_25348), .b(n_25347), .o(n_25349) );
na02f80 g544876 ( .a(n_23229), .b(n_22926), .o(n_22927) );
no02f80 g544877 ( .a(n_25652), .b(n_25651), .o(n_25653) );
in01f80 g544878 ( .a(n_24084), .o(n_24085) );
no02f80 g544879 ( .a(n_23804), .b(x_in_2_9), .o(n_24084) );
na02f80 g544880 ( .a(n_23804), .b(x_in_2_9), .o(n_24709) );
no02f80 g544881 ( .a(n_25649), .b(n_25648), .o(n_25650) );
in01f80 g544882 ( .a(n_24359), .o(n_24360) );
no02f80 g544883 ( .a(n_24083), .b(x_in_34_9), .o(n_24359) );
na02f80 g544884 ( .a(n_24083), .b(x_in_34_9), .o(n_25033) );
no02f80 g544885 ( .a(n_25646), .b(n_25645), .o(n_25647) );
no02f80 g544886 ( .a(n_25875), .b(n_25874), .o(n_25876) );
no02f80 g544887 ( .a(n_25345), .b(n_25344), .o(n_25346) );
na02f80 g544888 ( .a(n_25021), .b(x_in_8_12), .o(n_25932) );
in01f80 g544889 ( .a(n_25342), .o(n_25343) );
no02f80 g544890 ( .a(n_25021), .b(x_in_8_12), .o(n_25342) );
na02f80 g544891 ( .a(n_23796), .b(x_in_6_9), .o(n_24706) );
in01f80 g544892 ( .a(n_23802), .o(n_23803) );
no02f80 g544893 ( .a(n_23544), .b(x_in_18_9), .o(n_23802) );
na02f80 g544894 ( .a(n_23544), .b(x_in_18_9), .o(n_24399) );
no02f80 g544895 ( .a(n_22931), .b(n_22584), .o(n_22585) );
no02f80 g544896 ( .a(n_23800), .b(n_23799), .o(n_23801) );
na02f80 g544897 ( .a(n_23543), .b(n_23799), .o(n_24808) );
no02f80 g544898 ( .a(n_25643), .b(n_25642), .o(n_25644) );
in01f80 g544899 ( .a(n_23797), .o(n_23798) );
no02f80 g544900 ( .a(n_23542), .b(x_in_50_9), .o(n_23797) );
na02f80 g544901 ( .a(n_23542), .b(x_in_50_9), .o(n_24398) );
in01f80 g544902 ( .a(n_24081), .o(n_24082) );
no02f80 g544903 ( .a(n_23796), .b(x_in_6_9), .o(n_24081) );
no02f80 g544904 ( .a(n_25640), .b(n_25639), .o(n_25641) );
in01f80 g544905 ( .a(n_24079), .o(n_24080) );
no02f80 g544906 ( .a(n_23795), .b(x_in_10_9), .o(n_24079) );
no02f80 g544907 ( .a(n_23558), .b(n_23216), .o(n_23217) );
na02f80 g544908 ( .a(n_23795), .b(x_in_10_9), .o(n_24708) );
no02f80 g544909 ( .a(n_25340), .b(n_25339), .o(n_25341) );
in01f80 g544910 ( .a(n_24077), .o(n_24078) );
no02f80 g544911 ( .a(n_23794), .b(x_in_42_9), .o(n_24077) );
na02f80 g544912 ( .a(n_23794), .b(x_in_42_9), .o(n_24707) );
na02f80 g544913 ( .a(n_23533), .b(x_in_62_9), .o(n_24388) );
no02f80 g544914 ( .a(n_25337), .b(n_25336), .o(n_25338) );
in01f80 g544915 ( .a(n_24075), .o(n_24076) );
no02f80 g544916 ( .a(n_23793), .b(x_in_26_9), .o(n_24075) );
na02f80 g544917 ( .a(n_23793), .b(x_in_26_9), .o(n_24705) );
no02f80 g544918 ( .a(n_23559), .b(n_23214), .o(n_23215) );
no02f80 g544919 ( .a(n_25334), .b(n_25566), .o(n_25335) );
no02f80 g544920 ( .a(n_25332), .b(n_25331), .o(n_25333) );
in01f80 g544921 ( .a(n_23791), .o(n_23792) );
no02f80 g544922 ( .a(n_23541), .b(x_in_58_9), .o(n_23791) );
na02f80 g544923 ( .a(n_23541), .b(x_in_58_9), .o(n_24395) );
no02f80 g544924 ( .a(n_25637), .b(n_25636), .o(n_25638) );
na02f80 g544925 ( .a(n_23539), .b(x_in_2_10), .o(n_24396) );
in01f80 g544926 ( .a(n_24073), .o(n_24074) );
na02f80 g544927 ( .a(n_23790), .b(x_in_6_8), .o(n_24073) );
no02f80 g544928 ( .a(n_23790), .b(x_in_6_8), .o(n_24704) );
in01f80 g544929 ( .a(n_24071), .o(n_24072) );
na02f80 g544930 ( .a(n_23789), .b(n_23162), .o(n_24071) );
no02f80 g544931 ( .a(n_23557), .b(n_23212), .o(n_23213) );
no02f80 g544932 ( .a(n_25329), .b(n_25559), .o(n_25330) );
no02f80 g544933 ( .a(n_25327), .b(n_25326), .o(n_25328) );
in01f80 g544934 ( .a(n_24357), .o(n_24358) );
na02f80 g544935 ( .a(n_24070), .b(n_23444), .o(n_24357) );
na02f80 g544936 ( .a(n_23540), .b(x_in_22_10), .o(n_24389) );
na02f80 g544937 ( .a(n_23788), .b(x_in_22_9), .o(n_24703) );
in01f80 g544938 ( .a(n_24068), .o(n_24069) );
no02f80 g544939 ( .a(n_23788), .b(x_in_22_9), .o(n_24068) );
na02f80 g544940 ( .a(n_23206), .b(x_in_52_9), .o(n_24117) );
in01f80 g544941 ( .a(n_23786), .o(n_23787) );
no02f80 g544942 ( .a(n_23539), .b(x_in_2_10), .o(n_23786) );
in01f80 g544943 ( .a(n_23784), .o(n_23785) );
no02f80 g544944 ( .a(n_23540), .b(x_in_22_10), .o(n_23784) );
no02f80 g544945 ( .a(n_25324), .b(n_25323), .o(n_25325) );
na02f80 g544946 ( .a(n_23538), .b(x_in_54_9), .o(n_24400) );
in01f80 g544947 ( .a(n_23782), .o(n_23783) );
no02f80 g544948 ( .a(n_23538), .b(x_in_54_9), .o(n_23782) );
na02f80 g544949 ( .a(n_23772), .b(x_in_40_9), .o(n_24701) );
in01f80 g544950 ( .a(n_23780), .o(n_23781) );
no02f80 g544951 ( .a(n_23532), .b(x_in_14_9), .o(n_23780) );
no02f80 g544952 ( .a(n_25019), .b(n_25297), .o(n_25020) );
no02f80 g544953 ( .a(n_25624), .b(n_25623), .o(n_25625) );
na02f80 g544954 ( .a(n_23211), .b(x_in_54_10), .o(n_24119) );
in01f80 g544955 ( .a(n_23778), .o(n_23779) );
no02f80 g544956 ( .a(n_23537), .b(x_in_46_9), .o(n_23778) );
na02f80 g544957 ( .a(n_23537), .b(x_in_46_9), .o(n_24397) );
no02f80 g544958 ( .a(n_25321), .b(n_25320), .o(n_25322) );
no02f80 g544959 ( .a(n_25318), .b(n_25317), .o(n_25319) );
in01f80 g544960 ( .a(n_23776), .o(n_23777) );
no02f80 g544961 ( .a(n_23536), .b(x_in_30_9), .o(n_23776) );
na02f80 g544962 ( .a(n_23536), .b(x_in_30_9), .o(n_24394) );
in01f80 g544963 ( .a(n_23534), .o(n_23535) );
no02f80 g544964 ( .a(n_23211), .b(x_in_54_10), .o(n_23534) );
no02f80 g544965 ( .a(n_25315), .b(n_25314), .o(n_25316) );
in01f80 g544966 ( .a(n_23774), .o(n_23775) );
no02f80 g544967 ( .a(n_23533), .b(x_in_62_9), .o(n_23774) );
no02f80 g544968 ( .a(n_23235), .b(n_22924), .o(n_22925) );
na02f80 g544969 ( .a(n_23532), .b(x_in_14_9), .o(n_24401) );
in01f80 g544970 ( .a(n_25617), .o(n_25618) );
no02f80 g544971 ( .a(n_25305), .b(x_in_56_11), .o(n_25617) );
no02f80 g544972 ( .a(n_25615), .b(n_25614), .o(n_25616) );
na02f80 g544973 ( .a(n_23210), .b(x_in_14_10), .o(n_24113) );
no02f80 g544974 ( .a(n_25610), .b(n_25609), .o(n_25611) );
na02f80 g544975 ( .a(n_23773), .b(x_in_34_10), .o(n_24702) );
na02f80 g544976 ( .a(n_24356), .b(x_in_36_9), .o(n_25370) );
in01f80 g544977 ( .a(n_24688), .o(n_24689) );
no02f80 g544978 ( .a(n_24356), .b(x_in_36_9), .o(n_24688) );
in01f80 g544979 ( .a(n_23530), .o(n_23531) );
no02f80 g544980 ( .a(n_23210), .b(x_in_14_10), .o(n_23530) );
no02f80 g544981 ( .a(n_23234), .b(n_22922), .o(n_22923) );
no02f80 g544982 ( .a(n_25017), .b(n_25016), .o(n_25018) );
na02f80 g544983 ( .a(n_23209), .b(x_in_46_10), .o(n_24118) );
in01f80 g544984 ( .a(n_24066), .o(n_24067) );
no02f80 g544985 ( .a(n_23773), .b(x_in_34_10), .o(n_24066) );
in01f80 g544986 ( .a(n_23528), .o(n_23529) );
no02f80 g544987 ( .a(n_23209), .b(x_in_46_10), .o(n_23528) );
no02f80 g544988 ( .a(n_23233), .b(n_22920), .o(n_22921) );
in01f80 g544989 ( .a(n_24064), .o(n_24065) );
no02f80 g544990 ( .a(n_23772), .b(x_in_40_9), .o(n_24064) );
no02f80 g544991 ( .a(n_25598), .b(n_25597), .o(n_25599) );
na02f80 g544992 ( .a(n_23527), .b(x_in_16_10), .o(n_24387) );
in01f80 g544993 ( .a(n_23770), .o(n_23771) );
no02f80 g544994 ( .a(n_23527), .b(x_in_16_10), .o(n_23770) );
no02f80 g544995 ( .a(n_23232), .b(n_22918), .o(n_22919) );
no02f80 g544996 ( .a(n_25014), .b(FE_OFN1252_n_25296), .o(n_25015) );
na02f80 g544997 ( .a(n_23526), .b(x_in_12_10), .o(n_24386) );
no02f80 g544998 ( .a(n_26096), .b(n_26095), .o(n_26097) );
na02f80 g544999 ( .a(n_23523), .b(x_in_18_10), .o(n_24385) );
no02f80 g545000 ( .a(n_25312), .b(n_25311), .o(n_25313) );
na02f80 g545001 ( .a(n_23208), .b(x_in_30_10), .o(n_24116) );
in01f80 g545002 ( .a(n_23524), .o(n_23525) );
no02f80 g545003 ( .a(n_23208), .b(x_in_30_10), .o(n_23524) );
no02f80 g545004 ( .a(n_23231), .b(n_22916), .o(n_22917) );
in01f80 g545005 ( .a(n_23768), .o(n_23769) );
no02f80 g545006 ( .a(n_23523), .b(x_in_18_10), .o(n_23768) );
no02f80 g545007 ( .a(n_25595), .b(n_25594), .o(n_25596) );
na02f80 g545008 ( .a(n_23207), .b(x_in_62_10), .o(n_24115) );
in01f80 g545009 ( .a(n_23521), .o(n_23522) );
no02f80 g545010 ( .a(n_23207), .b(x_in_62_10), .o(n_23521) );
no02f80 g545011 ( .a(n_23230), .b(n_22914), .o(n_22915) );
in01f80 g545012 ( .a(n_23766), .o(n_23767) );
no02f80 g545013 ( .a(n_23526), .b(x_in_12_10), .o(n_23766) );
no02f80 g545014 ( .a(n_25592), .b(n_25591), .o(n_25593) );
in01f80 g545015 ( .a(n_23764), .o(n_23765) );
na02f80 g545016 ( .a(n_23520), .b(x_in_32_8), .o(n_23764) );
no02f80 g545017 ( .a(n_23520), .b(x_in_32_8), .o(n_24383) );
no02f80 g545018 ( .a(n_25309), .b(n_25308), .o(n_25310) );
in01f80 g545019 ( .a(n_23518), .o(n_23519) );
no02f80 g545020 ( .a(n_23206), .b(x_in_52_9), .o(n_23518) );
na02f80 g545021 ( .a(n_23516), .b(x_in_50_10), .o(n_24384) );
no02f80 g545022 ( .a(n_25589), .b(n_25588), .o(n_25590) );
no02f80 g545023 ( .a(n_25012), .b(n_25290), .o(n_25013) );
in01f80 g545024 ( .a(n_23762), .o(n_23763) );
no02f80 g545025 ( .a(n_23517), .b(x_in_16_9), .o(n_23762) );
na02f80 g545026 ( .a(n_23517), .b(x_in_16_9), .o(n_24379) );
no02f80 g545027 ( .a(n_25010), .b(n_25009), .o(n_25011) );
in01f80 g545028 ( .a(n_23760), .o(n_23761) );
no02f80 g545029 ( .a(n_23516), .b(x_in_50_10), .o(n_23760) );
in01f80 g545030 ( .a(n_24354), .o(n_24355) );
no02f80 g545031 ( .a(n_24063), .b(x_in_48_8), .o(n_24354) );
na02f80 g545032 ( .a(n_24063), .b(x_in_48_8), .o(n_25031) );
no02f80 g545033 ( .a(n_25007), .b(n_25006), .o(n_25008) );
na02f80 g545034 ( .a(n_25005), .b(x_in_8_11), .o(n_25930) );
in01f80 g545035 ( .a(n_25306), .o(n_25307) );
no02f80 g545036 ( .a(n_25005), .b(x_in_8_11), .o(n_25306) );
no02f80 g545037 ( .a(n_25586), .b(n_25585), .o(n_25587) );
no02f80 g545038 ( .a(n_24100), .b(n_23758), .o(n_23759) );
na02f80 g545039 ( .a(n_23757), .b(x_in_40_8), .o(n_24700) );
in01f80 g545040 ( .a(n_24061), .o(n_24062) );
no02f80 g545041 ( .a(n_23757), .b(x_in_40_8), .o(n_24061) );
na02f80 g545042 ( .a(n_23515), .b(x_in_32_9), .o(n_24378) );
in01f80 g545043 ( .a(n_23755), .o(n_23756) );
no02f80 g545044 ( .a(n_23515), .b(x_in_32_9), .o(n_23755) );
na02f80 g545045 ( .a(n_25305), .b(x_in_56_11), .o(n_26179) );
no02f80 g545046 ( .a(n_24686), .b(n_24685), .o(n_24687) );
na02f80 g545047 ( .a(n_25004), .b(x_in_44_12), .o(n_25929) );
in01f80 g545048 ( .a(n_25303), .o(n_25304) );
no02f80 g545049 ( .a(n_25004), .b(x_in_44_12), .o(n_25303) );
no02f80 g545050 ( .a(n_24692), .b(n_24352), .o(n_24353) );
in01f80 g545051 ( .a(n_25858), .o(n_25859) );
na02f80 g545052 ( .a(n_25584), .b(n_24975), .o(n_25858) );
no02f80 g545053 ( .a(n_25002), .b(n_25295), .o(n_25003) );
na02f80 g545054 ( .a(n_23514), .b(x_in_10_10), .o(n_24377) );
na02f80 g545055 ( .a(n_25001), .b(x_in_56_10), .o(n_25928) );
in01f80 g545056 ( .a(n_25301), .o(n_25302) );
no02f80 g545057 ( .a(n_25001), .b(x_in_56_10), .o(n_25301) );
in01f80 g545058 ( .a(n_23753), .o(n_23754) );
no02f80 g545059 ( .a(n_23514), .b(x_in_10_10), .o(n_23753) );
na02f80 g545060 ( .a(n_24347), .b(x_in_20_9), .o(n_25371) );
na02f80 g545061 ( .a(n_24060), .b(x_in_48_9), .o(n_25030) );
in01f80 g545062 ( .a(n_24350), .o(n_24351) );
no02f80 g545063 ( .a(n_24060), .b(x_in_48_9), .o(n_24350) );
no02f80 g545064 ( .a(n_25582), .b(n_25581), .o(n_25583) );
na02f80 g545065 ( .a(n_23513), .b(x_in_42_10), .o(n_24376) );
in01f80 g545066 ( .a(n_24348), .o(n_24349) );
na02f80 g545067 ( .a(n_24059), .b(n_23427), .o(n_24348) );
in01f80 g545068 ( .a(n_24683), .o(n_24684) );
no02f80 g545069 ( .a(n_24347), .b(x_in_20_9), .o(n_24683) );
in01f80 g545070 ( .a(n_23751), .o(n_23752) );
no02f80 g545071 ( .a(n_23513), .b(x_in_42_10), .o(n_23751) );
in01f80 g545072 ( .a(n_24681), .o(n_24682) );
na02f80 g545073 ( .a(n_24346), .b(x_in_36_8), .o(n_24681) );
no02f80 g545074 ( .a(n_24346), .b(x_in_36_8), .o(n_25365) );
na02f80 g545075 ( .a(n_24099), .b(n_23749), .o(n_23750) );
no02f80 g545076 ( .a(n_25579), .b(n_25578), .o(n_25580) );
na02f80 g545077 ( .a(n_23509), .b(x_in_26_10), .o(n_24375) );
no02f80 g545078 ( .a(n_23511), .b(n_23510), .o(n_23512) );
na02f80 g545079 ( .a(n_23225), .b(n_22911), .o(n_22912) );
na02f80 g545080 ( .a(n_23205), .b(n_23510), .o(n_24463) );
no02f80 g545081 ( .a(n_25852), .b(n_26050), .o(n_25853) );
na02f80 g545082 ( .a(n_24345), .b(x_in_20_8), .o(n_25364) );
in01f80 g545083 ( .a(n_24679), .o(n_24680) );
no02f80 g545084 ( .a(n_24345), .b(x_in_20_8), .o(n_24679) );
in01f80 g545085 ( .a(n_23747), .o(n_23748) );
no02f80 g545086 ( .a(n_23509), .b(x_in_26_10), .o(n_23747) );
no02f80 g545087 ( .a(n_23507), .b(n_23506), .o(n_23508) );
na02f80 g545088 ( .a(n_23204), .b(n_23506), .o(n_24461) );
no02f80 g545089 ( .a(n_25850), .b(n_25849), .o(n_25851) );
in01f80 g545090 ( .a(n_23504), .o(n_23505) );
na02f80 g545091 ( .a(n_23203), .b(x_in_52_8), .o(n_23504) );
no02f80 g545092 ( .a(n_23203), .b(x_in_52_8), .o(n_24110) );
no02f80 g545093 ( .a(n_24677), .b(n_24991), .o(n_24678) );
in01f80 g545094 ( .a(n_24057), .o(n_24058) );
no02f80 g545095 ( .a(n_23746), .b(x_in_12_9), .o(n_24057) );
na02f80 g545096 ( .a(n_23746), .b(x_in_12_9), .o(n_24699) );
no02f80 g545097 ( .a(n_25576), .b(n_25575), .o(n_25577) );
na02f80 g545098 ( .a(n_23503), .b(x_in_58_10), .o(n_24374) );
no02f80 g545099 ( .a(n_24999), .b(n_25293), .o(n_25000) );
in01f80 g545100 ( .a(n_25573), .o(n_25574) );
na02f80 g545101 ( .a(n_25300), .b(n_24655), .o(n_25573) );
na02f80 g545102 ( .a(n_25299), .b(x_in_44_11), .o(n_26171) );
in01f80 g545103 ( .a(n_25571), .o(n_25572) );
no02f80 g545104 ( .a(n_25299), .b(x_in_44_11), .o(n_25571) );
in01f80 g545105 ( .a(n_23744), .o(n_23745) );
no02f80 g545106 ( .a(n_23503), .b(x_in_58_10), .o(n_23744) );
in01f80 g545107 ( .a(n_24343), .o(n_24344) );
na02f80 g545108 ( .a(n_24056), .b(n_23423), .o(n_24343) );
na02f80 g545109 ( .a(n_24055), .b(x_in_60_9), .o(n_25032) );
in01f80 g545110 ( .a(n_24341), .o(n_24342) );
no02f80 g545111 ( .a(n_24055), .b(x_in_60_9), .o(n_24341) );
no02f80 g545112 ( .a(n_23236), .b(n_22909), .o(n_22910) );
in01f80 g545113 ( .a(n_24675), .o(n_24676) );
no02f80 g545114 ( .a(n_24340), .b(x_in_60_8), .o(n_24675) );
na02f80 g545115 ( .a(n_24340), .b(x_in_60_8), .o(n_25372) );
no02f80 g545116 ( .a(n_23556), .b(n_23201), .o(n_23202) );
no02f80 g545117 ( .a(n_23227), .b(n_22907), .o(n_22908) );
no02f80 g545118 ( .a(n_22929), .b(n_22582), .o(n_22583) );
no02f80 g545119 ( .a(n_23825), .b(n_23501), .o(n_23502) );
no02f80 g545120 ( .a(n_25028), .b(n_24673), .o(n_24674) );
no02f80 g545121 ( .a(n_24338), .b(n_24337), .o(n_24339) );
in01f80 g545122 ( .a(n_24335), .o(n_24336) );
na02f80 g545123 ( .a(n_24338), .b(n_24054), .o(n_24335) );
no02f80 g545124 ( .a(n_23555), .b(n_23199), .o(n_23200) );
no02f80 g545125 ( .a(n_23153), .b(n_26312), .o(n_23743) );
no02f80 g545126 ( .a(n_23226), .b(n_22905), .o(n_22906) );
na02f80 g545127 ( .a(n_24098), .b(n_23741), .o(n_23742) );
no02f80 g545128 ( .a(n_23224), .b(n_22903), .o(n_22904) );
no02f80 g545129 ( .a(n_23553), .b(n_23197), .o(n_23198) );
no02f80 g545130 ( .a(n_22930), .b(n_22580), .o(n_22581) );
na02f80 g545131 ( .a(n_23208), .b(n_23495), .o(n_23196) );
na02f80 g545132 ( .a(n_23540), .b(n_23740), .o(n_23500) );
na02f80 g545133 ( .a(n_23142), .b(n_23740), .o(n_24740) );
na02f80 g545134 ( .a(n_23211), .b(n_23499), .o(n_23195) );
na02f80 g545135 ( .a(n_22865), .b(n_23499), .o(n_24451) );
na02f80 g545136 ( .a(n_23210), .b(n_23498), .o(n_23194) );
na02f80 g545137 ( .a(n_22864), .b(n_23498), .o(n_24448) );
na02f80 g545138 ( .a(n_22863), .b(n_23497), .o(n_24449) );
na02f80 g545139 ( .a(n_23207), .b(n_23496), .o(n_23193) );
na02f80 g545140 ( .a(n_22860), .b(n_23496), .o(n_24454) );
na02f80 g545141 ( .a(n_23209), .b(n_23497), .o(n_23192) );
na02f80 g545142 ( .a(n_22861), .b(n_23495), .o(n_24450) );
na02f80 g545143 ( .a(n_23526), .b(n_23739), .o(n_23494) );
na02f80 g545144 ( .a(n_23141), .b(n_23739), .o(n_24739) );
no02f80 g545145 ( .a(n_23823), .b(n_23492), .o(n_23493) );
no02f80 g545146 ( .a(n_23223), .b(n_22901), .o(n_22902) );
no02f80 g545147 ( .a(n_23222), .b(n_22899), .o(n_22900) );
na02f80 g545148 ( .a(n_23554), .b(n_23190), .o(n_23191) );
no02f80 g545149 ( .a(n_24333), .b(n_24332), .o(n_24334) );
na02f80 g545150 ( .a(n_24053), .b(n_24332), .o(n_25378) );
na02f80 g545151 ( .a(n_24997), .b(n_25004), .o(n_24998) );
na02f80 g545152 ( .a(n_24997), .b(n_24672), .o(n_25943) );
no02f80 g545153 ( .a(n_24670), .b(n_24669), .o(n_24671) );
na02f80 g545154 ( .a(n_24996), .b(n_24320), .o(n_28633) );
no02f80 g545155 ( .a(n_23221), .b(n_22897), .o(n_22898) );
no02f80 g545156 ( .a(n_23220), .b(n_22895), .o(n_22896) );
no02f80 g545157 ( .a(n_23219), .b(n_22893), .o(n_22894) );
no02f80 g545158 ( .a(n_23737), .b(n_23736), .o(n_23738) );
na02f80 g545159 ( .a(n_23491), .b(n_23736), .o(n_25051) );
no02f80 g545160 ( .a(n_23218), .b(n_22891), .o(n_22892) );
no02f80 g545161 ( .a(n_23548), .b(n_23188), .o(n_23189) );
no02f80 g545162 ( .a(n_22555), .b(n_23188), .o(n_24148) );
na02f80 g545163 ( .a(n_25021), .b(n_25298), .o(n_24995) );
na02f80 g545164 ( .a(n_24628), .b(n_25298), .o(n_26169) );
na02f80 g545165 ( .a(n_23822), .b(n_23489), .o(n_23490) );
na02f80 g545166 ( .a(n_23237), .b(n_22889), .o(n_22890) );
no02f80 g545167 ( .a(n_25567), .b(n_25844), .o(n_25568) );
no02f80 g545168 ( .a(n_23487), .b(n_23486), .o(n_23488) );
no02f80 g545169 ( .a(n_23487), .b(n_22769), .o(n_24736) );
na02f80 g545170 ( .a(n_23186), .b(n_23485), .o(n_23187) );
in01f80 g545171 ( .a(n_23735), .o(n_24434) );
no02f80 g545172 ( .a(n_23539), .b(n_23485), .o(n_23735) );
na02f80 g545173 ( .a(n_23483), .b(n_23734), .o(n_23484) );
in01f80 g545174 ( .a(n_24052), .o(n_24732) );
no02f80 g545175 ( .a(n_23773), .b(n_23734), .o(n_24052) );
na02f80 g545176 ( .a(n_23481), .b(n_23480), .o(n_23482) );
na02f80 g545177 ( .a(n_23481), .b(n_22765), .o(n_24433) );
na02f80 g545178 ( .a(n_23478), .b(n_23477), .o(n_23479) );
in01f80 g545179 ( .a(n_26210), .o(n_25845) );
oa12f80 g545180 ( .a(n_23118), .b(n_25566), .c(n_23708), .o(n_26210) );
na02f80 g545181 ( .a(n_23478), .b(n_22764), .o(n_24432) );
no02f80 g545182 ( .a(n_23732), .b(n_23731), .o(n_23733) );
in01f80 g545183 ( .a(n_23730), .o(n_24429) );
na02f80 g545184 ( .a(n_23476), .b(n_23731), .o(n_23730) );
na02f80 g545185 ( .a(n_23184), .b(n_23475), .o(n_23185) );
in01f80 g545186 ( .a(n_23729), .o(n_24426) );
no02f80 g545187 ( .a(n_23514), .b(n_23475), .o(n_23729) );
na02f80 g545188 ( .a(n_23182), .b(n_23474), .o(n_23183) );
in01f80 g545189 ( .a(n_23728), .o(n_24423) );
no02f80 g545190 ( .a(n_23513), .b(n_23474), .o(n_23728) );
na02f80 g545191 ( .a(n_23180), .b(n_23473), .o(n_23181) );
in01f80 g545192 ( .a(n_23727), .o(n_24420) );
no02f80 g545193 ( .a(n_23509), .b(n_23473), .o(n_23727) );
na02f80 g545194 ( .a(n_23471), .b(n_23470), .o(n_23472) );
na02f80 g545195 ( .a(n_23468), .b(n_23726), .o(n_23469) );
in01f80 g545196 ( .a(n_25960), .o(n_25565) );
oa12f80 g545197 ( .a(n_22822), .b(n_25297), .c(n_23449), .o(n_25960) );
na02f80 g545198 ( .a(n_23471), .b(n_22763), .o(n_24419) );
in01f80 g545199 ( .a(n_26473), .o(n_26066) );
oa12f80 g545200 ( .a(n_23685), .b(n_24322), .c(n_25844), .o(n_26473) );
in01f80 g545201 ( .a(n_24051), .o(n_24726) );
no02f80 g545202 ( .a(n_23796), .b(n_23726), .o(n_24051) );
in01f80 g545203 ( .a(n_25957), .o(n_25564) );
oa12f80 g545204 ( .a(n_22545), .b(FE_OFN1252_n_25296), .c(n_23160), .o(n_25957) );
in01f80 g545205 ( .a(n_23725), .o(n_24416) );
no02f80 g545206 ( .a(n_23515), .b(n_23467), .o(n_23725) );
na02f80 g545207 ( .a(n_23178), .b(n_23467), .o(n_23179) );
no02f80 g545208 ( .a(n_22887), .b(n_22886), .o(n_22888) );
no02f80 g545209 ( .a(n_22887), .b(n_22204), .o(n_24139) );
na02f80 g545210 ( .a(n_23465), .b(n_23464), .o(n_23466) );
na02f80 g545211 ( .a(n_23465), .b(n_22762), .o(n_24415) );
na02f80 g545212 ( .a(n_24049), .b(n_24048), .o(n_24050) );
na02f80 g545213 ( .a(n_24049), .b(n_23379), .o(n_25048) );
no02f80 g545214 ( .a(n_23462), .b(n_23461), .o(n_23463) );
in01f80 g545215 ( .a(n_23460), .o(n_24132) );
na02f80 g545216 ( .a(n_23177), .b(n_23461), .o(n_23460) );
na02f80 g545217 ( .a(n_23723), .b(n_23722), .o(n_23724) );
na02f80 g545218 ( .a(n_23723), .b(n_23092), .o(n_24722) );
in01f80 g545219 ( .a(n_25950), .o(n_25563) );
oa12f80 g545220 ( .a(n_22795), .b(n_23429), .c(n_25295), .o(n_25950) );
na02f80 g545221 ( .a(n_24993), .b(n_25294), .o(n_24994) );
no02f80 g545222 ( .a(n_25305), .b(n_25294), .o(n_25976) );
no02f80 g545223 ( .a(n_23175), .b(n_23174), .o(n_23176) );
no02f80 g545224 ( .a(n_23175), .b(n_22476), .o(n_24410) );
ao12f80 g545225 ( .a(n_9555), .b(n_22885), .c(n_11590), .o(n_23842) );
na02f80 g545226 ( .a(n_24046), .b(n_24331), .o(n_24047) );
no02f80 g545227 ( .a(n_24356), .b(n_24331), .o(n_25376) );
na02f80 g545228 ( .a(n_24329), .b(n_24328), .o(n_24330) );
na02f80 g545229 ( .a(n_24329), .b(n_23664), .o(n_25375) );
na02f80 g545230 ( .a(n_22883), .b(n_23173), .o(n_22884) );
in01f80 g545231 ( .a(n_23459), .o(n_24128) );
no02f80 g545232 ( .a(n_23206), .b(n_23173), .o(n_23459) );
no02f80 g545233 ( .a(n_23171), .b(n_23170), .o(n_23172) );
no02f80 g545234 ( .a(n_23171), .b(n_22472), .o(n_24406) );
in01f80 g545235 ( .a(n_25945), .o(n_25562) );
oa12f80 g545236 ( .a(n_23098), .b(n_25293), .c(n_23700), .o(n_25945) );
ao22s80 g545237 ( .a(n_21192), .b(n_21563), .c(x_out_44_32), .d(FE_OFN318_n_27400), .o(n_22273) );
na02f80 g545238 ( .a(n_23720), .b(n_24045), .o(n_23721) );
in01f80 g545239 ( .a(n_24327), .o(n_25041) );
no02f80 g545240 ( .a(n_24055), .b(n_24045), .o(n_24327) );
in01f80 g545241 ( .a(n_26753), .o(n_26348) );
oa12f80 g545242 ( .a(n_23451), .b(n_22844), .c(n_25251), .o(n_26753) );
in01f80 g545243 ( .a(n_26750), .o(n_26347) );
oa12f80 g545244 ( .a(n_23710), .b(n_23124), .c(n_25250), .o(n_26750) );
in01f80 g545245 ( .a(n_26747), .o(n_26346) );
oa12f80 g545246 ( .a(n_23709), .b(n_23122), .c(n_25248), .o(n_26747) );
in01f80 g545247 ( .a(n_26744), .o(n_26345) );
oa12f80 g545248 ( .a(n_23704), .b(n_23120), .c(n_25247), .o(n_26744) );
in01f80 g545249 ( .a(n_26512), .o(n_26065) );
oa12f80 g545250 ( .a(n_23448), .b(n_24914), .c(n_22836), .o(n_26512) );
in01f80 g545251 ( .a(n_26509), .o(n_26064) );
oa12f80 g545252 ( .a(n_23447), .b(n_24913), .c(n_22834), .o(n_26509) );
in01f80 g545253 ( .a(n_26505), .o(n_26063) );
oa12f80 g545254 ( .a(n_23446), .b(n_24912), .c(n_22832), .o(n_26505) );
in01f80 g545255 ( .a(n_26502), .o(n_26062) );
oa12f80 g545256 ( .a(n_23707), .b(n_24911), .c(n_23116), .o(n_26502) );
in01f80 g545257 ( .a(n_26061), .o(n_26982) );
oa12f80 g545258 ( .a(n_21886), .b(n_25833), .c(n_21111), .o(n_26061) );
in01f80 g545259 ( .a(n_26498), .o(n_26060) );
oa12f80 g545260 ( .a(n_23701), .b(n_23112), .c(n_24909), .o(n_26498) );
in01f80 g545261 ( .a(n_26734), .o(n_26344) );
oa12f80 g545262 ( .a(n_23439), .b(n_22828), .c(n_25246), .o(n_26734) );
in01f80 g545263 ( .a(n_26495), .o(n_26059) );
oa12f80 g545264 ( .a(n_23445), .b(n_22826), .c(n_24908), .o(n_26495) );
in01f80 g545265 ( .a(n_26731), .o(n_26343) );
oa12f80 g545266 ( .a(n_23711), .b(n_23126), .c(n_25244), .o(n_26731) );
in01f80 g545267 ( .a(n_26492), .o(n_26058) );
oa12f80 g545268 ( .a(n_23442), .b(n_22820), .c(n_24907), .o(n_26492) );
in01f80 g545269 ( .a(n_26486), .o(n_26057) );
oa12f80 g545270 ( .a(n_23452), .b(n_22818), .c(n_24906), .o(n_26486) );
in01f80 g545271 ( .a(n_26728), .o(n_26342) );
oa12f80 g545272 ( .a(n_23440), .b(n_22816), .c(n_25243), .o(n_26728) );
in01f80 g545273 ( .a(n_26489), .o(n_26056) );
oa12f80 g545274 ( .a(n_23441), .b(n_22814), .c(n_24905), .o(n_26489) );
in01f80 g545275 ( .a(n_25843), .o(n_26689) );
oa12f80 g545276 ( .a(n_21049), .b(n_25555), .c(n_20701), .o(n_25843) );
in01f80 g545277 ( .a(n_26205), .o(n_25842) );
oa12f80 g545278 ( .a(n_23438), .b(n_22812), .c(n_24580), .o(n_26205) );
in01f80 g545279 ( .a(n_27233), .o(n_26946) );
oa12f80 g545280 ( .a(n_23705), .b(n_23108), .c(n_25798), .o(n_27233) );
in01f80 g545281 ( .a(n_26725), .o(n_26341) );
oa12f80 g545282 ( .a(n_23437), .b(n_22809), .c(n_25242), .o(n_26725) );
in01f80 g545283 ( .a(n_26483), .o(n_26055) );
oa12f80 g545284 ( .a(n_23436), .b(n_22807), .c(n_24904), .o(n_26483) );
oa12f80 g545285 ( .a(n_12463), .b(n_23169), .c(n_13641), .o(n_24125) );
in01f80 g545286 ( .a(n_26722), .o(n_26340) );
oa12f80 g545287 ( .a(n_23435), .b(n_22805), .c(n_25241), .o(n_26722) );
in01f80 g545288 ( .a(n_26480), .o(n_26054) );
oa12f80 g545289 ( .a(n_23433), .b(n_22803), .c(n_24903), .o(n_26480) );
in01f80 g545290 ( .a(n_26719), .o(n_26339) );
oa12f80 g545291 ( .a(n_23434), .b(n_22800), .c(n_25240), .o(n_26719) );
in01f80 g545292 ( .a(n_26202), .o(n_25841) );
oa12f80 g545293 ( .a(n_23702), .b(n_23106), .c(n_24579), .o(n_26202) );
in01f80 g545294 ( .a(n_25561), .o(n_26457) );
oa12f80 g545295 ( .a(n_18483), .b(n_25287), .c(n_17902), .o(n_25561) );
in01f80 g545296 ( .a(n_26199), .o(n_25840) );
oa12f80 g545297 ( .a(n_23703), .b(n_23104), .c(n_24576), .o(n_26199) );
in01f80 g545298 ( .a(n_26716), .o(n_26338) );
oa12f80 g545299 ( .a(n_23430), .b(n_22797), .c(n_25239), .o(n_26716) );
in01f80 g545300 ( .a(n_25292), .o(n_26188) );
oa12f80 g545301 ( .a(n_3154), .b(n_24988), .c(n_2154), .o(n_25292) );
in01f80 g545302 ( .a(n_26053), .o(n_26980) );
oa12f80 g545303 ( .a(n_23282), .b(n_25831), .c(n_22636), .o(n_26053) );
in01f80 g545304 ( .a(n_25954), .o(n_25560) );
oa12f80 g545305 ( .a(n_24031), .b(n_23397), .c(n_24222), .o(n_25954) );
in01f80 g545306 ( .a(n_26737), .o(n_26337) );
oa12f80 g545307 ( .a(n_23706), .b(n_23110), .c(n_25245), .o(n_26737) );
in01f80 g545308 ( .a(n_25838), .o(n_26691) );
oa12f80 g545309 ( .a(n_22125), .b(n_25557), .c(n_21446), .o(n_25838) );
in01f80 g545310 ( .a(n_25291), .o(n_26186) );
oa12f80 g545311 ( .a(n_22129), .b(n_24986), .c(n_21432), .o(n_25291) );
ao12f80 g545312 ( .a(n_13622), .b(n_23168), .c(n_14266), .o(n_24124) );
in01f80 g545313 ( .a(n_26713), .o(n_26336) );
oa12f80 g545314 ( .a(n_23428), .b(n_25238), .c(n_22793), .o(n_26713) );
in01f80 g545315 ( .a(n_27003), .o(n_26623) );
oa12f80 g545316 ( .a(n_24323), .b(n_23672), .c(n_25521), .o(n_27003) );
in01f80 g545317 ( .a(n_25837), .o(n_26686) );
oa12f80 g545318 ( .a(n_22128), .b(n_25553), .c(n_21428), .o(n_25837) );
in01f80 g545319 ( .a(n_26710), .o(n_26335) );
oa12f80 g545320 ( .a(n_23425), .b(n_25237), .c(n_22788), .o(n_26710) );
in01f80 g545321 ( .a(n_26994), .o(n_26622) );
oa12f80 g545322 ( .a(n_24656), .b(n_23962), .c(n_25519), .o(n_26994) );
in01f80 g545323 ( .a(n_26705), .o(n_26334) );
oa12f80 g545324 ( .a(n_23424), .b(n_25236), .c(n_22784), .o(n_26705) );
oa12f80 g545325 ( .a(FE_OFN1113_rst), .b(n_22270), .c(n_22578), .o(n_22579) );
in01f80 g545326 ( .a(n_25836), .o(n_26684) );
oa12f80 g545327 ( .a(n_23274), .b(n_25551), .c(n_22633), .o(n_25836) );
in01f80 g545328 ( .a(n_25835), .o(n_26682) );
oa12f80 g545329 ( .a(n_22123), .b(n_25549), .c(n_21423), .o(n_25835) );
in01f80 g545330 ( .a(n_26468), .o(n_26052) );
oa12f80 g545331 ( .a(n_23450), .b(n_24901), .c(n_22781), .o(n_26468) );
in01f80 g545332 ( .a(n_26740), .o(n_26333) );
oa12f80 g545333 ( .a(n_24035), .b(n_23384), .c(n_25235), .o(n_26740) );
in01f80 g545334 ( .a(n_26756), .o(n_26332) );
oa12f80 g545335 ( .a(n_24036), .b(n_23382), .c(n_25234), .o(n_26756) );
oa12f80 g545336 ( .a(n_22881), .b(n_1213), .c(FE_OFN116_n_27449), .o(n_22882) );
in01f80 g545337 ( .a(n_23563), .o(n_23167) );
ao12f80 g545338 ( .a(n_10815), .b(n_22880), .c(n_12052), .o(n_23563) );
ao22s80 g545339 ( .a(n_24992), .b(x_in_5_15), .c(n_23952), .d(x_in_4_14), .o(n_25703) );
ao12f80 g545340 ( .a(n_9531), .b(n_22577), .c(n_11520), .o(n_23239) );
ao12f80 g545341 ( .a(n_12470), .b(n_23166), .c(n_13662), .o(n_23835) );
ao12f80 g545342 ( .a(n_22775), .b(n_23418), .c(n_25290), .o(n_26193) );
ao12f80 g545343 ( .a(n_22506), .b(n_24991), .c(n_23151), .o(n_25939) );
oa12f80 g545344 ( .a(n_9104), .b(n_24990), .c(n_10789), .o(n_25700) );
oa12f80 g545345 ( .a(n_11144), .b(n_24044), .c(n_12732), .o(n_24694) );
ao12f80 g545346 ( .a(n_23421), .b(n_23420), .c(n_23419), .o(n_24043) );
in01f80 g545347 ( .a(n_23561), .o(n_23827) );
ao12f80 g545348 ( .a(n_22272), .b(n_22577), .c(n_22271), .o(n_23561) );
ao22s80 g545349 ( .a(n_22143), .b(n_25833), .c(n_22142), .d(n_24910), .o(n_25834) );
ao12f80 g545350 ( .a(n_22566), .b(n_22567), .c(n_22565), .o(n_23165) );
ao22s80 g545351 ( .a(n_24571), .b(n_23694), .c(n_25559), .d(x_in_6_7), .o(n_26466) );
in01f80 g545352 ( .a(n_23830), .o(n_24121) );
ao12f80 g545353 ( .a(n_22573), .b(n_22880), .c(n_22572), .o(n_23830) );
oa12f80 g545354 ( .a(n_22869), .b(n_22879), .c(n_23149), .o(n_24120) );
ao22s80 g545355 ( .a(n_22410), .b(n_25557), .c(n_22409), .d(n_24578), .o(n_25558) );
ao22s80 g545356 ( .a(n_25555), .b(n_21394), .c(n_24577), .d(n_21393), .o(n_25556) );
in01f80 g545357 ( .a(n_23719), .o(n_24712) );
oa12f80 g545358 ( .a(n_22873), .b(n_23166), .c(n_22872), .o(n_23719) );
ao12f80 g545359 ( .a(n_24034), .b(n_24033), .c(n_24032), .o(n_24668) );
ao12f80 g545360 ( .a(n_24653), .b(n_24992), .c(n_24652), .o(n_25289) );
in01f80 g545361 ( .a(n_24114), .o(n_24381) );
ao12f80 g545362 ( .a(n_22878), .b(n_23169), .c(n_22877), .o(n_24114) );
ao22s80 g545363 ( .a(n_25287), .b(n_18770), .c(n_24223), .d(n_18769), .o(n_25288) );
ao12f80 g545364 ( .a(n_23432), .b(n_23715), .c(n_23431), .o(n_24042) );
ao22s80 g545365 ( .a(n_24988), .b(n_3616), .c(n_23947), .d(n_3615), .o(n_24989) );
in01f80 g545366 ( .a(n_25926), .o(n_26180) );
ao12f80 g545367 ( .a(n_24651), .b(n_24990), .c(n_24650), .o(n_25926) );
ao12f80 g545368 ( .a(n_23699), .b(n_24038), .c(n_23698), .o(n_24326) );
oa12f80 g545369 ( .a(n_23697), .b(n_24044), .c(n_23696), .o(n_25029) );
ao12f80 g545370 ( .a(n_23156), .b(n_23155), .c(n_23154), .o(n_23718) );
in01f80 g545371 ( .a(n_23458), .o(n_24104) );
ao12f80 g545372 ( .a(n_22571), .b(n_22574), .c(n_22570), .o(n_23458) );
ao12f80 g545373 ( .a(n_23417), .b(n_23416), .c(n_23415), .o(n_24041) );
in01f80 g545374 ( .a(n_24102), .o(n_23717) );
oa12f80 g545375 ( .a(n_22876), .b(n_23168), .c(n_22875), .o(n_24102) );
ao22s80 g545376 ( .a(n_25831), .b(n_23604), .c(n_24902), .d(n_23603), .o(n_25832) );
ao22s80 g545377 ( .a(n_22419), .b(n_24986), .c(n_22418), .d(n_23946), .o(n_24987) );
ao22s80 g545378 ( .a(n_22417), .b(n_25553), .c(n_22416), .d(n_24575), .o(n_25554) );
in01f80 g545379 ( .a(n_23836), .o(n_23457) );
oa12f80 g545380 ( .a(n_22569), .b(n_22885), .c(n_22568), .o(n_23836) );
ao22s80 g545381 ( .a(n_25231), .b(n_24311), .c(n_26050), .d(x_in_36_7), .o(n_26993) );
ao22s80 g545382 ( .a(n_25551), .b(n_23602), .c(n_24574), .d(n_23601), .o(n_25552) );
oa12f80 g545383 ( .a(n_22871), .b(n_22870), .c(n_23150), .o(n_24109) );
ao22s80 g545384 ( .a(n_22406), .b(n_25549), .c(n_22405), .d(n_24573), .o(n_25550) );
oa22f80 g545385 ( .a(n_23082), .b(FE_OFN411_n_28303), .c(n_1023), .d(FE_OFN129_n_27449), .o(n_24040) );
oa22f80 g545386 ( .a(n_22193), .b(FE_OFN412_n_28303), .c(n_816), .d(FE_OFN91_n_27449), .o(n_23164) );
oa22f80 g545387 ( .a(n_24568), .b(FE_OFN157_n_28014), .c(n_481), .d(FE_OFN96_n_27449), .o(n_25548) );
oa22f80 g545388 ( .a(n_24038), .b(FE_OFN406_n_28303), .c(n_1833), .d(FE_OFN99_n_27449), .o(n_24039) );
oa22f80 g545389 ( .a(n_24054), .b(FE_OFN406_n_28303), .c(n_1045), .d(n_28607), .o(n_24325) );
oa22f80 g545390 ( .a(n_22471), .b(FE_OFN248_n_4162), .c(n_291), .d(FE_OFN92_n_27449), .o(n_23456) );
oa22f80 g545391 ( .a(n_24221), .b(FE_OFN410_n_28303), .c(n_1714), .d(FE_OFN63_n_27012), .o(n_25286) );
oa22f80 g545392 ( .a(n_22874), .b(FE_OFN249_n_4162), .c(n_1709), .d(FE_OFN65_n_27012), .o(n_23163) );
oa22f80 g545393 ( .a(n_23148), .b(FE_OFN409_n_28303), .c(n_1787), .d(FE_OFN355_n_4860), .o(n_23455) );
oa22f80 g545394 ( .a(FE_OFN452_n_23152), .b(FE_OFN411_n_28303), .c(n_499), .d(n_27709), .o(n_23454) );
oa22f80 g545395 ( .a(n_24217), .b(FE_OFN251_n_4162), .c(n_1696), .d(FE_OFN93_n_27449), .o(n_25284) );
oa22f80 g545396 ( .a(n_23662), .b(FE_OFN248_n_4162), .c(n_1741), .d(FE_OFN60_n_27012), .o(n_24667) );
oa22f80 g545397 ( .a(n_23715), .b(FE_OFN404_n_28303), .c(n_403), .d(FE_OFN286_n_29266), .o(n_23716) );
oa22f80 g545398 ( .a(n_23943), .b(FE_OFN410_n_28303), .c(n_518), .d(FE_OFN286_n_29266), .o(n_24985) );
oa22f80 g545399 ( .a(n_23081), .b(n_4280), .c(n_899), .d(n_28607), .o(n_24037) );
oa22f80 g545400 ( .a(FE_OFN426_n_23661), .b(FE_OFN406_n_28303), .c(n_1182), .d(n_28607), .o(n_24666) );
oa22f80 g545401 ( .a(n_23372), .b(FE_OFN404_n_28303), .c(n_908), .d(n_29261), .o(n_24324) );
oa22f80 g545402 ( .a(n_22757), .b(FE_OFN405_n_28303), .c(n_785), .d(FE_OFN89_n_27449), .o(n_23714) );
oa22f80 g545403 ( .a(n_22756), .b(FE_OFN409_n_28303), .c(n_729), .d(FE_OFN125_n_27449), .o(n_23713) );
oa22f80 g545404 ( .a(n_24566), .b(FE_OFN412_n_28303), .c(n_400), .d(FE_OFN65_n_27012), .o(n_25547) );
oa22f80 g545405 ( .a(n_23659), .b(FE_OFN251_n_4162), .c(n_1136), .d(FE_OFN93_n_27449), .o(n_24665) );
oa22f80 g545406 ( .a(n_23657), .b(FE_OFN248_n_4162), .c(n_612), .d(FE_OFN90_n_27449), .o(n_24663) );
oa22f80 g545407 ( .a(n_24214), .b(FE_OFN247_n_4162), .c(n_477), .d(FE_OFN134_n_27449), .o(n_25283) );
oa22f80 g545408 ( .a(n_21562), .b(n_4162), .c(n_453), .d(FE_OFN116_n_27449), .o(n_22576) );
oa22f80 g545409 ( .a(n_23941), .b(FE_OFN249_n_4162), .c(n_1554), .d(FE_OFN1111_rst), .o(n_24983) );
oa22f80 g545410 ( .a(n_24211), .b(FE_OFN249_n_4162), .c(n_1899), .d(FE_OFN1111_rst), .o(n_25282) );
oa22f80 g545411 ( .a(n_24209), .b(FE_OFN402_n_28303), .c(n_1525), .d(FE_OFN1123_rst), .o(n_25280) );
ao22s80 g545412 ( .a(n_23663), .b(x_in_24_15), .c(n_24030), .d(n_2545), .o(n_28849) );
no02f80 g545441 ( .a(n_22574), .b(n_8911), .o(n_22575) );
na02f80 g545442 ( .a(n_23452), .b(n_22819), .o(n_25315) );
na02f80 g545443 ( .a(n_24036), .b(n_23383), .o(n_25652) );
na02f80 g545444 ( .a(n_23711), .b(n_23127), .o(n_25589) );
na02f80 g545445 ( .a(n_23451), .b(n_22845), .o(n_25649) );
na02f80 g545446 ( .a(n_24323), .b(n_23673), .o(n_25875) );
na02f80 g545447 ( .a(n_23710), .b(n_23125), .o(n_25646) );
na02f80 g545448 ( .a(n_23450), .b(n_22782), .o(n_25345) );
in01f80 g545449 ( .a(n_25278), .o(n_25279) );
na02f80 g545450 ( .a(n_24982), .b(n_24277), .o(n_25278) );
no02f80 g545451 ( .a(n_22823), .b(n_23449), .o(n_25019) );
na02f80 g545452 ( .a(n_23709), .b(n_23123), .o(n_25643) );
na02f80 g545453 ( .a(n_23448), .b(n_22837), .o(n_25340) );
na02f80 g545454 ( .a(n_23447), .b(n_22835), .o(n_25337) );
no02f80 g545455 ( .a(n_23119), .b(n_23708), .o(n_25334) );
na02f80 g545456 ( .a(n_23446), .b(n_22833), .o(n_25332) );
na02f80 g545457 ( .a(n_24035), .b(n_23385), .o(n_25637) );
na02f80 g545458 ( .a(n_23707), .b(n_23117), .o(n_25348) );
na02f80 g545459 ( .a(n_22879), .b(x_in_38_12), .o(n_23789) );
in01f80 g545460 ( .a(n_23161), .o(n_23162) );
no02f80 g545461 ( .a(n_22879), .b(x_in_38_12), .o(n_23161) );
no02f80 g545462 ( .a(n_22880), .b(n_22572), .o(n_22573) );
na02f80 g545463 ( .a(n_23445), .b(n_22827), .o(n_25327) );
in01f80 g545464 ( .a(n_23443), .o(n_23444) );
no02f80 g545465 ( .a(n_23159), .b(x_in_38_11), .o(n_23443) );
na02f80 g545466 ( .a(n_23706), .b(n_23111), .o(n_25624) );
na02f80 g545467 ( .a(n_23442), .b(n_22821), .o(n_25318) );
na02f80 g545468 ( .a(n_23441), .b(n_22815), .o(n_25321) );
in01f80 g545469 ( .a(n_25276), .o(n_25277) );
na02f80 g545470 ( .a(n_24981), .b(n_24259), .o(n_25276) );
na02f80 g545471 ( .a(n_23440), .b(n_22817), .o(n_25615) );
na02f80 g545472 ( .a(n_23439), .b(n_22829), .o(n_25610) );
no02f80 g545473 ( .a(n_24033), .b(n_24032), .o(n_24034) );
no02f80 g545474 ( .a(n_23686), .b(n_24322), .o(n_25567) );
na02f80 g545475 ( .a(n_23438), .b(n_22813), .o(n_25017) );
na02f80 g545476 ( .a(n_23437), .b(n_22810), .o(n_25598) );
no02f80 g545477 ( .a(n_22546), .b(n_23160), .o(n_25014) );
na02f80 g545478 ( .a(n_23705), .b(n_23109), .o(n_26096) );
no02f80 g545479 ( .a(n_23169), .b(n_22877), .o(n_22878) );
na02f80 g545480 ( .a(n_23436), .b(n_22808), .o(n_25312) );
na02f80 g545481 ( .a(n_23435), .b(n_22806), .o(n_25595) );
na02f80 g545482 ( .a(n_23704), .b(n_23121), .o(n_25640) );
na02f80 g545483 ( .a(n_23434), .b(n_22801), .o(n_25592) );
na02f80 g545484 ( .a(n_23433), .b(n_22804), .o(n_25309) );
na02f80 g545485 ( .a(n_23159), .b(x_in_38_11), .o(n_24070) );
no02f80 g545486 ( .a(n_23715), .b(n_23431), .o(n_23432) );
no02f80 g545487 ( .a(n_22758), .b(n_23431), .o(n_24380) );
na02f80 g545488 ( .a(n_23703), .b(n_23105), .o(n_25010) );
na02f80 g545489 ( .a(n_23702), .b(n_23107), .o(n_25007) );
in01f80 g545490 ( .a(n_24661), .o(n_24662) );
na02f80 g545491 ( .a(n_24321), .b(n_23681), .o(n_24661) );
in01f80 g545492 ( .a(n_24979), .o(n_24980) );
na02f80 g545493 ( .a(n_24660), .b(n_23978), .o(n_24979) );
na02f80 g545494 ( .a(n_23430), .b(n_22798), .o(n_25586) );
in01f80 g545495 ( .a(n_25274), .o(n_25275) );
na02f80 g545496 ( .a(n_24978), .b(n_24237), .o(n_25274) );
na02f80 g545497 ( .a(n_24031), .b(n_23398), .o(n_24686) );
in01f80 g545498 ( .a(n_24976), .o(n_24977) );
na02f80 g545499 ( .a(n_24659), .b(n_23972), .o(n_24976) );
na02f80 g545500 ( .a(n_24658), .b(x_in_24_13), .o(n_25584) );
in01f80 g545501 ( .a(n_24974), .o(n_24975) );
no02f80 g545502 ( .a(n_24658), .b(x_in_24_13), .o(n_24974) );
na02f80 g545503 ( .a(n_24030), .b(n_24029), .o(n_24996) );
in01f80 g545504 ( .a(n_24319), .o(n_24320) );
no02f80 g545505 ( .a(n_24030), .b(n_24029), .o(n_24319) );
na02f80 g545506 ( .a(n_23168), .b(n_22875), .o(n_22876) );
no02f80 g545507 ( .a(n_22796), .b(n_23429), .o(n_25002) );
in01f80 g545508 ( .a(n_24972), .o(n_24973) );
na02f80 g545509 ( .a(n_24657), .b(n_23968), .o(n_24972) );
na02f80 g545510 ( .a(n_23428), .b(n_22794), .o(n_25582) );
in01f80 g545511 ( .a(n_24317), .o(n_24318) );
na02f80 g545512 ( .a(n_24028), .b(n_23392), .o(n_24317) );
na02f80 g545513 ( .a(n_23158), .b(x_in_28_12), .o(n_24059) );
in01f80 g545514 ( .a(n_23426), .o(n_23427) );
no02f80 g545515 ( .a(n_23158), .b(x_in_28_12), .o(n_23426) );
na02f80 g545516 ( .a(n_23701), .b(n_23113), .o(n_25324) );
na02f80 g545517 ( .a(n_23425), .b(n_22789), .o(n_25579) );
na02f80 g545518 ( .a(n_24656), .b(n_23963), .o(n_25850) );
na02f80 g545519 ( .a(n_23424), .b(n_22785), .o(n_25576) );
no02f80 g545520 ( .a(n_23099), .b(n_23700), .o(n_24999) );
na02f80 g545521 ( .a(n_24316), .b(x_in_44_10), .o(n_25300) );
in01f80 g545522 ( .a(n_24654), .o(n_24655) );
no02f80 g545523 ( .a(n_24316), .b(x_in_44_10), .o(n_24654) );
na02f80 g545524 ( .a(n_23157), .b(x_in_28_11), .o(n_24056) );
in01f80 g545525 ( .a(n_23422), .o(n_23423) );
no02f80 g545526 ( .a(n_23157), .b(x_in_28_11), .o(n_23422) );
na02f80 g545527 ( .a(n_23378), .b(n_24019), .o(n_25028) );
no02f80 g545528 ( .a(n_22577), .b(n_22271), .o(n_22272) );
no02f80 g545529 ( .a(n_24038), .b(n_23698), .o(n_23699) );
no02f80 g545530 ( .a(n_23080), .b(n_23698), .o(n_24338) );
no02f80 g545531 ( .a(n_23155), .b(n_23154), .o(n_23156) );
in01f80 g545532 ( .a(n_24107), .o(n_23153) );
na02f80 g545533 ( .a(n_22874), .b(n_23154), .o(n_24107) );
no02f80 g545534 ( .a(n_24992), .b(n_24652), .o(n_24653) );
na02f80 g545535 ( .a(n_23166), .b(n_22872), .o(n_22873) );
no02f80 g545536 ( .a(n_24990), .b(n_24650), .o(n_24651) );
no02f80 g545537 ( .a(n_23420), .b(n_23419), .o(n_23421) );
na02f80 g545538 ( .a(n_23152), .b(n_23419), .o(n_24370) );
na02f80 g545539 ( .a(n_24044), .b(n_23696), .o(n_23697) );
na02f80 g545540 ( .a(n_22776), .b(n_23418), .o(n_25012) );
na02f80 g545541 ( .a(n_22507), .b(n_23151), .o(n_24677) );
no02f80 g545542 ( .a(n_22574), .b(n_22570), .o(n_22571) );
na02f80 g545543 ( .a(n_22870), .b(n_23150), .o(n_22871) );
no02f80 g545544 ( .a(n_23158), .b(n_23150), .o(n_24106) );
na02f80 g545545 ( .a(n_22885), .b(n_22568), .o(n_22569) );
na02f80 g545546 ( .a(n_22470), .b(n_23149), .o(n_24105) );
na02f80 g545547 ( .a(n_22879), .b(n_23149), .o(n_22869) );
na02f80 g545548 ( .a(n_22270), .b(FE_OFN1113_rst), .o(n_22881) );
no02f80 g545549 ( .a(n_22567), .b(n_21916), .o(n_23826) );
no02f80 g545550 ( .a(n_22567), .b(n_22565), .o(n_22566) );
in01f80 g545551 ( .a(FE_OFN542_n_23570), .o(n_21979) );
ao22s80 g545552 ( .a(n_20475), .b(n_9618), .c(n_2835), .d(x_in_13_15), .o(n_23570) );
oa12f80 g545553 ( .a(n_12929), .b(n_23695), .c(n_14462), .o(n_24692) );
no02f80 g545554 ( .a(n_23416), .b(n_23415), .o(n_23417) );
in01f80 g545555 ( .a(n_23414), .o(n_24101) );
na02f80 g545556 ( .a(n_23148), .b(n_23415), .o(n_23414) );
in01f80 g545557 ( .a(n_25823), .o(n_26673) );
oa12f80 g545558 ( .a(n_23362), .b(n_22729), .c(n_25539), .o(n_25823) );
oa12f80 g545559 ( .a(n_13220), .b(n_22564), .c(n_14292), .o(n_23559) );
oa12f80 g545560 ( .a(n_16386), .b(n_22563), .c(n_16904), .o(n_23558) );
ao12f80 g545561 ( .a(n_15563), .b(n_21978), .c(n_16266), .o(n_22931) );
oa12f80 g545562 ( .a(n_15344), .b(n_22562), .c(n_14782), .o(n_23557) );
oa12f80 g545563 ( .a(n_15431), .b(n_22269), .c(n_14770), .o(n_23235) );
in01f80 g545564 ( .a(n_25273), .o(n_26160) );
oa12f80 g545565 ( .a(n_23651), .b(n_23016), .c(n_24949), .o(n_25273) );
oa12f80 g545566 ( .a(n_15355), .b(n_22268), .c(n_14727), .o(n_23234) );
ao12f80 g545567 ( .a(n_14746), .b(n_22267), .c(n_15400), .o(n_23233) );
ao12f80 g545568 ( .a(n_15145), .b(n_22266), .c(n_14385), .o(n_23232) );
ao12f80 g545569 ( .a(n_14718), .b(n_22265), .c(n_15388), .o(n_23231) );
oa12f80 g545570 ( .a(n_15376), .b(n_22264), .c(n_14692), .o(n_23230) );
in01f80 g545571 ( .a(n_24647), .o(n_25691) );
oa12f80 g545572 ( .a(n_23071), .b(n_24312), .c(n_22423), .o(n_24647) );
in01f80 g545573 ( .a(n_22868), .o(n_23819) );
oa12f80 g545574 ( .a(n_13158), .b(n_22561), .c(n_14314), .o(n_22868) );
in01f80 g545575 ( .a(n_25543), .o(n_26432) );
oa12f80 g545576 ( .a(n_23359), .b(n_22679), .c(n_25260), .o(n_25543) );
ao12f80 g545577 ( .a(n_15793), .b(n_23147), .c(n_16472), .o(n_24100) );
in01f80 g545578 ( .a(n_25272), .o(n_26150) );
oa12f80 g545579 ( .a(n_23356), .b(n_22671), .c(n_24932), .o(n_25272) );
in01f80 g545580 ( .a(n_25271), .o(n_26147) );
oa12f80 g545581 ( .a(n_23064), .b(n_22413), .c(n_24928), .o(n_25271) );
ao12f80 g545582 ( .a(n_15780), .b(n_23146), .c(n_16471), .o(n_24099) );
oa12f80 g545583 ( .a(n_11427), .b(n_22263), .c(n_12481), .o(n_23229) );
ao12f80 g545584 ( .a(n_12932), .b(n_22262), .c(n_12250), .o(n_23225) );
ao12f80 g545585 ( .a(n_15085), .b(n_22261), .c(n_14222), .o(n_23236) );
oa12f80 g545586 ( .a(n_14724), .b(n_22560), .c(n_15389), .o(n_23556) );
oa12f80 g545587 ( .a(n_14360), .b(n_22260), .c(n_15136), .o(n_23227) );
ao12f80 g545588 ( .a(n_11511), .b(n_21977), .c(n_12047), .o(n_22929) );
oa12f80 g545589 ( .a(n_16089), .b(n_22867), .c(n_16674), .o(n_23825) );
oa12f80 g545590 ( .a(n_15291), .b(n_22559), .c(n_16032), .o(n_23555) );
ao12f80 g545591 ( .a(n_13198), .b(n_22259), .c(n_14391), .o(n_23226) );
oa12f80 g545592 ( .a(n_13189), .b(n_23145), .c(n_14364), .o(n_24098) );
oa12f80 g545593 ( .a(n_10936), .b(n_22855), .c(n_9175), .o(n_23822) );
oa12f80 g545594 ( .a(n_14958), .b(n_22258), .c(n_13999), .o(n_23224) );
oa12f80 g545595 ( .a(n_11342), .b(n_24026), .c(n_12827), .o(n_24027) );
ao12f80 g545596 ( .a(n_14425), .b(n_22558), .c(n_15160), .o(n_23553) );
oa12f80 g545597 ( .a(n_11787), .b(n_21976), .c(n_10652), .o(n_22930) );
oa12f80 g545598 ( .a(n_13167), .b(n_22866), .c(n_14329), .o(n_23823) );
oa12f80 g545599 ( .a(n_14260), .b(n_22257), .c(n_15104), .o(n_23223) );
ao12f80 g545600 ( .a(n_14913), .b(n_22256), .c(n_13905), .o(n_23222) );
ao12f80 g545601 ( .a(n_12495), .b(n_22557), .c(n_11518), .o(n_23554) );
oa12f80 g545602 ( .a(n_15526), .b(n_22255), .c(n_16259), .o(n_23221) );
ao12f80 g545603 ( .a(n_14908), .b(n_22254), .c(n_13884), .o(n_23220) );
oa12f80 g545604 ( .a(n_14936), .b(n_22253), .c(n_13964), .o(n_23219) );
oa12f80 g545605 ( .a(n_10663), .b(n_22252), .c(n_11798), .o(n_23218) );
ao12f80 g545606 ( .a(n_10801), .b(n_22251), .c(n_11185), .o(n_23237) );
ao12f80 g545607 ( .a(n_22772), .b(n_22771), .c(n_22770), .o(n_23413) );
ao12f80 g545608 ( .a(n_24286), .b(n_24285), .c(n_24284), .o(n_24971) );
in01f80 g545609 ( .a(n_23204), .o(n_23507) );
ao12f80 g545610 ( .a(n_21975), .b(n_22263), .c(n_21974), .o(n_23204) );
oa12f80 g545611 ( .a(n_22504), .b(n_22503), .c(n_22502), .o(n_23804) );
ao12f80 g545612 ( .a(n_24283), .b(n_24282), .c(n_24281), .o(n_24970) );
oa12f80 g545613 ( .a(n_22768), .b(n_22767), .c(n_22766), .o(n_24083) );
ao12f80 g545614 ( .a(n_23381), .b(n_23692), .c(n_23380), .o(n_24025) );
ao12f80 g545615 ( .a(n_24593), .b(n_24592), .c(n_24591), .o(n_25270) );
ao12f80 g545616 ( .a(n_24280), .b(n_24279), .c(n_24278), .o(n_24969) );
ao12f80 g545617 ( .a(n_24018), .b(n_24017), .c(n_24016), .o(n_24646) );
ao22s80 g545618 ( .a(n_23650), .b(n_25539), .c(n_23649), .d(n_24556), .o(n_25540) );
in01f80 g545619 ( .a(n_23468), .o(n_23796) );
ao12f80 g545620 ( .a(n_22248), .b(n_22563), .c(n_22247), .o(n_23468) );
oa12f80 g545621 ( .a(n_22216), .b(n_22215), .c(n_22501), .o(n_23544) );
ao12f80 g545622 ( .a(n_22841), .b(n_23134), .c(n_22840), .o(n_23412) );
ao12f80 g545623 ( .a(n_24275), .b(n_24274), .c(n_24273), .o(n_24968) );
oa12f80 g545624 ( .a(n_22214), .b(n_22213), .c(n_22500), .o(n_23542) );
ao12f80 g545625 ( .a(n_22499), .b(n_22498), .c(n_22497), .o(n_23144) );
ao12f80 g545626 ( .a(n_24272), .b(n_24271), .c(n_24270), .o(n_24967) );
oa12f80 g545627 ( .a(n_22496), .b(n_22495), .c(n_22494), .o(n_23795) );
ao12f80 g545628 ( .a(n_24014), .b(n_24013), .c(n_24012), .o(n_24645) );
oa12f80 g545629 ( .a(n_22493), .b(n_22492), .c(n_22491), .o(n_23794) );
ao12f80 g545630 ( .a(n_23966), .b(n_23965), .c(n_23964), .o(n_24644) );
oa12f80 g545631 ( .a(n_22490), .b(n_22489), .c(n_22488), .o(n_23793) );
in01f80 g545632 ( .a(n_23487), .o(n_23143) );
oa12f80 g545633 ( .a(n_22246), .b(n_22564), .c(n_22245), .o(n_23487) );
ao12f80 g545634 ( .a(n_24269), .b(n_24268), .c(n_24572), .o(n_24965) );
ao12f80 g545635 ( .a(n_24011), .b(n_24010), .c(n_24009), .o(n_24643) );
ao12f80 g545636 ( .a(n_24267), .b(n_24266), .c(n_24265), .o(n_24964) );
ao12f80 g545637 ( .a(n_23992), .b(n_23991), .c(n_23990), .o(n_24642) );
ao12f80 g545638 ( .a(n_24006), .b(n_24005), .c(n_24004), .o(n_24641) );
oa12f80 g545639 ( .a(n_23094), .b(n_23694), .c(x_in_6_7), .o(n_25329) );
in01f80 g545640 ( .a(n_23540), .o(n_23142) );
oa12f80 g545641 ( .a(n_22244), .b(n_22562), .c(n_22243), .o(n_23540) );
oa12f80 g545642 ( .a(n_22520), .b(n_22519), .c(n_22778), .o(n_23788) );
in01f80 g545643 ( .a(n_22883), .o(n_23206) );
ao12f80 g545644 ( .a(n_21570), .b(n_21978), .c(n_21569), .o(n_22883) );
ao12f80 g545645 ( .a(n_23961), .b(n_23960), .c(n_23959), .o(n_24639) );
oa12f80 g545646 ( .a(n_22233), .b(n_22232), .c(n_22518), .o(n_23538) );
ao12f80 g545647 ( .a(n_24003), .b(n_24002), .c(n_24001), .o(n_24638) );
ao12f80 g545648 ( .a(n_24008), .b(n_24007), .c(n_24218), .o(n_24637) );
oa12f80 g545649 ( .a(n_22229), .b(n_22228), .c(n_22514), .o(n_23532) );
ao12f80 g545650 ( .a(n_24289), .b(n_24288), .c(n_24287), .o(n_24957) );
in01f80 g545651 ( .a(n_23211), .o(n_22865) );
oa12f80 g545652 ( .a(n_21973), .b(n_22269), .c(n_21972), .o(n_23211) );
oa12f80 g545653 ( .a(n_22231), .b(n_22230), .c(n_22515), .o(n_23537) );
ao12f80 g545654 ( .a(n_24000), .b(n_23999), .c(n_23998), .o(n_24636) );
oa12f80 g545655 ( .a(n_22227), .b(n_22226), .c(n_22517), .o(n_23536) );
ao12f80 g545656 ( .a(n_23997), .b(n_23996), .c(n_23995), .o(n_24635) );
oa12f80 g545657 ( .a(n_22225), .b(n_22224), .c(n_22516), .o(n_23533) );
ao12f80 g545658 ( .a(n_23989), .b(n_23988), .c(n_23987), .o(n_24634) );
in01f80 g545659 ( .a(n_23186), .o(n_23539) );
ao12f80 g545660 ( .a(n_21953), .b(n_22258), .c(n_21952), .o(n_23186) );
ao12f80 g545661 ( .a(n_24257), .b(n_24256), .c(n_24255), .o(n_24951) );
in01f80 g545662 ( .a(n_23210), .o(n_22864) );
oa12f80 g545663 ( .a(n_21963), .b(n_22268), .c(n_21962), .o(n_23210) );
ao22s80 g545664 ( .a(n_23933), .b(n_24949), .c(n_23932), .d(n_23931), .o(n_24950) );
ao12f80 g545665 ( .a(n_24254), .b(n_24253), .c(n_24252), .o(n_24948) );
in01f80 g545666 ( .a(n_23483), .o(n_23773) );
ao12f80 g545667 ( .a(n_22235), .b(n_22558), .c(n_22234), .o(n_23483) );
ao12f80 g545668 ( .a(n_24590), .b(n_24589), .c(n_24900), .o(n_25265) );
ao12f80 g545669 ( .a(n_23951), .b(n_23950), .c(n_24225), .o(n_24633) );
in01f80 g545670 ( .a(n_23209), .o(n_22863) );
oa12f80 g545671 ( .a(n_21971), .b(n_22267), .c(n_21970), .o(n_23209) );
in01f80 g545672 ( .a(n_23171), .o(n_22862) );
oa12f80 g545673 ( .a(n_21955), .b(n_22259), .c(n_21954), .o(n_23171) );
ao12f80 g545674 ( .a(n_24251), .b(n_24250), .c(n_24249), .o(n_24946) );
in01f80 g545675 ( .a(n_23465), .o(n_23527) );
ao12f80 g545676 ( .a(n_21969), .b(n_22266), .c(n_21968), .o(n_23465) );
ao12f80 g545677 ( .a(n_23986), .b(n_24219), .c(n_23985), .o(n_24632) );
in01f80 g545678 ( .a(n_24053), .o(n_24333) );
ao12f80 g545679 ( .a(n_22780), .b(n_23145), .c(n_22779), .o(n_24053) );
in01f80 g545680 ( .a(n_23526), .o(n_23141) );
oa12f80 g545681 ( .a(n_22239), .b(n_22560), .c(n_22238), .o(n_23526) );
ao12f80 g545682 ( .a(n_24917), .b(n_24916), .c(n_24915), .o(n_25538) );
in01f80 g545683 ( .a(n_23481), .o(n_23523) );
ao12f80 g545684 ( .a(n_21957), .b(n_22260), .c(n_21956), .o(n_23481) );
ao12f80 g545685 ( .a(n_23984), .b(n_23983), .c(n_23982), .o(n_24631) );
in01f80 g545686 ( .a(n_23208), .o(n_22861) );
oa12f80 g545687 ( .a(n_21967), .b(n_22265), .c(n_21966), .o(n_23208) );
ao12f80 g545688 ( .a(n_24248), .b(n_24247), .c(n_24246), .o(n_24945) );
in01f80 g545689 ( .a(n_23207), .o(n_22860) );
oa12f80 g545690 ( .a(n_21965), .b(n_22264), .c(n_21964), .o(n_23207) );
oa12f80 g545691 ( .a(n_22212), .b(n_22211), .c(n_22487), .o(n_23541) );
ao12f80 g545692 ( .a(n_24245), .b(n_24244), .c(n_24243), .o(n_24944) );
in01f80 g545693 ( .a(n_23543), .o(n_23800) );
ao12f80 g545694 ( .a(n_22221), .b(n_22557), .c(n_22220), .o(n_23543) );
oa12f80 g545695 ( .a(n_22209), .b(n_22483), .c(n_22208), .o(n_23520) );
ao12f80 g545696 ( .a(n_23981), .b(n_23980), .c(n_23979), .o(n_24630) );
in01f80 g545697 ( .a(n_23478), .o(n_23516) );
ao12f80 g545698 ( .a(n_21943), .b(n_22253), .c(n_21942), .o(n_23478) );
ao12f80 g545699 ( .a(n_22207), .b(n_22206), .c(n_22205), .o(n_22859) );
ao12f80 g545700 ( .a(n_23689), .b(n_23688), .c(n_23687), .o(n_24315) );
oa12f80 g545701 ( .a(n_22203), .b(n_22202), .c(n_22482), .o(n_23517) );
ao12f80 g545702 ( .a(n_23684), .b(n_23683), .c(n_23682), .o(n_24314) );
in01f80 g545703 ( .a(n_24049), .o(n_24060) );
ao12f80 g545704 ( .a(n_22511), .b(n_22866), .c(n_22510), .o(n_24049) );
oa12f80 g545705 ( .a(n_22761), .b(n_22760), .c(n_23093), .o(n_24063) );
ao12f80 g545706 ( .a(n_23949), .b(n_23948), .c(n_24224), .o(n_24629) );
ao12f80 g545707 ( .a(n_22201), .b(n_22200), .c(n_22199), .o(n_22858) );
in01f80 g545708 ( .a(n_23177), .o(n_23462) );
ao12f80 g545709 ( .a(n_21941), .b(n_22251), .c(n_21940), .o(n_23177) );
ao22s80 g545710 ( .a(n_23361), .b(n_24312), .c(n_23360), .d(n_23344), .o(n_24313) );
oa12f80 g545711 ( .a(n_23669), .b(n_23668), .c(n_23953), .o(n_25005) );
in01f80 g545712 ( .a(n_23476), .o(n_23732) );
ao12f80 g545713 ( .a(n_22241), .b(n_22561), .c(n_22240), .o(n_23476) );
in01f80 g545714 ( .a(n_25021), .o(n_24628) );
oa12f80 g545715 ( .a(n_23691), .b(n_23690), .c(n_23956), .o(n_25021) );
ao12f80 g545716 ( .a(n_24242), .b(n_24241), .c(n_24240), .o(n_24940) );
ao22s80 g545717 ( .a(n_23648), .b(n_25260), .c(n_23647), .d(n_24205), .o(n_25261) );
in01f80 g545718 ( .a(n_23723), .o(n_23772) );
ao12f80 g545719 ( .a(n_22237), .b(n_22559), .c(n_22236), .o(n_23723) );
oa12f80 g545720 ( .a(n_22481), .b(n_22480), .c(n_22759), .o(n_23757) );
in01f80 g545721 ( .a(n_23178), .o(n_23515) );
ao12f80 g545722 ( .a(n_21947), .b(n_22255), .c(n_21946), .o(n_23178) );
ao12f80 g545723 ( .a(n_23396), .b(n_23395), .c(n_23394), .o(n_24024) );
in01f80 g545724 ( .a(n_24672), .o(n_25004) );
ao12f80 g545725 ( .a(n_23406), .b(n_23695), .c(n_23405), .o(n_24672) );
in01f80 g545726 ( .a(n_22887), .o(n_22556) );
oa12f80 g545727 ( .a(n_21568), .b(n_21977), .c(n_21567), .o(n_22887) );
ao12f80 g545728 ( .a(n_23970), .b(n_23969), .c(n_24215), .o(n_24626) );
in01f80 g545729 ( .a(n_23184), .o(n_23514) );
ao12f80 g545730 ( .a(n_21951), .b(n_22257), .c(n_21950), .o(n_23184) );
oa12f80 g545731 ( .a(n_23667), .b(n_23666), .c(n_23665), .o(n_25001) );
in01f80 g545732 ( .a(n_24993), .o(n_25305) );
ao12f80 g545733 ( .a(n_23675), .b(n_24026), .c(n_23674), .o(n_24993) );
ao12f80 g545734 ( .a(n_22479), .b(n_22478), .c(n_22477), .o(n_23140) );
in01f80 g545735 ( .a(n_23175), .o(n_22857) );
oa12f80 g545736 ( .a(n_21939), .b(n_22252), .c(n_21938), .o(n_23175) );
in01f80 g545737 ( .a(n_24329), .o(n_24347) );
ao12f80 g545738 ( .a(n_22792), .b(n_23147), .c(n_22791), .o(n_24329) );
ao22s80 g545739 ( .a(n_23646), .b(n_24932), .c(n_23645), .d(n_23930), .o(n_24933) );
ao12f80 g545740 ( .a(n_24235), .b(n_24234), .c(n_24233), .o(n_24930) );
ao22s80 g545741 ( .a(n_23355), .b(n_24928), .c(n_23354), .d(n_23929), .o(n_24929) );
in01f80 g545742 ( .a(n_23182), .o(n_23513) );
ao12f80 g545743 ( .a(n_21949), .b(n_22256), .c(n_21948), .o(n_23182) );
ao12f80 g545744 ( .a(n_22219), .b(n_22218), .c(n_22217), .o(n_22856) );
in01f80 g545745 ( .a(n_22555), .o(n_23548) );
oa12f80 g545746 ( .a(n_21566), .b(n_21976), .c(n_21565), .o(n_22555) );
in01f80 g545747 ( .a(n_24046), .o(n_24356) );
ao12f80 g545748 ( .a(n_22787), .b(n_23146), .c(n_22786), .o(n_24046) );
ao12f80 g545749 ( .a(n_24264), .b(n_24263), .c(n_24262), .o(n_24927) );
oa12f80 g545750 ( .a(n_23090), .b(n_23091), .c(n_23089), .o(n_24346) );
ao12f80 g545751 ( .a(n_24232), .b(n_24231), .c(n_24230), .o(n_24926) );
in01f80 g545752 ( .a(n_23491), .o(n_23737) );
ao22s80 g545753 ( .a(n_21915), .b(n_11588), .c(n_22855), .d(n_11589), .o(n_23491) );
in01f80 g545754 ( .a(n_23180), .o(n_23509) );
ao12f80 g545755 ( .a(n_21945), .b(n_22254), .c(n_21944), .o(n_23180) );
ao12f80 g545756 ( .a(n_22528), .b(n_22850), .c(n_22527), .o(n_23139) );
in01f80 g545757 ( .a(n_23205), .o(n_23511) );
ao12f80 g545758 ( .a(n_21961), .b(n_22262), .c(n_21960), .o(n_23205) );
ao12f80 g545759 ( .a(n_24588), .b(n_24587), .c(n_24586), .o(n_25259) );
oa12f80 g545760 ( .a(n_23670), .b(n_24311), .c(x_in_36_7), .o(n_25852) );
oa12f80 g545761 ( .a(n_23088), .b(n_23087), .c(n_23375), .o(n_24345) );
ao12f80 g545762 ( .a(n_22525), .b(n_22853), .c(n_22524), .o(n_23138) );
ao12f80 g545763 ( .a(n_24585), .b(n_24584), .c(n_24583), .o(n_25258) );
oa12f80 g545764 ( .a(n_22486), .b(n_22485), .c(n_22484), .o(n_23790) );
oa12f80 g545765 ( .a(n_21935), .b(n_22197), .c(n_21934), .o(n_23203) );
ao12f80 g545766 ( .a(n_22475), .b(n_22474), .c(n_22473), .o(n_23137) );
ao12f80 g545767 ( .a(n_23390), .b(n_23389), .c(n_23388), .o(n_24023) );
oa12f80 g545768 ( .a(n_22513), .b(n_22512), .c(n_22777), .o(n_23746) );
ao12f80 g545769 ( .a(n_24229), .b(n_24228), .c(n_24227), .o(n_24925) );
in01f80 g545770 ( .a(n_23471), .o(n_23503) );
ao12f80 g545771 ( .a(n_21959), .b(n_22261), .c(n_21958), .o(n_23471) );
ao12f80 g545772 ( .a(n_23958), .b(n_23957), .c(n_24212), .o(n_24625) );
in01f80 g545773 ( .a(n_25299), .o(n_24924) );
oa12f80 g545774 ( .a(n_23955), .b(n_23954), .c(n_24020), .o(n_25299) );
ao12f80 g545775 ( .a(n_22774), .b(n_23130), .c(n_22773), .o(n_23411) );
in01f80 g545776 ( .a(n_23720), .o(n_24055) );
ao12f80 g545777 ( .a(n_22522), .b(n_22867), .c(n_22521), .o(n_23720) );
oa12f80 g545778 ( .a(n_23086), .b(n_23085), .c(n_23084), .o(n_24340) );
oa22f80 g545779 ( .a(n_22167), .b(FE_OFN251_n_4162), .c(n_646), .d(FE_OFN14_n_29068), .o(n_23136) );
oa22f80 g545780 ( .a(n_23638), .b(FE_OFN251_n_4162), .c(n_1530), .d(FE_OFN14_n_29068), .o(n_24624) );
oa22f80 g545781 ( .a(n_22853), .b(FE_OFN247_n_4162), .c(n_915), .d(FE_OFN364_n_4860), .o(n_22854) );
oa22f80 g545782 ( .a(FE_OFN434_n_23637), .b(n_28608), .c(n_1067), .d(n_28928), .o(n_24623) );
oa22f80 g545783 ( .a(n_23928), .b(FE_OFN247_n_4162), .c(n_1403), .d(FE_OFN134_n_27449), .o(n_24923) );
oa22f80 g545784 ( .a(n_23060), .b(FE_OFN244_n_4162), .c(n_366), .d(FE_OFN139_n_27449), .o(n_24022) );
oa22f80 g545785 ( .a(FE_OFN728_n_23636), .b(FE_OFN230_n_4162), .c(n_504), .d(n_28607), .o(n_24621) );
oa22f80 g545786 ( .a(n_23342), .b(FE_OFN267_n_4280), .c(n_803), .d(FE_OFN329_n_4860), .o(n_24310) );
oa22f80 g545787 ( .a(n_24204), .b(FE_OFN406_n_28303), .c(n_1003), .d(FE_OFN360_n_4860), .o(n_25257) );
oa22f80 g545788 ( .a(n_22435), .b(FE_OFN179_n_27681), .c(n_1201), .d(FE_OFN1174_n_4860), .o(n_23410) );
oa22f80 g545789 ( .a(n_23635), .b(FE_OFN179_n_27681), .c(n_1412), .d(FE_OFN131_n_27449), .o(n_24620) );
oa22f80 g545790 ( .a(n_22434), .b(n_4162), .c(n_1332), .d(FE_OFN116_n_27449), .o(n_23409) );
oa22f80 g545791 ( .a(n_23634), .b(FE_OFN235_n_4162), .c(n_131), .d(FE_OFN114_n_27449), .o(n_24619) );
oa22f80 g545792 ( .a(n_23341), .b(FE_OFN410_n_28303), .c(n_1781), .d(FE_OFN350_n_4860), .o(n_24309) );
oa22f80 g545793 ( .a(n_23340), .b(FE_OFN400_n_28303), .c(n_324), .d(FE_OFN1114_rst), .o(n_24308) );
oa22f80 g545794 ( .a(n_22505), .b(FE_OFN268_n_4280), .c(n_1603), .d(FE_OFN330_n_4860), .o(n_22852) );
oa22f80 g545795 ( .a(n_23633), .b(FE_OFN257_n_4280), .c(n_1351), .d(FE_OFN1108_rst), .o(n_24618) );
oa22f80 g545796 ( .a(n_23339), .b(n_28303), .c(n_244), .d(FE_OFN1109_rst), .o(n_24307) );
oa22f80 g545797 ( .a(n_23632), .b(FE_OFN409_n_28303), .c(n_1360), .d(FE_OFN65_n_27012), .o(n_24617) );
oa22f80 g545798 ( .a(n_23338), .b(FE_OFN267_n_4280), .c(n_391), .d(FE_OFN113_n_27449), .o(n_24306) );
oa22f80 g545799 ( .a(n_23337), .b(FE_OFN411_n_28303), .c(n_1879), .d(n_29104), .o(n_24305) );
oa22f80 g545800 ( .a(FE_OFN650_n_23576), .b(n_28303), .c(n_1370), .d(n_29104), .o(n_24304) );
oa22f80 g545801 ( .a(n_23281), .b(FE_OFN417_n_28303), .c(n_475), .d(FE_OFN101_n_27449), .o(n_24303) );
oa22f80 g545802 ( .a(FE_OFN807_n_23617), .b(n_23291), .c(n_362), .d(n_27449), .o(n_24616) );
oa22f80 g545803 ( .a(n_23631), .b(FE_OFN404_n_28303), .c(n_951), .d(FE_OFN133_n_27449), .o(n_24614) );
oa22f80 g545804 ( .a(n_23453), .b(FE_OFN236_n_4162), .c(n_1225), .d(FE_OFN125_n_27449), .o(n_24302) );
oa22f80 g545805 ( .a(FE_OFN849_n_23567), .b(n_21988), .c(n_1200), .d(FE_OFN56_n_27012), .o(n_24301) );
oa22f80 g545806 ( .a(n_23248), .b(FE_OFN266_n_4280), .c(n_1193), .d(n_29261), .o(n_24300) );
oa22f80 g545807 ( .a(n_23333), .b(n_21988), .c(n_282), .d(FE_OFN347_n_4860), .o(n_24299) );
oa22f80 g545808 ( .a(n_23639), .b(FE_OFN230_n_4162), .c(n_1419), .d(FE_OFN352_n_4860), .o(n_24613) );
oa22f80 g545809 ( .a(n_22198), .b(n_4162), .c(n_106), .d(FE_OFN115_n_27449), .o(n_22554) );
oa22f80 g545810 ( .a(n_23630), .b(FE_OFN247_n_4162), .c(n_1907), .d(FE_OFN128_n_27449), .o(n_24612) );
oa22f80 g545811 ( .a(FE_OFN1005_n_23624), .b(FE_OFN235_n_4162), .c(n_1682), .d(n_27709), .o(n_24611) );
oa22f80 g545812 ( .a(n_22850), .b(FE_OFN234_n_4162), .c(n_493), .d(FE_OFN286_n_29266), .o(n_22851) );
oa22f80 g545813 ( .a(n_23927), .b(n_28303), .c(n_1310), .d(FE_OFN68_n_27012), .o(n_24921) );
oa22f80 g545814 ( .a(n_22196), .b(FE_OFN175_n_26184), .c(n_779), .d(FE_OFN74_n_27012), .o(n_22553) );
oa22f80 g545815 ( .a(FE_OFN556_n_23580), .b(FE_OFN405_n_28303), .c(n_1683), .d(n_29264), .o(n_24610) );
oa22f80 g545816 ( .a(n_23640), .b(FE_OFN236_n_4162), .c(n_565), .d(FE_OFN357_n_4860), .o(n_24609) );
oa22f80 g545817 ( .a(n_23336), .b(FE_OFN239_n_4162), .c(n_1443), .d(FE_OFN130_n_27449), .o(n_24298) );
oa22f80 g545818 ( .a(n_23692), .b(n_23291), .c(n_596), .d(FE_OFN95_n_27449), .o(n_23693) );
oa22f80 g545819 ( .a(n_24200), .b(FE_OFN244_n_4162), .c(n_562), .d(FE_OFN361_n_4860), .o(n_25256) );
oa22f80 g545820 ( .a(n_23335), .b(FE_OFN413_n_28303), .c(n_496), .d(FE_OFN350_n_4860), .o(n_24297) );
oa22f80 g545821 ( .a(n_23629), .b(FE_OFN411_n_28303), .c(n_1943), .d(FE_OFN129_n_27449), .o(n_24608) );
oa22f80 g545822 ( .a(n_23628), .b(FE_OFN293_n_3069), .c(n_1573), .d(FE_OFN89_n_27449), .o(n_24606) );
oa22f80 g545823 ( .a(n_23134), .b(FE_OFN311_n_3069), .c(n_633), .d(FE_OFN134_n_27449), .o(n_23135) );
oa22f80 g545824 ( .a(n_23334), .b(FE_OFN313_n_3069), .c(n_720), .d(FE_OFN131_n_27449), .o(n_24296) );
oa22f80 g545825 ( .a(n_21490), .b(FE_OFN297_n_3069), .c(n_392), .d(FE_OFN142_n_27449), .o(n_22552) );
oa22f80 g545826 ( .a(n_23627), .b(FE_OFN417_n_28303), .c(n_1614), .d(FE_OFN142_n_27449), .o(n_24605) );
oa22f80 g545827 ( .a(n_23332), .b(FE_OFN181_n_27681), .c(n_1184), .d(FE_OFN136_n_27449), .o(n_24295) );
oa22f80 g545828 ( .a(n_23626), .b(FE_OFN180_n_27681), .c(n_1710), .d(FE_OFN134_n_27449), .o(n_24604) );
oa22f80 g545829 ( .a(FE_OFN891_n_22165), .b(n_21988), .c(n_643), .d(n_28928), .o(n_23133) );
oa22f80 g545830 ( .a(n_23331), .b(n_29496), .c(n_25), .d(n_28928), .o(n_24294) );
oa22f80 g545831 ( .a(n_22164), .b(n_21988), .c(n_37), .d(FE_OFN1118_rst), .o(n_23132) );
oa22f80 g545832 ( .a(n_23625), .b(FE_OFN308_n_3069), .c(n_418), .d(FE_OFN114_n_27449), .o(n_24603) );
oa22f80 g545833 ( .a(n_23926), .b(FE_OFN295_n_3069), .c(n_345), .d(FE_OFN360_n_4860), .o(n_24920) );
oa22f80 g545834 ( .a(n_23330), .b(FE_OFN264_n_4280), .c(n_1341), .d(FE_OFN65_n_27012), .o(n_24293) );
oa22f80 g545835 ( .a(n_21936), .b(FE_OFN296_n_3069), .c(n_1477), .d(FE_OFN104_n_27449), .o(n_22250) );
oa22f80 g545836 ( .a(n_24020), .b(FE_OFN312_n_3069), .c(n_1166), .d(FE_OFN113_n_27449), .o(n_24021) );
oa22f80 g545837 ( .a(n_23329), .b(FE_OFN313_n_3069), .c(n_659), .d(FE_OFN142_n_27449), .o(n_24292) );
oa22f80 g545838 ( .a(n_21910), .b(FE_OFN414_n_28303), .c(n_825), .d(FE_OFN353_n_4860), .o(n_22849) );
oa22f80 g545839 ( .a(FE_OFN997_n_23622), .b(n_21988), .c(n_1631), .d(n_27449), .o(n_24601) );
oa22f80 g545840 ( .a(FE_OFN514_n_23620), .b(n_21988), .c(n_322), .d(n_27449), .o(n_24600) );
oa22f80 g545841 ( .a(n_21911), .b(FE_OFN413_n_28303), .c(n_1569), .d(FE_OFN138_n_27449), .o(n_22848) );
oa22f80 g545842 ( .a(n_23619), .b(FE_OFN413_n_28303), .c(n_687), .d(FE_OFN104_n_27449), .o(n_24598) );
oa22f80 g545843 ( .a(n_21909), .b(FE_OFN300_n_3069), .c(n_1955), .d(FE_OFN1110_rst), .o(n_22847) );
oa22f80 g545844 ( .a(n_23616), .b(FE_OFN184_n_29402), .c(n_820), .d(FE_OFN326_n_4860), .o(n_24596) );
oa22f80 g545845 ( .a(n_23130), .b(FE_OFN183_n_29402), .c(n_1526), .d(FE_OFN80_n_27012), .o(n_23131) );
oa22f80 g545846 ( .a(n_22162), .b(FE_OFN175_n_26184), .c(n_955), .d(FE_OFN75_n_27012), .o(n_23129) );
oa22f80 g545847 ( .a(n_23924), .b(FE_OFN148_n_25677), .c(n_1578), .d(FE_OFN105_n_27449), .o(n_24919) );
oa22f80 g545848 ( .a(n_21937), .b(FE_OFN150_n_25677), .c(n_1405), .d(FE_OFN326_n_4860), .o(n_22249) );
oa22f80 g545849 ( .a(n_22161), .b(FE_OFN402_n_28303), .c(n_31), .d(FE_OFN364_n_4860), .o(n_23128) );
oa22f80 g545850 ( .a(n_23923), .b(FE_OFN311_n_3069), .c(n_1596), .d(FE_OFN1123_rst), .o(n_24918) );
oa22f80 g545851 ( .a(n_21907), .b(FE_OFN410_n_28303), .c(n_1272), .d(FE_OFN135_n_27449), .o(n_22846) );
oa22f80 g545852 ( .a(n_23328), .b(FE_OFN183_n_29402), .c(n_693), .d(FE_OFN130_n_27449), .o(n_24291) );
oa22f80 g545853 ( .a(n_23615), .b(n_4280), .c(n_1386), .d(FE_OFN105_n_27449), .o(n_24595) );
oa22f80 g545854 ( .a(n_23327), .b(FE_OFN310_n_3069), .c(n_1249), .d(FE_OFN134_n_27449), .o(n_24290) );
oa22f80 g545855 ( .a(n_22432), .b(FE_OFN256_n_4280), .c(n_266), .d(FE_OFN1123_rst), .o(n_23408) );
ao22s80 g545856 ( .a(n_24019), .b(x_in_4_12), .c(n_23656), .d(n_16444), .o(n_24670) );
na02f80 g545933 ( .a(n_23690), .b(n_23956), .o(n_23691) );
no02f80 g545934 ( .a(n_23695), .b(n_23405), .o(n_23406) );
na02f80 g545935 ( .a(n_23096), .b(x_in_60_8), .o(n_24035) );
no02f80 g545936 ( .a(n_24288), .b(n_24287), .o(n_24289) );
no02f80 g545937 ( .a(n_24285), .b(n_24284), .o(n_24286) );
no02f80 g545938 ( .a(n_22263), .b(n_21974), .o(n_21975) );
in01f80 g545939 ( .a(n_22844), .o(n_22845) );
no02f80 g545940 ( .a(n_22551), .b(x_in_2_8), .o(n_22844) );
in01f80 g545941 ( .a(n_23126), .o(n_23127) );
no02f80 g545942 ( .a(n_22824), .b(x_in_40_8), .o(n_23126) );
na02f80 g545943 ( .a(n_22551), .b(x_in_2_8), .o(n_23451) );
no02f80 g545944 ( .a(n_24282), .b(n_24281), .o(n_24283) );
in01f80 g545945 ( .a(n_23124), .o(n_23125) );
no02f80 g545946 ( .a(n_22843), .b(x_in_34_8), .o(n_23124) );
na02f80 g545947 ( .a(n_22843), .b(x_in_34_8), .o(n_23710) );
no02f80 g545948 ( .a(n_24592), .b(n_24591), .o(n_24593) );
no02f80 g545949 ( .a(n_24279), .b(n_24278), .o(n_24280) );
no02f80 g545950 ( .a(n_24017), .b(n_24016), .o(n_24018) );
na02f80 g545951 ( .a(n_24015), .b(x_in_8_11), .o(n_24982) );
in01f80 g545952 ( .a(n_24276), .o(n_24277) );
no02f80 g545953 ( .a(n_24015), .b(x_in_8_11), .o(n_24276) );
no02f80 g545954 ( .a(n_22563), .b(n_22247), .o(n_22248) );
in01f80 g545955 ( .a(n_23122), .o(n_23123) );
no02f80 g545956 ( .a(n_22842), .b(x_in_18_8), .o(n_23122) );
na02f80 g545957 ( .a(n_22842), .b(x_in_18_8), .o(n_23709) );
no02f80 g545958 ( .a(n_23134), .b(n_22840), .o(n_22841) );
no02f80 g545959 ( .a(n_22166), .b(n_22840), .o(n_23799) );
no02f80 g545960 ( .a(n_24274), .b(n_24273), .o(n_24275) );
in01f80 g545961 ( .a(n_23120), .o(n_23121) );
no02f80 g545962 ( .a(n_22839), .b(x_in_50_8), .o(n_23120) );
na02f80 g545963 ( .a(n_22839), .b(x_in_50_8), .o(n_23704) );
in01f80 g545964 ( .a(n_23118), .o(n_23119) );
na02f80 g545965 ( .a(n_22838), .b(x_in_6_8), .o(n_23118) );
no02f80 g545966 ( .a(n_22838), .b(x_in_6_8), .o(n_23708) );
no02f80 g545967 ( .a(n_24271), .b(n_24270), .o(n_24272) );
in01f80 g545968 ( .a(n_22836), .o(n_22837) );
no02f80 g545969 ( .a(n_22550), .b(x_in_10_8), .o(n_22836) );
na02f80 g545970 ( .a(n_22550), .b(x_in_10_8), .o(n_23448) );
no02f80 g545971 ( .a(n_24013), .b(n_24012), .o(n_24014) );
in01f80 g545972 ( .a(n_22834), .o(n_22835) );
no02f80 g545973 ( .a(n_22549), .b(x_in_42_8), .o(n_22834) );
na02f80 g545974 ( .a(n_22549), .b(x_in_42_8), .o(n_23447) );
in01f80 g545975 ( .a(n_22832), .o(n_22833) );
no02f80 g545976 ( .a(n_22548), .b(x_in_26_8), .o(n_22832) );
na02f80 g545977 ( .a(n_22564), .b(n_22245), .o(n_22246) );
na02f80 g545978 ( .a(n_22548), .b(x_in_26_8), .o(n_23446) );
no02f80 g545979 ( .a(n_24268), .b(n_24572), .o(n_24269) );
no02f80 g545980 ( .a(n_24010), .b(n_24009), .o(n_24011) );
in01f80 g545981 ( .a(n_23116), .o(n_23117) );
no02f80 g545982 ( .a(n_22831), .b(x_in_58_8), .o(n_23116) );
no02f80 g545983 ( .a(n_24266), .b(n_24265), .o(n_24267) );
na02f80 g545984 ( .a(n_22831), .b(x_in_58_8), .o(n_23707) );
na02f80 g545985 ( .a(n_23993), .b(x_in_56_10), .o(n_24981) );
in01f80 g545986 ( .a(n_23403), .o(n_23404) );
na02f80 g545987 ( .a(n_23115), .b(n_22455), .o(n_23403) );
no02f80 g545988 ( .a(n_24007), .b(n_24218), .o(n_24008) );
no02f80 g545989 ( .a(n_24005), .b(n_24004), .o(n_24006) );
in01f80 g545990 ( .a(n_23401), .o(n_23402) );
na02f80 g545991 ( .a(n_23114), .b(n_22463), .o(n_23401) );
na02f80 g545992 ( .a(n_22562), .b(n_22243), .o(n_22244) );
na02f80 g545993 ( .a(n_22830), .b(x_in_22_8), .o(n_23701) );
in01f80 g545994 ( .a(n_23112), .o(n_23113) );
no02f80 g545995 ( .a(n_22830), .b(x_in_22_8), .o(n_23112) );
na02f80 g545996 ( .a(n_22547), .b(x_in_2_9), .o(n_23439) );
in01f80 g545997 ( .a(n_22828), .o(n_22829) );
no02f80 g545998 ( .a(n_22547), .b(x_in_2_9), .o(n_22828) );
in01f80 g545999 ( .a(n_22545), .o(n_22546) );
na02f80 g546000 ( .a(n_22242), .b(x_in_52_8), .o(n_22545) );
no02f80 g546001 ( .a(n_21978), .b(n_21569), .o(n_21570) );
no02f80 g546002 ( .a(n_22242), .b(x_in_52_8), .o(n_23160) );
na02f80 g546003 ( .a(n_22544), .b(x_in_54_8), .o(n_23445) );
in01f80 g546004 ( .a(n_22826), .o(n_22827) );
no02f80 g546005 ( .a(n_22544), .b(x_in_54_8), .o(n_22826) );
na02f80 g546006 ( .a(n_22825), .b(x_in_22_9), .o(n_23706) );
in01f80 g546007 ( .a(n_23110), .o(n_23111) );
no02f80 g546008 ( .a(n_22825), .b(x_in_22_9), .o(n_23110) );
no02f80 g546009 ( .a(n_24002), .b(n_24001), .o(n_24003) );
na02f80 g546010 ( .a(n_22824), .b(x_in_40_8), .o(n_23711) );
no02f80 g546011 ( .a(n_24263), .b(n_24262), .o(n_24264) );
no02f80 g546012 ( .a(n_22543), .b(x_in_14_8), .o(n_23449) );
in01f80 g546013 ( .a(n_22822), .o(n_22823) );
na02f80 g546014 ( .a(n_22543), .b(x_in_14_8), .o(n_22822) );
na02f80 g546015 ( .a(n_22542), .b(x_in_46_8), .o(n_23442) );
na02f80 g546016 ( .a(n_22269), .b(n_21972), .o(n_21973) );
in01f80 g546017 ( .a(n_22820), .o(n_22821) );
no02f80 g546018 ( .a(n_22542), .b(x_in_46_8), .o(n_22820) );
no02f80 g546019 ( .a(n_23999), .b(n_23998), .o(n_24000) );
in01f80 g546020 ( .a(n_22818), .o(n_22819) );
no02f80 g546021 ( .a(n_22532), .b(x_in_30_8), .o(n_22818) );
na02f80 g546022 ( .a(n_22541), .b(x_in_54_9), .o(n_23440) );
in01f80 g546023 ( .a(n_22816), .o(n_22817) );
no02f80 g546024 ( .a(n_22541), .b(x_in_54_9), .o(n_22816) );
no02f80 g546025 ( .a(n_23996), .b(n_23995), .o(n_23997) );
na02f80 g546026 ( .a(n_22540), .b(x_in_62_8), .o(n_23441) );
in01f80 g546027 ( .a(n_22814), .o(n_22815) );
no02f80 g546028 ( .a(n_22540), .b(x_in_62_8), .o(n_22814) );
in01f80 g546029 ( .a(n_24260), .o(n_24261) );
na02f80 g546030 ( .a(n_23994), .b(n_23366), .o(n_24260) );
in01f80 g546031 ( .a(n_24258), .o(n_24259) );
no02f80 g546032 ( .a(n_23993), .b(x_in_56_10), .o(n_24258) );
no02f80 g546033 ( .a(n_23991), .b(n_23990), .o(n_23992) );
no02f80 g546034 ( .a(n_24256), .b(n_24255), .o(n_24257) );
no02f80 g546035 ( .a(n_24253), .b(n_24252), .o(n_24254) );
no02f80 g546036 ( .a(n_23400), .b(x_in_36_8), .o(n_24322) );
na02f80 g546037 ( .a(n_22539), .b(x_in_14_9), .o(n_23438) );
in01f80 g546038 ( .a(n_22812), .o(n_22813) );
no02f80 g546039 ( .a(n_22539), .b(x_in_14_9), .o(n_22812) );
na02f80 g546040 ( .a(n_22811), .b(x_in_34_9), .o(n_23705) );
in01f80 g546041 ( .a(n_23108), .o(n_23109) );
no02f80 g546042 ( .a(n_22811), .b(x_in_34_9), .o(n_23108) );
na02f80 g546043 ( .a(n_22267), .b(n_21970), .o(n_21971) );
na02f80 g546044 ( .a(n_22538), .b(x_in_46_9), .o(n_23437) );
in01f80 g546045 ( .a(n_22809), .o(n_22810) );
no02f80 g546046 ( .a(n_22538), .b(x_in_46_9), .o(n_22809) );
no02f80 g546047 ( .a(n_24250), .b(n_24249), .o(n_24251) );
no02f80 g546048 ( .a(n_22266), .b(n_21968), .o(n_21969) );
na02f80 g546049 ( .a(n_22537), .b(x_in_16_9), .o(n_23436) );
in01f80 g546050 ( .a(n_22807), .o(n_22808) );
no02f80 g546051 ( .a(n_22537), .b(x_in_16_9), .o(n_22807) );
no02f80 g546052 ( .a(n_23988), .b(n_23987), .o(n_23989) );
no02f80 g546053 ( .a(n_24219), .b(n_23985), .o(n_23986) );
no02f80 g546054 ( .a(n_24916), .b(n_24915), .o(n_24917) );
no02f80 g546055 ( .a(n_23983), .b(n_23982), .o(n_23984) );
na02f80 g546056 ( .a(n_22265), .b(n_21966), .o(n_21967) );
na02f80 g546057 ( .a(n_22536), .b(x_in_30_9), .o(n_23435) );
in01f80 g546058 ( .a(n_22805), .o(n_22806) );
no02f80 g546059 ( .a(n_22536), .b(x_in_30_9), .o(n_22805) );
na02f80 g546060 ( .a(n_22535), .b(x_in_18_9), .o(n_23433) );
in01f80 g546061 ( .a(n_22803), .o(n_22804) );
no02f80 g546062 ( .a(n_22535), .b(x_in_18_9), .o(n_22803) );
no02f80 g546063 ( .a(n_24247), .b(n_24246), .o(n_24248) );
na02f80 g546064 ( .a(n_22264), .b(n_21964), .o(n_21965) );
na02f80 g546065 ( .a(n_22802), .b(x_in_12_9), .o(n_23702) );
in01f80 g546066 ( .a(n_23106), .o(n_23107) );
no02f80 g546067 ( .a(n_22802), .b(x_in_12_9), .o(n_23106) );
na02f80 g546068 ( .a(n_22534), .b(x_in_62_9), .o(n_23434) );
in01f80 g546069 ( .a(n_22800), .o(n_22801) );
no02f80 g546070 ( .a(n_22534), .b(x_in_62_9), .o(n_22800) );
no02f80 g546071 ( .a(n_24244), .b(n_24243), .o(n_24245) );
no02f80 g546072 ( .a(n_23980), .b(n_23979), .o(n_23981) );
no02f80 g546073 ( .a(n_23688), .b(n_23687), .o(n_23689) );
in01f80 g546074 ( .a(n_23104), .o(n_23105) );
no02f80 g546075 ( .a(n_22799), .b(x_in_16_8), .o(n_23104) );
na02f80 g546076 ( .a(n_22799), .b(x_in_16_8), .o(n_23703) );
in01f80 g546077 ( .a(n_23685), .o(n_23686) );
na02f80 g546078 ( .a(n_23400), .b(x_in_36_8), .o(n_23685) );
na02f80 g546079 ( .a(n_22533), .b(x_in_50_9), .o(n_23430) );
no02f80 g546080 ( .a(n_23683), .b(n_23682), .o(n_23684) );
in01f80 g546081 ( .a(n_22797), .o(n_22798) );
no02f80 g546082 ( .a(n_22533), .b(x_in_50_9), .o(n_22797) );
na02f80 g546083 ( .a(n_23399), .b(x_in_48_7), .o(n_24321) );
in01f80 g546084 ( .a(n_23680), .o(n_23681) );
no02f80 g546085 ( .a(n_23399), .b(x_in_48_7), .o(n_23680) );
no02f80 g546086 ( .a(n_24589), .b(n_24900), .o(n_24590) );
na02f80 g546087 ( .a(n_23679), .b(x_in_8_10), .o(n_24660) );
in01f80 g546088 ( .a(n_23977), .o(n_23978) );
no02f80 g546089 ( .a(n_23679), .b(x_in_8_10), .o(n_23977) );
no02f80 g546090 ( .a(n_22561), .b(n_22240), .o(n_22241) );
na02f80 g546091 ( .a(n_22532), .b(x_in_30_8), .o(n_23452) );
no02f80 g546092 ( .a(n_24241), .b(n_24240), .o(n_24242) );
na02f80 g546093 ( .a(n_23103), .b(x_in_40_7), .o(n_24031) );
in01f80 g546094 ( .a(n_23397), .o(n_23398) );
no02f80 g546095 ( .a(n_23103), .b(x_in_40_7), .o(n_23397) );
in01f80 g546096 ( .a(n_24238), .o(n_24239) );
na02f80 g546097 ( .a(n_23976), .b(n_23358), .o(n_24238) );
in01f80 g546098 ( .a(n_22795), .o(n_22796) );
na02f80 g546099 ( .a(n_22531), .b(x_in_32_8), .o(n_22795) );
no02f80 g546100 ( .a(n_22531), .b(x_in_32_8), .o(n_23429) );
na02f80 g546101 ( .a(n_23975), .b(x_in_44_11), .o(n_24978) );
no02f80 g546102 ( .a(n_23395), .b(n_23394), .o(n_23396) );
in01f80 g546103 ( .a(n_24236), .o(n_24237) );
no02f80 g546104 ( .a(n_23975), .b(x_in_44_11), .o(n_24236) );
in01f80 g546105 ( .a(n_23973), .o(n_23974) );
na02f80 g546106 ( .a(n_23678), .b(n_23067), .o(n_23973) );
na02f80 g546107 ( .a(n_23677), .b(x_in_24_12), .o(n_24659) );
in01f80 g546108 ( .a(n_23971), .o(n_23972) );
no02f80 g546109 ( .a(n_23677), .b(x_in_24_12), .o(n_23971) );
no02f80 g546110 ( .a(n_23969), .b(n_24215), .o(n_23970) );
na02f80 g546111 ( .a(n_23676), .b(x_in_56_9), .o(n_24657) );
in01f80 g546112 ( .a(n_23967), .o(n_23968) );
no02f80 g546113 ( .a(n_23676), .b(x_in_56_9), .o(n_23967) );
no02f80 g546114 ( .a(n_24026), .b(n_23674), .o(n_23675) );
na02f80 g546115 ( .a(n_22530), .b(x_in_10_9), .o(n_23428) );
in01f80 g546116 ( .a(n_22793), .o(n_22794) );
no02f80 g546117 ( .a(n_22530), .b(x_in_10_9), .o(n_22793) );
no02f80 g546118 ( .a(n_23147), .b(n_22791), .o(n_22792) );
na02f80 g546119 ( .a(n_23393), .b(x_in_20_8), .o(n_24323) );
in01f80 g546120 ( .a(n_23672), .o(n_23673) );
no02f80 g546121 ( .a(n_23393), .b(x_in_20_8), .o(n_23672) );
na02f80 g546122 ( .a(n_22268), .b(n_21962), .o(n_21963) );
na02f80 g546123 ( .a(n_23102), .b(x_in_48_8), .o(n_24028) );
in01f80 g546124 ( .a(n_23391), .o(n_23392) );
no02f80 g546125 ( .a(n_23102), .b(x_in_48_8), .o(n_23391) );
no02f80 g546126 ( .a(n_24234), .b(n_24233), .o(n_24235) );
in01f80 g546127 ( .a(n_23100), .o(n_23101) );
na02f80 g546128 ( .a(n_22790), .b(n_22180), .o(n_23100) );
no02f80 g546129 ( .a(n_23965), .b(n_23964), .o(n_23966) );
na02f80 g546130 ( .a(n_22529), .b(x_in_42_9), .o(n_23425) );
in01f80 g546131 ( .a(n_22788), .o(n_22789) );
no02f80 g546132 ( .a(n_22529), .b(x_in_42_9), .o(n_22788) );
no02f80 g546133 ( .a(n_23146), .b(n_22786), .o(n_22787) );
no02f80 g546134 ( .a(n_24231), .b(n_24230), .o(n_24232) );
no02f80 g546135 ( .a(n_22850), .b(n_22527), .o(n_22528) );
no02f80 g546136 ( .a(n_22262), .b(n_21960), .o(n_21961) );
no02f80 g546137 ( .a(n_21908), .b(n_22527), .o(n_23510) );
no02f80 g546138 ( .a(n_24587), .b(n_24586), .o(n_24588) );
na02f80 g546139 ( .a(n_23671), .b(x_in_20_7), .o(n_24656) );
in01f80 g546140 ( .a(n_23962), .o(n_23963) );
no02f80 g546141 ( .a(n_23671), .b(x_in_20_7), .o(n_23962) );
in01f80 g546142 ( .a(n_22784), .o(n_22785) );
no02f80 g546143 ( .a(n_22526), .b(x_in_26_9), .o(n_22784) );
na02f80 g546144 ( .a(n_22526), .b(x_in_26_9), .o(n_23424) );
no02f80 g546145 ( .a(n_22853), .b(n_22524), .o(n_22525) );
no02f80 g546146 ( .a(n_21912), .b(n_22524), .o(n_23506) );
no02f80 g546147 ( .a(n_24584), .b(n_24583), .o(n_24585) );
no02f80 g546148 ( .a(n_23960), .b(n_23959), .o(n_23961) );
no02f80 g546149 ( .a(n_23389), .b(n_23388), .o(n_23390) );
no02f80 g546150 ( .a(n_22783), .b(x_in_12_8), .o(n_23700) );
in01f80 g546151 ( .a(n_23098), .o(n_23099) );
na02f80 g546152 ( .a(n_22783), .b(x_in_12_8), .o(n_23098) );
no02f80 g546153 ( .a(n_24228), .b(n_24227), .o(n_24229) );
no02f80 g546154 ( .a(n_22261), .b(n_21958), .o(n_21959) );
no02f80 g546155 ( .a(n_20875), .b(FE_OFN369_n_26312), .o(n_21192) );
no02f80 g546156 ( .a(n_23957), .b(n_24212), .o(n_23958) );
in01f80 g546157 ( .a(n_24581), .o(n_24582) );
na02f80 g546158 ( .a(n_24226), .b(n_23642), .o(n_24581) );
in01f80 g546159 ( .a(n_23386), .o(n_23387) );
na02f80 g546160 ( .a(n_23097), .b(n_22440), .o(n_23386) );
na02f80 g546161 ( .a(n_22523), .b(x_in_58_9), .o(n_23450) );
in01f80 g546162 ( .a(n_22781), .o(n_22782) );
no02f80 g546163 ( .a(n_22523), .b(x_in_58_9), .o(n_22781) );
in01f80 g546164 ( .a(n_23384), .o(n_23385) );
no02f80 g546165 ( .a(n_23096), .b(x_in_60_8), .o(n_23384) );
na02f80 g546166 ( .a(n_23095), .b(x_in_60_7), .o(n_24036) );
in01f80 g546167 ( .a(n_23382), .o(n_23383) );
no02f80 g546168 ( .a(n_23095), .b(x_in_60_7), .o(n_23382) );
na02f80 g546169 ( .a(n_22560), .b(n_22238), .o(n_22239) );
na02f80 g546170 ( .a(n_21977), .b(n_21567), .o(n_21568) );
no02f80 g546171 ( .a(n_22260), .b(n_21956), .o(n_21957) );
na02f80 g546172 ( .a(n_23343), .b(n_23956), .o(n_24990) );
no02f80 g546173 ( .a(n_22867), .b(n_22521), .o(n_22522) );
no02f80 g546174 ( .a(n_22559), .b(n_22236), .o(n_22237) );
na02f80 g546175 ( .a(n_22259), .b(n_21954), .o(n_21955) );
no02f80 g546176 ( .a(n_23145), .b(n_22779), .o(n_22780) );
no02f80 g546177 ( .a(n_22258), .b(n_21952), .o(n_21953) );
no02f80 g546178 ( .a(n_22558), .b(n_22234), .o(n_22235) );
na02f80 g546179 ( .a(n_21976), .b(n_21565), .o(n_21566) );
na02f80 g546180 ( .a(n_22519), .b(n_22778), .o(n_22520) );
na02f80 g546181 ( .a(n_22232), .b(n_22518), .o(n_22233) );
no02f80 g546182 ( .a(n_22541), .b(n_22518), .o(n_23499) );
na02f80 g546183 ( .a(n_22230), .b(n_22515), .o(n_22231) );
na02f80 g546184 ( .a(n_22228), .b(n_22514), .o(n_22229) );
na02f80 g546185 ( .a(n_22226), .b(n_22517), .o(n_22227) );
no02f80 g546186 ( .a(n_22536), .b(n_22517), .o(n_23495) );
na02f80 g546187 ( .a(n_22224), .b(n_22516), .o(n_22225) );
no02f80 g546188 ( .a(n_22534), .b(n_22516), .o(n_23496) );
no02f80 g546189 ( .a(n_22825), .b(n_22778), .o(n_23740) );
no02f80 g546190 ( .a(n_22538), .b(n_22515), .o(n_23497) );
no02f80 g546191 ( .a(n_22539), .b(n_22514), .o(n_23498) );
na02f80 g546192 ( .a(n_22512), .b(n_22777), .o(n_22513) );
no02f80 g546193 ( .a(n_22802), .b(n_22777), .o(n_23739) );
no02f80 g546194 ( .a(n_22866), .b(n_22510), .o(n_22511) );
no02f80 g546195 ( .a(n_22257), .b(n_21950), .o(n_21951) );
no02f80 g546196 ( .a(n_22256), .b(n_21948), .o(n_21949) );
no02f80 g546197 ( .a(n_23692), .b(n_23380), .o(n_23381) );
no02f80 g546198 ( .a(FE_OFN753_n_22913), .b(n_23380), .o(n_24332) );
na02f80 g546199 ( .a(n_22509), .b(n_22508), .o(n_23418) );
in01f80 g546200 ( .a(n_22775), .o(n_22776) );
no02f80 g546201 ( .a(n_22509), .b(n_22508), .o(n_22775) );
na02f80 g546202 ( .a(n_24311), .b(x_in_36_7), .o(n_23670) );
na02f80 g546203 ( .a(n_22223), .b(n_22222), .o(n_23151) );
in01f80 g546204 ( .a(n_22506), .o(n_22507) );
no02f80 g546205 ( .a(n_22223), .b(n_22222), .o(n_22506) );
na02f80 g546206 ( .a(n_23954), .b(n_24020), .o(n_23955) );
no02f80 g546207 ( .a(n_23954), .b(n_23975), .o(n_24997) );
na02f80 g546208 ( .a(n_23694), .b(x_in_6_7), .o(n_23094) );
no02f80 g546209 ( .a(n_22557), .b(n_22220), .o(n_22221) );
no02f80 g546210 ( .a(n_22255), .b(n_21946), .o(n_21947) );
no02f80 g546211 ( .a(n_22254), .b(n_21944), .o(n_21945) );
no02f80 g546212 ( .a(n_22253), .b(n_21942), .o(n_21943) );
no02f80 g546213 ( .a(n_22251), .b(n_21940), .o(n_21941) );
no02f80 g546214 ( .a(n_23130), .b(n_22773), .o(n_22774) );
no02f80 g546215 ( .a(n_22163), .b(n_22773), .o(n_23736) );
na02f80 g546216 ( .a(n_22252), .b(n_21938), .o(n_21939) );
no02f80 g546217 ( .a(n_22218), .b(n_22217), .o(n_22219) );
na02f80 g546218 ( .a(n_21937), .b(n_22217), .o(n_23188) );
na02f80 g546219 ( .a(n_23668), .b(n_23953), .o(n_23669) );
no02f80 g546220 ( .a(n_24015), .b(n_23953), .o(n_25298) );
na02f80 g546221 ( .a(n_23945), .b(n_23944), .o(n_23952) );
no02f80 g546222 ( .a(n_23950), .b(n_24225), .o(n_23951) );
no02f80 g546223 ( .a(n_23948), .b(n_24224), .o(n_23949) );
no02f80 g546224 ( .a(n_22771), .b(n_22770), .o(n_22772) );
in01f80 g546225 ( .a(n_22769), .o(n_23486) );
na02f80 g546226 ( .a(n_22505), .b(n_22770), .o(n_22769) );
na02f80 g546227 ( .a(n_22503), .b(n_21832), .o(n_23485) );
na02f80 g546228 ( .a(n_22503), .b(n_22502), .o(n_22504) );
na02f80 g546229 ( .a(n_22767), .b(n_22120), .o(n_23734) );
na02f80 g546230 ( .a(n_22767), .b(n_22766), .o(n_22768) );
in01f80 g546231 ( .a(n_22765), .o(n_23480) );
no02f80 g546232 ( .a(n_22535), .b(n_22501), .o(n_22765) );
na02f80 g546233 ( .a(n_22215), .b(n_22501), .o(n_22216) );
na02f80 g546234 ( .a(n_22213), .b(n_22500), .o(n_22214) );
in01f80 g546235 ( .a(n_22764), .o(n_23477) );
no02f80 g546236 ( .a(n_22533), .b(n_22500), .o(n_22764) );
no02f80 g546237 ( .a(n_22498), .b(n_22497), .o(n_22499) );
no02f80 g546238 ( .a(n_22498), .b(n_21827), .o(n_23731) );
na02f80 g546239 ( .a(n_22495), .b(n_22494), .o(n_22496) );
na02f80 g546240 ( .a(n_22495), .b(n_21829), .o(n_23475) );
na02f80 g546241 ( .a(n_22492), .b(n_22491), .o(n_22493) );
na02f80 g546242 ( .a(n_22492), .b(n_21830), .o(n_23474) );
na02f80 g546243 ( .a(n_22489), .b(n_21828), .o(n_23473) );
na02f80 g546244 ( .a(n_22489), .b(n_22488), .o(n_22490) );
in01f80 g546245 ( .a(n_22763), .o(n_23470) );
no02f80 g546246 ( .a(n_22523), .b(n_22487), .o(n_22763) );
na02f80 g546247 ( .a(n_22211), .b(n_22487), .o(n_22212) );
na02f80 g546248 ( .a(n_22485), .b(n_22484), .o(n_22486) );
in01f80 g546249 ( .a(n_25016), .o(n_24580) );
oa12f80 g546250 ( .a(n_21526), .b(n_22189), .c(n_24225), .o(n_25016) );
ao12f80 g546251 ( .a(n_10825), .b(n_22210), .c(n_12060), .o(n_23169) );
in01f80 g546252 ( .a(n_25006), .o(n_24579) );
oa12f80 g546253 ( .a(n_21867), .b(n_22446), .c(n_24224), .o(n_25006) );
na02f80 g546254 ( .a(n_22483), .b(n_21820), .o(n_23467) );
na02f80 g546255 ( .a(n_22483), .b(n_22208), .o(n_22209) );
no02f80 g546256 ( .a(n_22206), .b(n_22205), .o(n_22207) );
in01f80 g546257 ( .a(n_22204), .o(n_22886) );
na02f80 g546258 ( .a(n_21936), .b(n_22205), .o(n_22204) );
in01f80 g546259 ( .a(n_22762), .o(n_23464) );
no02f80 g546260 ( .a(n_22537), .b(n_22482), .o(n_22762) );
na02f80 g546261 ( .a(n_22202), .b(n_22482), .o(n_22203) );
in01f80 g546262 ( .a(n_23379), .o(n_24048) );
no02f80 g546263 ( .a(n_23102), .b(n_23093), .o(n_23379) );
na02f80 g546264 ( .a(n_22760), .b(n_23093), .o(n_22761) );
no02f80 g546265 ( .a(n_22200), .b(n_22199), .o(n_22201) );
no02f80 g546266 ( .a(n_22200), .b(n_21466), .o(n_23461) );
na02f80 g546267 ( .a(n_22485), .b(n_21826), .o(n_23726) );
in01f80 g546268 ( .a(n_23092), .o(n_23722) );
no02f80 g546269 ( .a(n_22824), .b(n_22759), .o(n_23092) );
na02f80 g546270 ( .a(n_22480), .b(n_22759), .o(n_22481) );
na02f80 g546271 ( .a(n_23666), .b(n_23665), .o(n_23667) );
na02f80 g546272 ( .a(n_23666), .b(n_22976), .o(n_25294) );
no02f80 g546273 ( .a(n_22478), .b(n_22477), .o(n_22479) );
in01f80 g546274 ( .a(n_22476), .o(n_23174) );
na02f80 g546275 ( .a(n_22198), .b(n_22477), .o(n_22476) );
ao12f80 g546276 ( .a(n_16074), .b(n_23377), .c(n_23376), .o(n_23378) );
na02f80 g546277 ( .a(n_23091), .b(n_22392), .o(n_24331) );
na02f80 g546278 ( .a(n_23091), .b(n_23089), .o(n_23090) );
in01f80 g546279 ( .a(n_23664), .o(n_24328) );
no02f80 g546280 ( .a(n_23393), .b(n_23375), .o(n_23664) );
na02f80 g546281 ( .a(n_23087), .b(n_23375), .o(n_23088) );
na02f80 g546282 ( .a(n_22197), .b(n_21461), .o(n_23173) );
na02f80 g546283 ( .a(n_22197), .b(n_21934), .o(n_21935) );
no02f80 g546284 ( .a(n_22474), .b(n_22473), .o(n_22475) );
in01f80 g546285 ( .a(n_22472), .o(n_23170) );
na02f80 g546286 ( .a(n_22196), .b(n_22473), .o(n_22472) );
na02f80 g546287 ( .a(n_23085), .b(n_22386), .o(n_24045) );
na02f80 g546288 ( .a(n_23085), .b(n_23084), .o(n_23086) );
in01f80 g546289 ( .a(n_25648), .o(n_25251) );
oa12f80 g546290 ( .a(n_22750), .b(n_22153), .c(n_23919), .o(n_25648) );
in01f80 g546291 ( .a(n_25645), .o(n_25250) );
oa12f80 g546292 ( .a(n_23065), .b(n_22425), .c(n_23918), .o(n_25645) );
in01f80 g546293 ( .a(n_25642), .o(n_25248) );
oa12f80 g546294 ( .a(n_22465), .b(n_21895), .c(n_23917), .o(n_25642) );
in01f80 g546295 ( .a(n_25639), .o(n_25247) );
oa12f80 g546296 ( .a(n_22456), .b(n_21890), .c(n_23916), .o(n_25639) );
in01f80 g546297 ( .a(n_25339), .o(n_24914) );
oa12f80 g546298 ( .a(n_22748), .b(n_23600), .c(n_22148), .o(n_25339) );
in01f80 g546299 ( .a(n_25336), .o(n_24913) );
oa12f80 g546300 ( .a(n_22747), .b(n_23599), .c(n_22146), .o(n_25336) );
in01f80 g546301 ( .a(n_25331), .o(n_24912) );
oa12f80 g546302 ( .a(n_22737), .b(n_23598), .c(n_22144), .o(n_25331) );
in01f80 g546303 ( .a(n_25347), .o(n_24911) );
oa12f80 g546304 ( .a(n_22464), .b(n_23597), .c(n_21874), .o(n_25347) );
in01f80 g546305 ( .a(n_24910), .o(n_25833) );
oa12f80 g546306 ( .a(n_21061), .b(n_24567), .c(n_20696), .o(n_24910) );
ao12f80 g546307 ( .a(n_24570), .b(n_22749), .c(n_24569), .o(n_25559) );
oa12f80 g546308 ( .a(n_12474), .b(n_21933), .c(n_13659), .o(n_22880) );
in01f80 g546309 ( .a(n_24578), .o(n_25557) );
oa12f80 g546310 ( .a(n_21398), .b(n_24220), .c(n_21002), .o(n_24578) );
in01f80 g546311 ( .a(n_25323), .o(n_24909) );
oa12f80 g546312 ( .a(n_22745), .b(n_22139), .c(n_23595), .o(n_25323) );
in01f80 g546313 ( .a(n_25609), .o(n_25246) );
oa12f80 g546314 ( .a(n_22457), .b(n_21847), .c(n_23915), .o(n_25609) );
in01f80 g546315 ( .a(n_25326), .o(n_24908) );
oa12f80 g546316 ( .a(n_22453), .b(n_21883), .c(n_23594), .o(n_25326) );
in01f80 g546317 ( .a(n_25623), .o(n_25245) );
oa12f80 g546318 ( .a(n_22460), .b(n_21881), .c(n_23913), .o(n_25623) );
in01f80 g546319 ( .a(n_25588), .o(n_25244) );
oa12f80 g546320 ( .a(n_22736), .b(n_22151), .c(n_23912), .o(n_25588) );
in01f80 g546321 ( .a(n_25317), .o(n_24907) );
oa12f80 g546322 ( .a(n_22461), .b(n_21845), .c(n_23593), .o(n_25317) );
in01f80 g546323 ( .a(n_25314), .o(n_24906) );
oa12f80 g546324 ( .a(n_22459), .b(n_21878), .c(n_23592), .o(n_25314) );
in01f80 g546325 ( .a(n_25614), .o(n_25243) );
oa12f80 g546326 ( .a(n_22190), .b(n_21530), .c(n_23914), .o(n_25614) );
in01f80 g546327 ( .a(n_25320), .o(n_24905) );
oa12f80 g546328 ( .a(n_22458), .b(n_21876), .c(n_23591), .o(n_25320) );
in01f80 g546329 ( .a(n_24577), .o(n_25555) );
oa12f80 g546330 ( .a(n_20428), .b(n_24216), .c(n_20026), .o(n_24577) );
in01f80 g546331 ( .a(n_26095), .o(n_25798) );
oa12f80 g546332 ( .a(n_22744), .b(n_22137), .c(n_24528), .o(n_26095) );
in01f80 g546333 ( .a(n_25597), .o(n_25242) );
oa12f80 g546334 ( .a(n_22187), .b(n_21524), .c(n_23911), .o(n_25597) );
in01f80 g546335 ( .a(n_25311), .o(n_24904) );
oa12f80 g546336 ( .a(n_22452), .b(n_21871), .c(n_23590), .o(n_25311) );
in01f80 g546337 ( .a(n_25594), .o(n_25241) );
oa12f80 g546338 ( .a(n_22186), .b(n_21521), .c(n_23910), .o(n_25594) );
in01f80 g546339 ( .a(n_25308), .o(n_24903) );
oa12f80 g546340 ( .a(n_22451), .b(n_21869), .c(n_23589), .o(n_25308) );
in01f80 g546341 ( .a(n_25591), .o(n_25240) );
oa12f80 g546342 ( .a(n_22185), .b(n_21517), .c(n_23909), .o(n_25591) );
in01f80 g546343 ( .a(n_24223), .o(n_25287) );
oa12f80 g546344 ( .a(n_17696), .b(n_23942), .c(n_17055), .o(n_24223) );
oa12f80 g546345 ( .a(n_22743), .b(n_22135), .c(n_23271), .o(n_25290) );
in01f80 g546346 ( .a(n_25009), .o(n_24576) );
oa12f80 g546347 ( .a(n_22447), .b(n_21864), .c(n_23270), .o(n_25009) );
in01f80 g546348 ( .a(n_25585), .o(n_25239) );
oa12f80 g546349 ( .a(n_22445), .b(n_21862), .c(n_23908), .o(n_25585) );
in01f80 g546350 ( .a(n_23947), .o(n_24988) );
oa12f80 g546351 ( .a(n_3060), .b(n_23660), .c(n_2164), .o(n_23947) );
in01f80 g546352 ( .a(n_24902), .o(n_25831) );
oa12f80 g546353 ( .a(n_22042), .b(n_24565), .c(n_21629), .o(n_24902) );
in01f80 g546354 ( .a(n_24685), .o(n_24222) );
oa12f80 g546355 ( .a(n_22740), .b(n_22132), .c(n_22974), .o(n_24685) );
in01f80 g546356 ( .a(n_23946), .o(n_24986) );
oa12f80 g546357 ( .a(n_21430), .b(n_23658), .c(n_20748), .o(n_23946) );
oa12f80 g546358 ( .a(n_13124), .b(n_22195), .c(n_14267), .o(n_23168) );
in01f80 g546359 ( .a(n_25581), .o(n_25238) );
oa12f80 g546360 ( .a(n_22444), .b(n_23907), .c(n_21858), .o(n_25581) );
in01f80 g546361 ( .a(n_24575), .o(n_25553) );
oa12f80 g546362 ( .a(n_20737), .b(n_24213), .c(n_20340), .o(n_24575) );
in01f80 g546363 ( .a(n_25874), .o(n_25521) );
oa12f80 g546364 ( .a(n_23363), .b(n_22669), .c(n_24194), .o(n_25874) );
in01f80 g546365 ( .a(n_25578), .o(n_25237) );
oa12f80 g546366 ( .a(n_22443), .b(n_23906), .c(n_21854), .o(n_25578) );
ao12f80 g546367 ( .a(n_25230), .b(n_23643), .c(n_25229), .o(n_26050) );
in01f80 g546368 ( .a(n_25849), .o(n_25519) );
oa12f80 g546369 ( .a(n_23353), .b(n_22663), .c(n_24193), .o(n_25849) );
in01f80 g546370 ( .a(n_25575), .o(n_25236) );
oa12f80 g546371 ( .a(n_22441), .b(n_23905), .c(n_21849), .o(n_25575) );
oa12f80 g546372 ( .a(n_22442), .b(n_22973), .c(n_21843), .o(n_24991) );
in01f80 g546373 ( .a(n_24574), .o(n_25551) );
oa12f80 g546374 ( .a(n_22353), .b(n_24210), .c(n_21658), .o(n_24574) );
in01f80 g546375 ( .a(n_24573), .o(n_25549) );
oa12f80 g546376 ( .a(n_21348), .b(n_24208), .c(n_20991), .o(n_24573) );
in01f80 g546377 ( .a(n_25344), .o(n_24901) );
oa12f80 g546378 ( .a(n_22466), .b(n_23587), .c(n_21841), .o(n_25344) );
in01f80 g546379 ( .a(n_25636), .o(n_25235) );
oa12f80 g546380 ( .a(n_23074), .b(n_22407), .c(n_23904), .o(n_25636) );
in01f80 g546381 ( .a(n_25651), .o(n_25234) );
oa12f80 g546382 ( .a(n_23364), .b(n_22655), .c(n_23903), .o(n_25651) );
oa12f80 g546383 ( .a(n_12268), .b(n_21564), .c(n_12943), .o(n_22577) );
in01f80 g546384 ( .a(n_24030), .o(n_23663) );
oa12f80 g546385 ( .a(n_2546), .b(n_23374), .c(n_23075), .o(n_24030) );
oa12f80 g546386 ( .a(n_10841), .b(n_22194), .c(n_12064), .o(n_23166) );
ao12f80 g546387 ( .a(n_12705), .b(n_23083), .c(n_14021), .o(n_24044) );
oa12f80 g546388 ( .a(n_23945), .b(n_23376), .c(n_23944), .o(n_24992) );
ao12f80 g546389 ( .a(n_2097), .b(n_23373), .c(n_23345), .o(n_24033) );
ao12f80 g546390 ( .a(n_22652), .b(n_24900), .c(n_23349), .o(n_25844) );
ao12f80 g546391 ( .a(n_12497), .b(n_21932), .c(n_11532), .o(n_22574) );
oa12f80 g546392 ( .a(n_12936), .b(n_21931), .c(n_14085), .o(n_22885) );
ao12f80 g546393 ( .a(n_22437), .b(n_22752), .c(n_22436), .o(n_23082) );
in01f80 g546394 ( .a(n_22567), .o(n_22193) );
oa12f80 g546395 ( .a(n_21189), .b(n_21564), .c(n_21188), .o(n_22567) );
ao22s80 g546396 ( .a(n_23586), .b(n_22433), .c(n_24572), .d(x_in_6_7), .o(n_25566) );
ao12f80 g546397 ( .a(n_21919), .b(n_21918), .c(n_21917), .o(n_22471) );
oa12f80 g546398 ( .a(n_22746), .b(n_24570), .c(n_24569), .o(n_24571) );
in01f80 g546399 ( .a(n_22879), .o(n_22470) );
oa12f80 g546400 ( .a(n_21560), .b(n_21933), .c(n_21559), .o(n_22879) );
oa12f80 g546401 ( .a(n_21921), .b(n_21920), .c(n_22174), .o(n_23159) );
ao22s80 g546402 ( .a(n_21400), .b(n_24567), .c(n_21399), .d(n_23596), .o(n_24568) );
ao22s80 g546403 ( .a(n_21735), .b(n_24220), .c(n_21734), .d(n_23273), .o(n_24221) );
ao22s80 g546404 ( .a(n_23264), .b(n_21544), .c(n_24219), .d(x_in_52_7), .o(n_25296) );
ao22s80 g546405 ( .a(n_23259), .b(n_22591), .c(n_24218), .d(x_in_14_7), .o(n_25297) );
in01f80 g546406 ( .a(n_23152), .o(n_23420) );
ao12f80 g546407 ( .a(n_21929), .b(n_22194), .c(n_21928), .o(n_23152) );
ao22s80 g546408 ( .a(n_24216), .b(n_20756), .c(n_23272), .d(n_20755), .o(n_24217) );
ao12f80 g546409 ( .a(n_23073), .b(n_23373), .c(n_23072), .o(n_23662) );
in01f80 g546410 ( .a(n_22758), .o(n_23715) );
oa12f80 g546411 ( .a(n_21924), .b(n_22210), .c(n_21923), .o(n_22758) );
ao22s80 g546412 ( .a(n_23942), .b(n_17905), .c(n_22975), .d(n_17904), .o(n_23943) );
ao12f80 g546413 ( .a(n_22450), .b(n_22449), .c(n_22448), .o(n_23081) );
in01f80 g546414 ( .a(n_21563), .o(n_22270) );
ao12f80 g546415 ( .a(n_20473), .b(n_20474), .c(n_20472), .o(n_21563) );
ao22s80 g546416 ( .a(n_23660), .b(n_3707), .c(n_22650), .d(n_3706), .o(n_23661) );
ao12f80 g546417 ( .a(n_22735), .b(n_22734), .c(n_22733), .o(n_23372) );
in01f80 g546418 ( .a(n_23080), .o(n_24038) );
oa12f80 g546419 ( .a(n_22183), .b(n_22182), .c(n_22181), .o(n_23080) );
in01f80 g546420 ( .a(n_24054), .o(n_24337) );
ao12f80 g546421 ( .a(n_22742), .b(n_23083), .c(n_22741), .o(n_24054) );
ao22s80 g546422 ( .a(n_23256), .b(n_21900), .c(n_24215), .d(x_in_32_7), .o(n_25295) );
ao12f80 g546423 ( .a(n_22177), .b(n_22468), .c(n_22176), .o(n_22757) );
in01f80 g546424 ( .a(n_22874), .o(n_23155) );
ao12f80 g546425 ( .a(n_21556), .b(n_21932), .c(n_21555), .o(n_22874) );
oa12f80 g546426 ( .a(n_23351), .b(n_23374), .c(n_23350), .o(n_24658) );
ao12f80 g546427 ( .a(n_22173), .b(n_22172), .c(n_22171), .o(n_22756) );
in01f80 g546428 ( .a(n_23148), .o(n_23416) );
ao12f80 g546429 ( .a(n_21927), .b(n_22195), .c(n_21926), .o(n_23148) );
ao22s80 g546430 ( .a(n_24565), .b(n_22303), .c(n_23588), .d(n_22302), .o(n_24566) );
ao22s80 g546431 ( .a(n_21789), .b(n_23658), .c(n_21788), .d(n_22649), .o(n_23659) );
in01f80 g546432 ( .a(n_22870), .o(n_23158) );
ao12f80 g546433 ( .a(n_21558), .b(n_21931), .c(n_21557), .o(n_22870) );
ao22s80 g546434 ( .a(n_23377), .b(n_16655), .c(n_23656), .d(n_16654), .o(n_23657) );
oa12f80 g546435 ( .a(n_23644), .b(n_25230), .c(n_25229), .o(n_25231) );
ao22s80 g546436 ( .a(n_21034), .b(n_24213), .c(n_21033), .d(n_23269), .o(n_24214) );
ao22s80 g546437 ( .a(n_23251), .b(n_22731), .c(n_24212), .d(x_in_12_7), .o(n_25293) );
ao12f80 g546438 ( .a(n_20877), .b(n_21190), .c(n_20876), .o(n_21562) );
in01f80 g546439 ( .a(n_24316), .o(n_23941) );
oa12f80 g546440 ( .a(n_23063), .b(n_23348), .c(n_23070), .o(n_24316) );
ao22s80 g546441 ( .a(n_24210), .b(n_22632), .c(n_23268), .d(n_22631), .o(n_24211) );
oa12f80 g546442 ( .a(n_21922), .b(n_21925), .c(n_22175), .o(n_23157) );
ao22s80 g546443 ( .a(n_21657), .b(n_24208), .c(n_21656), .d(n_23267), .o(n_24209) );
oa22f80 g546444 ( .a(n_22115), .b(FE_OFN411_n_28303), .c(n_455), .d(FE_OFN192_n_28928), .o(n_23079) );
oa22f80 g546445 ( .a(n_21554), .b(FE_OFN267_n_4280), .c(n_245), .d(FE_OFN60_n_27012), .o(n_21930) );
oa22f80 g546446 ( .a(n_22438), .b(FE_OFN198_n_29637), .c(n_1156), .d(FE_OFN1112_rst), .o(n_22755) );
oa22f80 g546447 ( .a(n_21115), .b(FE_OFN199_n_29637), .c(n_1446), .d(FE_OFN92_n_27449), .o(n_22192) );
oa22f80 g546448 ( .a(FE_OFN1228_n_23261), .b(n_21988), .c(n_1692), .d(FE_OFN96_n_27449), .o(n_24207) );
oa22f80 g546449 ( .a(n_22972), .b(n_29698), .c(n_990), .d(FE_OFN336_n_4860), .o(n_23940) );
oa22f80 g546450 ( .a(n_22468), .b(n_21988), .c(n_1020), .d(FE_OFN347_n_4860), .o(n_22469) );
oa22f80 g546451 ( .a(n_21813), .b(FE_OFN409_n_28303), .c(n_1953), .d(FE_OFN355_n_4860), .o(n_22754) );
oa22f80 g546452 ( .a(n_22752), .b(FE_OFN411_n_28303), .c(n_1769), .d(FE_OFN364_n_4860), .o(n_22753) );
oa22f80 g546453 ( .a(n_22970), .b(FE_OFN314_n_3069), .c(n_508), .d(FE_OFN330_n_4860), .o(n_23939) );
oa22f80 g546454 ( .a(n_22384), .b(FE_OFN400_n_28303), .c(n_1304), .d(FE_OFN1114_rst), .o(n_23371) );
oa22f80 g546455 ( .a(n_22184), .b(FE_OFN294_n_3069), .c(n_792), .d(FE_OFN1119_rst), .o(n_22467) );
oa22f80 g546456 ( .a(n_22648), .b(FE_OFN295_n_3069), .c(n_1595), .d(FE_OFN15_n_29068), .o(n_23655) );
oa22f80 g546457 ( .a(n_22114), .b(FE_OFN253_n_4280), .c(n_218), .d(FE_OFN138_n_27449), .o(n_23078) );
oa22f80 g546458 ( .a(n_21190), .b(FE_OFN310_n_3069), .c(n_1857), .d(FE_OFN116_n_27449), .o(n_21191) );
oa22f80 g546459 ( .a(n_22382), .b(FE_OFN295_n_3069), .c(n_929), .d(FE_OFN76_n_27012), .o(n_23370) );
oa22f80 g546460 ( .a(n_22380), .b(FE_OFN307_n_3069), .c(n_1649), .d(FE_OFN1112_rst), .o(n_23369) );
oa22f80 g546461 ( .a(n_21814), .b(FE_OFN312_n_3069), .c(n_1271), .d(FE_OFN1106_rst), .o(n_22751) );
oa22f80 g546462 ( .a(n_22113), .b(FE_OFN306_n_3069), .c(n_1677), .d(rst), .o(n_23077) );
oa22f80 g546463 ( .a(n_23347), .b(FE_OFN312_n_3069), .c(n_1642), .d(FE_OFN1111_rst), .o(n_23653) );
oa22f80 g546464 ( .a(n_23253), .b(FE_OFN312_n_3069), .c(n_170), .d(FE_OFN330_n_4860), .o(n_24206) );
oa22f80 g546465 ( .a(n_22379), .b(FE_OFN186_n_29496), .c(n_54), .d(FE_OFN93_n_27449), .o(n_23367) );
oa22f80 g546466 ( .a(n_22646), .b(FE_OFN308_n_3069), .c(n_640), .d(FE_OFN114_n_27449), .o(n_23652) );
oa22f80 g546467 ( .a(FE_OFN686_n_22968), .b(FE_OFN292_n_3069), .c(n_398), .d(n_28607), .o(n_23938) );
oa22f80 g546468 ( .a(n_20464), .b(FE_OFN310_n_3069), .c(n_112), .d(FE_OFN353_n_4860), .o(n_21561) );
oa22f80 g546469 ( .a(n_22966), .b(FE_OFN412_n_28303), .c(n_1651), .d(FE_OFN113_n_27449), .o(n_23937) );
oa22f80 g546470 ( .a(n_22965), .b(FE_OFN312_n_3069), .c(n_73), .d(FE_OFN124_n_27449), .o(n_23936) );
oa22f80 g546471 ( .a(n_22963), .b(FE_OFN311_n_3069), .c(n_464), .d(FE_OFN80_n_27012), .o(n_23934) );
in01f80 g546501 ( .a(n_23365), .o(n_23366) );
no02f80 g546502 ( .a(n_23075), .b(x_in_24_13), .o(n_23365) );
na02f80 g546503 ( .a(n_23075), .b(x_in_24_13), .o(n_23994) );
na02f80 g546504 ( .a(n_23364), .b(n_22656), .o(n_24285) );
na02f80 g546505 ( .a(n_22750), .b(n_22154), .o(n_24282) );
na02f80 g546506 ( .a(n_23363), .b(n_22670), .o(n_24592) );
na02f80 g546507 ( .a(n_22466), .b(n_21842), .o(n_24017) );
na02f80 g546508 ( .a(n_22749), .b(n_22141), .o(n_24005) );
na02f80 g546509 ( .a(n_22465), .b(n_21896), .o(n_24274) );
na02f80 g546510 ( .a(n_22748), .b(n_22149), .o(n_24013) );
na02f80 g546511 ( .a(n_22747), .b(n_22147), .o(n_23965) );
na02f80 g546512 ( .a(n_23074), .b(n_22408), .o(n_24266) );
na02f80 g546513 ( .a(n_22464), .b(n_21875), .o(n_23991) );
na02f80 g546514 ( .a(n_22188), .b(x_in_38_11), .o(n_23115) );
no02f80 g546515 ( .a(n_22126), .b(x_in_6_7), .o(n_22746) );
na02f80 g546516 ( .a(n_21933), .b(n_21559), .o(n_21560) );
in01f80 g546517 ( .a(n_22462), .o(n_22463) );
no02f80 g546518 ( .a(n_22191), .b(x_in_38_10), .o(n_22462) );
na02f80 g546519 ( .a(n_22191), .b(x_in_38_10), .o(n_23114) );
na02f80 g546520 ( .a(n_22461), .b(n_21846), .o(n_23999) );
na02f80 g546521 ( .a(n_22460), .b(n_21882), .o(n_24288) );
na02f80 g546522 ( .a(n_22745), .b(n_22140), .o(n_23960) );
na02f80 g546523 ( .a(n_22459), .b(n_21879), .o(n_23996) );
in01f80 g546524 ( .a(n_23932), .o(n_23933) );
na02f80 g546525 ( .a(n_23651), .b(n_23017), .o(n_23932) );
na02f80 g546526 ( .a(n_22458), .b(n_21877), .o(n_23988) );
no02f80 g546527 ( .a(n_22194), .b(n_21928), .o(n_21929) );
in01f80 g546528 ( .a(n_23649), .o(n_23650) );
na02f80 g546529 ( .a(n_23362), .b(n_22730), .o(n_23649) );
na02f80 g546530 ( .a(n_22190), .b(n_21531), .o(n_24256) );
na02f80 g546531 ( .a(n_22457), .b(n_21848), .o(n_24253) );
no02f80 g546532 ( .a(n_23373), .b(n_23072), .o(n_23073) );
no02f80 g546533 ( .a(n_21527), .b(n_22189), .o(n_23950) );
na02f80 g546534 ( .a(n_22456), .b(n_21891), .o(n_24271) );
in01f80 g546535 ( .a(n_22454), .o(n_22455) );
no02f80 g546536 ( .a(n_22188), .b(x_in_38_11), .o(n_22454) );
na02f80 g546537 ( .a(n_22187), .b(n_21525), .o(n_24250) );
na02f80 g546538 ( .a(n_22453), .b(n_21884), .o(n_24002) );
na02f80 g546539 ( .a(n_22744), .b(n_22138), .o(n_24916) );
na02f80 g546540 ( .a(n_22452), .b(n_21872), .o(n_23983) );
na02f80 g546541 ( .a(n_22186), .b(n_21522), .o(n_24247) );
na02f80 g546542 ( .a(n_22185), .b(n_21518), .o(n_24244) );
na02f80 g546543 ( .a(n_22451), .b(n_21870), .o(n_23980) );
na02f80 g546544 ( .a(n_22743), .b(n_22136), .o(n_23688) );
no02f80 g546545 ( .a(n_22449), .b(n_22448), .o(n_22450) );
na02f80 g546546 ( .a(n_22184), .b(n_22448), .o(n_23431) );
na02f80 g546547 ( .a(n_22447), .b(n_21865), .o(n_23683) );
no02f80 g546548 ( .a(n_21868), .b(n_22446), .o(n_23948) );
in01f80 g546549 ( .a(n_23360), .o(n_23361) );
na02f80 g546550 ( .a(n_23071), .b(n_22424), .o(n_23360) );
na02f80 g546551 ( .a(n_22445), .b(n_21863), .o(n_24241) );
na02f80 g546552 ( .a(n_22182), .b(n_22181), .o(n_22183) );
no02f80 g546553 ( .a(n_23083), .b(n_22741), .o(n_22742) );
in01f80 g546554 ( .a(n_23647), .o(n_23648) );
na02f80 g546555 ( .a(n_23359), .b(n_22680), .o(n_23647) );
na02f80 g546556 ( .a(n_23070), .b(x_in_44_10), .o(n_23976) );
in01f80 g546557 ( .a(n_23357), .o(n_23358) );
no02f80 g546558 ( .a(n_23070), .b(x_in_44_10), .o(n_23357) );
na02f80 g546559 ( .a(n_22740), .b(n_22133), .o(n_23395) );
in01f80 g546560 ( .a(n_23068), .o(n_23069) );
na02f80 g546561 ( .a(n_22739), .b(n_22131), .o(n_23068) );
na02f80 g546562 ( .a(n_22738), .b(x_in_24_11), .o(n_23678) );
in01f80 g546563 ( .a(n_23066), .o(n_23067) );
no02f80 g546564 ( .a(n_22738), .b(x_in_24_11), .o(n_23066) );
no02f80 g546565 ( .a(n_22195), .b(n_21926), .o(n_21927) );
na02f80 g546566 ( .a(n_23065), .b(n_22426), .o(n_24279) );
na02f80 g546567 ( .a(n_22737), .b(n_22145), .o(n_24010) );
in01f80 g546568 ( .a(n_23645), .o(n_23646) );
na02f80 g546569 ( .a(n_23356), .b(n_22672), .o(n_23645) );
na02f80 g546570 ( .a(n_22444), .b(n_21859), .o(n_24234) );
na02f80 g546571 ( .a(n_21925), .b(x_in_28_11), .o(n_22790) );
in01f80 g546572 ( .a(n_23354), .o(n_23355) );
na02f80 g546573 ( .a(n_23064), .b(n_22414), .o(n_23354) );
in01f80 g546574 ( .a(n_22179), .o(n_22180) );
no02f80 g546575 ( .a(n_21925), .b(x_in_28_11), .o(n_22179) );
na02f80 g546576 ( .a(n_22736), .b(n_22152), .o(n_24263) );
no02f80 g546577 ( .a(n_22984), .b(x_in_36_7), .o(n_23644) );
na02f80 g546578 ( .a(n_22443), .b(n_21855), .o(n_24231) );
na02f80 g546579 ( .a(n_23643), .b(n_22983), .o(n_24587) );
na02f80 g546580 ( .a(n_23353), .b(n_22664), .o(n_24584) );
na02f80 g546581 ( .a(n_22442), .b(n_21844), .o(n_23389) );
na02f80 g546582 ( .a(n_22441), .b(n_21850), .o(n_24228) );
no02f80 g546583 ( .a(n_21190), .b(n_20876), .o(n_20877) );
in01f80 g546584 ( .a(n_20875), .o(n_22578) );
no02f80 g546585 ( .a(n_20107), .b(n_20876), .o(n_20875) );
na02f80 g546586 ( .a(n_23352), .b(x_in_44_9), .o(n_24226) );
in01f80 g546587 ( .a(n_23641), .o(n_23642) );
no02f80 g546588 ( .a(n_23352), .b(x_in_44_9), .o(n_23641) );
na02f80 g546589 ( .a(n_22178), .b(x_in_28_10), .o(n_23097) );
in01f80 g546590 ( .a(n_22439), .o(n_22440) );
no02f80 g546591 ( .a(n_22178), .b(x_in_28_10), .o(n_22439) );
na02f80 g546592 ( .a(n_22210), .b(n_21923), .o(n_21924) );
na02f80 g546593 ( .a(n_21564), .b(n_21188), .o(n_21189) );
na02f80 g546594 ( .a(n_20474), .b(n_9619), .o(n_20475) );
no02f80 g546595 ( .a(n_22734), .b(n_22733), .o(n_22735) );
na02f80 g546596 ( .a(n_22438), .b(n_22733), .o(n_23698) );
no02f80 g546597 ( .a(n_22468), .b(n_22176), .o(n_22177) );
no02f80 g546598 ( .a(n_21457), .b(n_22176), .o(n_23154) );
no02f80 g546599 ( .a(n_20474), .b(n_20472), .o(n_20473) );
no02f80 g546600 ( .a(n_22752), .b(n_22436), .o(n_22437) );
no02f80 g546601 ( .a(n_21812), .b(n_22436), .o(n_23419) );
na02f80 g546602 ( .a(n_23374), .b(n_23350), .o(n_23351) );
na02f80 g546603 ( .a(n_22653), .b(n_23349), .o(n_24589) );
na02f80 g546604 ( .a(n_23348), .b(n_23070), .o(n_23063) );
na02f80 g546605 ( .a(n_23348), .b(n_23347), .o(n_23954) );
na02f80 g546606 ( .a(n_21925), .b(n_22175), .o(n_21922) );
na02f80 g546607 ( .a(n_21456), .b(n_22175), .o(n_23150) );
no02f80 g546608 ( .a(n_21931), .b(n_21557), .o(n_21558) );
no02f80 g546609 ( .a(n_22188), .b(n_22174), .o(n_23149) );
na02f80 g546610 ( .a(n_21920), .b(n_22174), .o(n_21921) );
in01f80 g546611 ( .a(n_24019), .o(n_23346) );
na02f80 g546612 ( .a(n_23377), .b(n_23062), .o(n_24019) );
no02f80 g546613 ( .a(n_21932), .b(n_21555), .o(n_21556) );
no02f80 g546614 ( .a(n_21918), .b(n_21917), .o(n_21919) );
in01f80 g546615 ( .a(n_21916), .o(n_22565) );
na02f80 g546616 ( .a(n_21554), .b(n_21917), .o(n_21916) );
na03f80 g546617 ( .a(n_23345), .b(n_23373), .c(n_2210), .o(n_23945) );
oa12f80 g546618 ( .a(n_12343), .b(n_22732), .c(n_12342), .o(n_23695) );
no02f80 g546619 ( .a(n_22172), .b(n_22171), .o(n_22173) );
no02f80 g546620 ( .a(n_22172), .b(n_21411), .o(n_23415) );
in01f80 g546621 ( .a(n_21915), .o(n_22855) );
ao12f80 g546622 ( .a(n_9143), .b(n_21553), .c(n_7882), .o(n_21915) );
in01f80 g546623 ( .a(n_24556), .o(n_25539) );
oa12f80 g546624 ( .a(n_22368), .b(n_21754), .c(n_24203), .o(n_24556) );
ao12f80 g546625 ( .a(n_15857), .b(n_21552), .c(n_16495), .o(n_22563) );
ao12f80 g546626 ( .a(n_13218), .b(n_21551), .c(n_14448), .o(n_22564) );
oa12f80 g546627 ( .a(n_15560), .b(n_20874), .c(n_16268), .o(n_21978) );
oa12f80 g546628 ( .a(n_14780), .b(n_21550), .c(n_15416), .o(n_22562) );
oa12f80 g546629 ( .a(n_14768), .b(n_21187), .c(n_15410), .o(n_22269) );
in01f80 g546630 ( .a(n_23931), .o(n_24949) );
oa12f80 g546631 ( .a(n_22367), .b(n_21711), .c(n_23623), .o(n_23931) );
oa12f80 g546632 ( .a(n_14750), .b(n_21186), .c(n_15409), .o(n_22268) );
oa12f80 g546633 ( .a(n_14745), .b(n_21185), .c(n_15399), .o(n_22267) );
ao12f80 g546634 ( .a(n_14384), .b(n_21184), .c(n_15144), .o(n_22266) );
oa12f80 g546635 ( .a(n_14717), .b(n_21183), .c(n_15387), .o(n_22265) );
oa12f80 g546636 ( .a(n_14691), .b(n_21182), .c(n_15369), .o(n_22264) );
in01f80 g546637 ( .a(n_23344), .o(n_24312) );
oa12f80 g546638 ( .a(n_22098), .b(n_23061), .c(n_21371), .o(n_23344) );
ao12f80 g546639 ( .a(n_13156), .b(n_21549), .c(n_14315), .o(n_22561) );
in01f80 g546640 ( .a(n_24205), .o(n_25260) );
oa12f80 g546641 ( .a(n_22097), .b(n_23925), .c(n_21369), .o(n_24205) );
oa12f80 g546642 ( .a(n_16104), .b(n_22170), .c(n_16682), .o(n_23147) );
in01f80 g546643 ( .a(n_23930), .o(n_24932) );
oa12f80 g546644 ( .a(n_22095), .b(n_21359), .c(n_23621), .o(n_23930) );
ao12f80 g546645 ( .a(n_12292), .b(n_23058), .c(n_12951), .o(n_24026) );
in01f80 g546646 ( .a(n_23929), .o(n_24928) );
oa12f80 g546647 ( .a(n_22094), .b(n_23618), .c(n_21357), .o(n_23929) );
oa12f80 g546648 ( .a(n_15505), .b(n_22169), .c(n_16252), .o(n_23146) );
ao12f80 g546649 ( .a(n_11485), .b(n_21181), .c(n_12482), .o(n_22263) );
ao12f80 g546650 ( .a(n_12252), .b(n_21180), .c(n_12472), .o(n_22262) );
ao12f80 g546651 ( .a(n_14218), .b(n_21179), .c(n_15116), .o(n_22261) );
ao12f80 g546652 ( .a(n_14723), .b(n_21548), .c(n_15375), .o(n_22560) );
oa12f80 g546653 ( .a(n_11504), .b(n_20873), .c(n_12488), .o(n_21977) );
ao12f80 g546654 ( .a(n_14353), .b(n_21178), .c(n_15133), .o(n_22260) );
ao12f80 g546655 ( .a(n_15859), .b(n_21914), .c(n_16492), .o(n_22867) );
ao12f80 g546656 ( .a(n_14655), .b(n_21547), .c(n_15350), .o(n_22559) );
oa12f80 g546657 ( .a(n_13649), .b(n_21177), .c(n_14399), .o(n_22259) );
ao12f80 g546658 ( .a(n_13187), .b(n_22168), .c(n_14365), .o(n_23145) );
oa12f80 g546659 ( .a(n_14446), .b(n_21176), .c(n_15170), .o(n_22258) );
oa12f80 g546660 ( .a(n_14420), .b(n_21546), .c(n_15157), .o(n_22558) );
oa12f80 g546661 ( .a(n_10654), .b(n_20872), .c(n_11788), .o(n_21976) );
ao12f80 g546662 ( .a(n_13637), .b(n_21913), .c(n_14670), .o(n_22866) );
in01f80 g546663 ( .a(n_23690), .o(n_23343) );
ao12f80 g546664 ( .a(n_10911), .b(n_23059), .c(n_12083), .o(n_23690) );
ao12f80 g546665 ( .a(n_14259), .b(n_21175), .c(n_15101), .o(n_22257) );
ao12f80 g546666 ( .a(n_13903), .b(n_21174), .c(n_14912), .o(n_22256) );
ao12f80 g546667 ( .a(n_11514), .b(n_21545), .c(n_12493), .o(n_22557) );
ao12f80 g546668 ( .a(n_15800), .b(n_21173), .c(n_16475), .o(n_22255) );
ao12f80 g546669 ( .a(n_13883), .b(n_21172), .c(n_14907), .o(n_22254) );
oa12f80 g546670 ( .a(n_13961), .b(n_21171), .c(n_14934), .o(n_22253) );
oa12f80 g546671 ( .a(n_7718), .b(n_21170), .c(n_9094), .o(n_22251) );
ao12f80 g546672 ( .a(n_10665), .b(n_21169), .c(n_11799), .o(n_22252) );
ao12f80 g546673 ( .a(n_21488), .b(n_21487), .c(n_21486), .o(n_22167) );
in01f80 g546674 ( .a(n_21912), .o(n_22853) );
oa12f80 g546675 ( .a(n_20871), .b(n_21181), .c(n_20870), .o(n_21912) );
ao12f80 g546676 ( .a(n_23045), .b(n_23044), .c(n_23043), .o(n_23638) );
oa12f80 g546677 ( .a(n_21136), .b(n_21135), .c(n_21485), .o(n_22551) );
ao12f80 g546678 ( .a(n_23042), .b(n_23041), .c(n_23040), .o(n_23637) );
oa12f80 g546679 ( .a(n_21476), .b(n_21475), .c(n_21831), .o(n_22843) );
ao12f80 g546680 ( .a(n_23285), .b(n_23284), .c(n_23283), .o(n_23928) );
ao12f80 g546681 ( .a(n_22399), .b(n_22398), .c(n_22397), .o(n_23060) );
ao12f80 g546682 ( .a(n_23039), .b(n_23038), .c(n_23037), .o(n_23636) );
ao12f80 g546683 ( .a(n_22728), .b(n_22727), .c(n_22726), .o(n_23342) );
ao22s80 g546684 ( .a(n_22641), .b(n_24203), .c(n_22640), .d(n_23247), .o(n_24204) );
oa12f80 g546685 ( .a(n_21134), .b(n_21133), .c(n_21483), .o(n_22550) );
ao12f80 g546686 ( .a(n_21894), .b(n_21893), .c(n_21892), .o(n_22435) );
ao12f80 g546687 ( .a(n_23036), .b(n_23035), .c(n_23034), .o(n_23635) );
oa12f80 g546688 ( .a(n_21460), .b(n_21459), .c(n_21458), .o(n_22839) );
in01f80 g546689 ( .a(n_22485), .o(n_22838) );
ao12f80 g546690 ( .a(n_21168), .b(n_21552), .c(n_21167), .o(n_22485) );
ao12f80 g546691 ( .a(n_21825), .b(n_21824), .c(n_21823), .o(n_22434) );
ao12f80 g546692 ( .a(n_23033), .b(n_23032), .c(n_23031), .o(n_23634) );
in01f80 g546693 ( .a(n_22505), .o(n_22771) );
ao12f80 g546694 ( .a(n_21166), .b(n_21551), .c(n_21165), .o(n_22505) );
ao12f80 g546695 ( .a(n_22719), .b(n_22718), .c(n_22717), .o(n_23341) );
oa12f80 g546696 ( .a(n_21132), .b(n_21131), .c(n_21484), .o(n_22549) );
ao12f80 g546697 ( .a(n_22667), .b(n_22666), .c(n_22665), .o(n_23340) );
ao12f80 g546698 ( .a(n_22987), .b(n_22986), .c(n_22985), .o(n_23633) );
ao12f80 g546699 ( .a(n_22725), .b(n_22724), .c(n_22723), .o(n_23339) );
ao12f80 g546700 ( .a(n_23030), .b(n_23029), .c(n_23028), .o(n_23632) );
oa12f80 g546701 ( .a(n_21481), .b(n_21480), .c(n_21479), .o(n_22831) );
ao12f80 g546702 ( .a(n_22710), .b(n_22709), .c(n_22708), .o(n_23338) );
oa12f80 g546703 ( .a(n_21822), .b(n_22433), .c(n_21821), .o(n_23694) );
ao12f80 g546704 ( .a(n_22722), .b(n_22721), .c(n_22720), .o(n_23337) );
oa12f80 g546705 ( .a(n_21464), .b(n_21463), .c(n_21462), .o(n_22842) );
oa12f80 g546706 ( .a(n_21494), .b(n_21533), .c(n_21838), .o(n_22830) );
in01f80 g546707 ( .a(n_22503), .o(n_22547) );
ao12f80 g546708 ( .a(n_20849), .b(n_21176), .c(n_20848), .o(n_22503) );
ao12f80 g546709 ( .a(n_22716), .b(n_22715), .c(n_22714), .o(n_23576) );
in01f80 g546710 ( .a(n_22197), .o(n_22242) );
ao12f80 g546711 ( .a(n_20471), .b(n_20874), .c(n_20470), .o(n_22197) );
in01f80 g546712 ( .a(n_22519), .o(n_22825) );
ao12f80 g546713 ( .a(n_21164), .b(n_21550), .c(n_21163), .o(n_22519) );
ao12f80 g546714 ( .a(n_22713), .b(n_22712), .c(n_22711), .o(n_23281) );
ao12f80 g546715 ( .a(n_23027), .b(n_23026), .c(n_23025), .o(n_23617) );
oa12f80 g546716 ( .a(n_21145), .b(n_21161), .c(n_21498), .o(n_22543) );
oa12f80 g546717 ( .a(n_21836), .b(n_22591), .c(x_in_14_7), .o(n_24007) );
ao12f80 g546718 ( .a(n_23024), .b(n_23023), .c(n_23022), .o(n_23631) );
oa12f80 g546719 ( .a(n_21143), .b(n_21160), .c(n_21497), .o(n_22542) );
ao12f80 g546720 ( .a(n_22704), .b(n_22703), .c(n_22702), .o(n_23567) );
oa12f80 g546721 ( .a(n_21142), .b(n_21159), .c(n_21495), .o(n_22532) );
in01f80 g546722 ( .a(n_22232), .o(n_22541) );
ao12f80 g546723 ( .a(n_20869), .b(n_21187), .c(n_20868), .o(n_22232) );
ao12f80 g546724 ( .a(n_22701), .b(n_22700), .c(n_22699), .o(n_23248) );
oa12f80 g546725 ( .a(n_21144), .b(n_21162), .c(n_21499), .o(n_22544) );
oa12f80 g546726 ( .a(n_21141), .b(n_21158), .c(n_21496), .o(n_22540) );
ao12f80 g546727 ( .a(n_22993), .b(n_22992), .c(n_22991), .o(n_23639) );
ao12f80 g546728 ( .a(n_23015), .b(n_23014), .c(n_23013), .o(n_23630) );
ao12f80 g546729 ( .a(n_22707), .b(n_22706), .c(n_22705), .o(n_23453) );
ao12f80 g546730 ( .a(n_23288), .b(n_23287), .c(n_23286), .o(n_23927) );
in01f80 g546731 ( .a(n_22228), .o(n_22539) );
ao12f80 g546732 ( .a(n_20867), .b(n_21186), .c(n_20866), .o(n_22228) );
in01f80 g546733 ( .a(n_22767), .o(n_22811) );
ao12f80 g546734 ( .a(n_21147), .b(n_21546), .c(n_21146), .o(n_22767) );
ao12f80 g546735 ( .a(n_23012), .b(n_23011), .c(n_23266), .o(n_23580) );
in01f80 g546736 ( .a(n_22196), .o(n_22474) );
ao12f80 g546737 ( .a(n_20851), .b(n_21177), .c(n_20850), .o(n_22196) );
in01f80 g546738 ( .a(n_22230), .o(n_22538) );
ao12f80 g546739 ( .a(n_20865), .b(n_21185), .c(n_20864), .o(n_22230) );
ao12f80 g546740 ( .a(n_23010), .b(n_23009), .c(n_23008), .o(n_23640) );
in01f80 g546741 ( .a(n_22202), .o(n_22537) );
ao12f80 g546742 ( .a(n_20863), .b(n_21184), .c(n_20862), .o(n_22202) );
ao12f80 g546743 ( .a(n_22695), .b(n_22694), .c(n_22693), .o(n_23336) );
in01f80 g546744 ( .a(FE_OFN753_n_22913), .o(n_23692) );
oa12f80 g546745 ( .a(n_21840), .b(n_22168), .c(n_21839), .o(n_22913) );
ao12f80 g546746 ( .a(n_23607), .b(n_23606), .c(n_23605), .o(n_24200) );
ao12f80 g546747 ( .a(n_22692), .b(n_22691), .c(n_22690), .o(n_23335) );
in01f80 g546748 ( .a(n_22226), .o(n_22536) );
ao12f80 g546749 ( .a(n_20861), .b(n_21183), .c(n_20860), .o(n_22226) );
in01f80 g546750 ( .a(n_22215), .o(n_22535) );
ao12f80 g546751 ( .a(n_20853), .b(n_21178), .c(n_20852), .o(n_22215) );
ao12f80 g546752 ( .a(n_23007), .b(n_23006), .c(n_23005), .o(n_23629) );
in01f80 g546753 ( .a(n_22512), .o(n_22802) );
ao12f80 g546754 ( .a(n_21153), .b(n_21548), .c(n_21152), .o(n_22512) );
in01f80 g546755 ( .a(n_22224), .o(n_22534) );
ao12f80 g546756 ( .a(n_20859), .b(n_21182), .c(n_20858), .o(n_22224) );
ao12f80 g546757 ( .a(n_23004), .b(n_23003), .c(n_23002), .o(n_23628) );
in01f80 g546758 ( .a(n_22166), .o(n_23134) );
oa12f80 g546759 ( .a(n_21140), .b(n_21545), .c(n_21139), .o(n_22166) );
ao12f80 g546760 ( .a(n_22686), .b(n_22685), .c(n_22684), .o(n_23334) );
ao12f80 g546761 ( .a(n_21129), .b(n_21900), .c(n_21473), .o(n_22509) );
ao12f80 g546762 ( .a(n_20833), .b(n_20832), .c(n_20831), .o(n_21490) );
ao12f80 g546763 ( .a(n_23001), .b(n_23000), .c(n_22999), .o(n_23627) );
oa12f80 g546764 ( .a(n_21472), .b(n_21471), .c(n_21470), .o(n_22799) );
ao12f80 g546765 ( .a(n_22689), .b(n_22688), .c(n_22687), .o(n_23333) );
ao12f80 g546766 ( .a(n_22683), .b(n_22682), .c(n_22681), .o(n_23332) );
in01f80 g546767 ( .a(n_22213), .o(n_22533) );
ao12f80 g546768 ( .a(n_20839), .b(n_21171), .c(n_20838), .o(n_22213) );
in01f80 g546769 ( .a(n_22760), .o(n_23102) );
ao12f80 g546770 ( .a(n_21492), .b(n_21913), .c(n_21491), .o(n_22760) );
oa12f80 g546771 ( .a(n_22119), .b(n_22118), .c(n_22117), .o(n_23399) );
ao12f80 g546772 ( .a(n_22998), .b(n_22997), .c(n_23265), .o(n_23626) );
ao12f80 g546773 ( .a(n_21469), .b(n_21468), .c(n_21467), .o(n_22165) );
in01f80 g546774 ( .a(n_22200), .o(n_21911) );
oa12f80 g546775 ( .a(n_20835), .b(n_21170), .c(n_20834), .o(n_22200) );
ao22s80 g546776 ( .a(n_22364), .b(n_23061), .c(n_22363), .d(n_22086), .o(n_23331) );
oa12f80 g546777 ( .a(n_22403), .b(n_22427), .c(n_22654), .o(n_23679) );
in01f80 g546778 ( .a(FE_OFN921_n_22498), .o(n_22164) );
oa12f80 g546779 ( .a(n_21157), .b(n_21549), .c(n_21156), .o(n_22498) );
in01f80 g546780 ( .a(n_23668), .o(n_24015) );
ao22s80 g546781 ( .a(n_23059), .b(n_12522), .c(n_22089), .d(n_12523), .o(n_23668) );
ao12f80 g546782 ( .a(n_22996), .b(n_22995), .c(n_22994), .o(n_23625) );
ao22s80 g546783 ( .a(n_22361), .b(n_23925), .c(n_22360), .d(n_22955), .o(n_23926) );
in01f80 g546784 ( .a(n_22480), .o(n_22824) );
ao12f80 g546785 ( .a(n_21151), .b(n_21547), .c(n_21150), .o(n_22480) );
oa12f80 g546786 ( .a(n_21819), .b(n_21818), .c(n_21817), .o(n_23103) );
in01f80 g546787 ( .a(n_22483), .o(n_22531) );
ao12f80 g546788 ( .a(n_20843), .b(n_21173), .c(n_20842), .o(n_22483) );
in01f80 g546789 ( .a(n_24020), .o(n_23975) );
ao12f80 g546790 ( .a(n_22421), .b(n_22732), .c(n_22420), .o(n_24020) );
ao12f80 g546791 ( .a(n_22678), .b(n_22677), .c(n_22676), .o(n_23330) );
oa12f80 g546792 ( .a(n_22402), .b(n_22401), .c(n_22400), .o(n_23677) );
ao22s80 g546793 ( .a(n_22639), .b(n_23623), .c(n_22638), .d(n_22630), .o(n_23624) );
in01f80 g546794 ( .a(n_21936), .o(n_22206) );
ao12f80 g546795 ( .a(n_20469), .b(n_20873), .c(n_20468), .o(n_21936) );
ao12f80 g546796 ( .a(n_22675), .b(n_22674), .c(n_22673), .o(n_23329) );
in01f80 g546797 ( .a(n_23666), .o(n_23993) );
ao22s80 g546798 ( .a(n_22085), .b(n_13501), .c(n_23058), .d(n_13500), .o(n_23666) );
oa12f80 g546799 ( .a(n_22394), .b(n_22393), .c(n_22651), .o(n_23676) );
in01f80 g546800 ( .a(n_22495), .o(n_22530) );
ao12f80 g546801 ( .a(n_20847), .b(n_21175), .c(n_20846), .o(n_22495) );
ao12f80 g546802 ( .a(n_21127), .b(n_21126), .c(n_21125), .o(n_21910) );
in01f80 g546803 ( .a(n_22198), .o(n_22478) );
ao12f80 g546804 ( .a(n_20837), .b(n_21169), .c(n_20836), .o(n_22198) );
in01f80 g546805 ( .a(n_23087), .o(n_23393) );
ao12f80 g546806 ( .a(n_21857), .b(n_22170), .c(n_21856), .o(n_23087) );
ao22s80 g546807 ( .a(n_22359), .b(n_23621), .c(n_22358), .d(n_22629), .o(n_23622) );
ao12f80 g546808 ( .a(n_22990), .b(n_22989), .c(n_22988), .o(n_23620) );
ao22s80 g546809 ( .a(n_22357), .b(n_23618), .c(n_22356), .d(n_22628), .o(n_23619) );
ao12f80 g546810 ( .a(n_21138), .b(n_21541), .c(n_21137), .o(n_21909) );
in01f80 g546811 ( .a(n_21937), .o(n_22218) );
ao12f80 g546812 ( .a(n_20467), .b(n_20872), .c(n_20466), .o(n_21937) );
in01f80 g546813 ( .a(n_22492), .o(n_22529) );
ao12f80 g546814 ( .a(n_20845), .b(n_21174), .c(n_20844), .o(n_22492) );
in01f80 g546815 ( .a(n_23091), .o(n_23400) );
ao12f80 g546816 ( .a(n_21853), .b(n_22169), .c(n_21852), .o(n_23091) );
oa12f80 g546817 ( .a(n_22391), .b(n_22396), .c(n_22390), .o(n_24311) );
in01f80 g546818 ( .a(n_22163), .o(n_23130) );
oa12f80 g546819 ( .a(n_21149), .b(n_21553), .c(n_21148), .o(n_22163) );
ao12f80 g546820 ( .a(n_22982), .b(n_22981), .c(n_22980), .o(n_23616) );
ao12f80 g546821 ( .a(n_21512), .b(n_21511), .c(n_21510), .o(n_22162) );
in01f80 g546822 ( .a(n_21908), .o(n_22850) );
oa12f80 g546823 ( .a(n_20857), .b(n_21180), .c(n_20856), .o(n_21908) );
ao12f80 g546824 ( .a(n_23280), .b(n_23279), .c(n_23278), .o(n_23924) );
oa12f80 g546825 ( .a(n_22389), .b(n_22388), .c(n_22387), .o(n_23671) );
in01f80 g546826 ( .a(n_22489), .o(n_22526) );
ao12f80 g546827 ( .a(n_20841), .b(n_21172), .c(n_20840), .o(n_22489) );
ao12f80 g546828 ( .a(n_21508), .b(n_21507), .c(n_21506), .o(n_22161) );
ao12f80 g546829 ( .a(n_23277), .b(n_23276), .c(n_23275), .o(n_23923) );
oa12f80 g546830 ( .a(n_21124), .b(n_21123), .c(n_21482), .o(n_22548) );
ao12f80 g546831 ( .a(n_20830), .b(n_21544), .c(n_21121), .o(n_22223) );
ao12f80 g546832 ( .a(n_21120), .b(n_21119), .c(n_21118), .o(n_21907) );
ao12f80 g546833 ( .a(n_22662), .b(n_22661), .c(n_22660), .o(n_23328) );
oa12f80 g546834 ( .a(n_21493), .b(n_21519), .c(n_21837), .o(n_22783) );
ao12f80 g546835 ( .a(n_22979), .b(n_22978), .c(n_22977), .o(n_23615) );
ao12f80 g546836 ( .a(n_22659), .b(n_22658), .c(n_22657), .o(n_23327) );
oa12f80 g546837 ( .a(n_22121), .b(n_22731), .c(x_in_12_7), .o(n_23957) );
in01f80 g546838 ( .a(n_22211), .o(n_22523) );
ao12f80 g546839 ( .a(n_20855), .b(n_21179), .c(n_20854), .o(n_22211) );
ao12f80 g546840 ( .a(n_21835), .b(n_21834), .c(n_21833), .o(n_22432) );
in01f80 g546841 ( .a(n_23085), .o(n_23096) );
ao12f80 g546842 ( .a(n_21501), .b(n_21914), .c(n_21500), .o(n_23085) );
oa12f80 g546843 ( .a(n_21816), .b(n_21815), .c(n_22116), .o(n_23095) );
oa22f80 g546844 ( .a(n_21410), .b(FE_OFN314_n_3069), .c(n_1255), .d(FE_OFN119_n_27449), .o(n_22431) );
oa22f80 g546845 ( .a(FE_OFN632_n_21154), .b(n_29691), .c(n_557), .d(FE_OFN69_n_27012), .o(n_21543) );
oa22f80 g546846 ( .a(n_22350), .b(FE_OFN314_n_3069), .c(n_874), .d(FE_OFN72_n_27012), .o(n_23326) );
oa22f80 g546847 ( .a(n_22349), .b(FE_OFN309_n_3069), .c(n_597), .d(FE_OFN69_n_27012), .o(n_23325) );
oa22f80 g546848 ( .a(n_22627), .b(FE_OFN311_n_3069), .c(n_1743), .d(FE_OFN134_n_27449), .o(n_23614) );
oa22f80 g546849 ( .a(n_22084), .b(FE_OFN313_n_3069), .c(n_1553), .d(FE_OFN361_n_4860), .o(n_23057) );
oa22f80 g546850 ( .a(n_22348), .b(FE_OFN313_n_3069), .c(n_138), .d(FE_OFN1124_rst), .o(n_23324) );
oa22f80 g546851 ( .a(n_22077), .b(FE_OFN248_n_4162), .c(n_1853), .d(FE_OFN113_n_27449), .o(n_23056) );
oa22f80 g546852 ( .a(n_22954), .b(FE_OFN234_n_4162), .c(n_637), .d(FE_OFN127_n_27449), .o(n_23922) );
oa22f80 g546853 ( .a(n_21409), .b(FE_OFN311_n_3069), .c(n_774), .d(FE_OFN134_n_27449), .o(n_22430) );
oa22f80 g546854 ( .a(n_22347), .b(FE_OFN313_n_3069), .c(n_569), .d(FE_OFN131_n_27449), .o(n_23323) );
oa22f80 g546855 ( .a(n_21091), .b(FE_OFN310_n_3069), .c(n_1307), .d(FE_OFN1114_rst), .o(n_22160) );
oa22f80 g546856 ( .a(n_22346), .b(FE_OFN308_n_3069), .c(n_333), .d(FE_OFN114_n_27449), .o(n_23322) );
oa22f80 g546857 ( .a(FE_OFN508_n_22083), .b(FE_OFN214_n_29687), .c(n_1786), .d(n_28362), .o(n_23055) );
oa22f80 g546858 ( .a(n_22082), .b(FE_OFN308_n_3069), .c(n_916), .d(FE_OFN326_n_4860), .o(n_23054) );
oa22f80 g546859 ( .a(n_21090), .b(FE_OFN219_n_23315), .c(n_1401), .d(rst), .o(n_22159) );
oa22f80 g546860 ( .a(n_22345), .b(FE_OFN303_n_3069), .c(n_862), .d(FE_OFN1108_rst), .o(n_23321) );
oa22f80 g546861 ( .a(n_22344), .b(n_4280), .c(n_1501), .d(FE_OFN105_n_27449), .o(n_23320) );
oa22f80 g546862 ( .a(n_22326), .b(FE_OFN314_n_3069), .c(n_240), .d(FE_OFN93_n_27449), .o(n_23319) );
oa22f80 g546863 ( .a(FE_OFN1019_n_22081), .b(n_21076), .c(n_1171), .d(n_27449), .o(n_23053) );
oa22f80 g546864 ( .a(n_22080), .b(n_21076), .c(n_443), .d(FE_OFN96_n_27449), .o(n_23052) );
oa22f80 g546865 ( .a(n_22343), .b(FE_OFN253_n_4280), .c(n_1733), .d(FE_OFN136_n_27449), .o(n_23318) );
oa22f80 g546866 ( .a(n_22342), .b(n_23315), .c(n_1409), .d(FE_OFN95_n_27449), .o(n_23317) );
oa22f80 g546867 ( .a(n_22341), .b(n_23315), .c(n_304), .d(FE_OFN136_n_27449), .o(n_23316) );
oa22f80 g546868 ( .a(n_22335), .b(FE_OFN306_n_3069), .c(n_748), .d(FE_OFN125_n_27449), .o(n_23314) );
oa22f80 g546869 ( .a(FE_OFN847_n_22340), .b(n_29691), .c(n_326), .d(n_27449), .o(n_23313) );
oa22f80 g546870 ( .a(n_22338), .b(FE_OFN310_n_3069), .c(n_867), .d(FE_OFN1114_rst), .o(n_23312) );
oa22f80 g546871 ( .a(n_22327), .b(FE_OFN293_n_3069), .c(n_1243), .d(FE_OFN89_n_27449), .o(n_23311) );
oa22f80 g546872 ( .a(n_22339), .b(FE_OFN292_n_3069), .c(n_677), .d(FE_OFN101_n_27449), .o(n_23310) );
oa22f80 g546873 ( .a(n_20805), .b(n_26184), .c(n_336), .d(FE_OFN353_n_4860), .o(n_21906) );
oa22f80 g546874 ( .a(n_22319), .b(FE_OFN310_n_3069), .c(n_1282), .d(FE_OFN353_n_4860), .o(n_23309) );
oa22f80 g546875 ( .a(n_22337), .b(FE_OFN265_n_4280), .c(n_522), .d(FE_OFN1182_rst), .o(n_23308) );
oa22f80 g546876 ( .a(n_21541), .b(FE_OFN266_n_4280), .c(n_380), .d(FE_OFN287_n_29266), .o(n_21542) );
oa22f80 g546877 ( .a(n_21155), .b(n_29698), .c(n_1430), .d(FE_OFN286_n_29266), .o(n_21540) );
oa22f80 g546878 ( .a(n_22626), .b(FE_OFN293_n_3069), .c(n_495), .d(n_29104), .o(n_23612) );
oa22f80 g546879 ( .a(n_22336), .b(FE_OFN260_n_4280), .c(n_357), .d(FE_OFN125_n_27449), .o(n_23307) );
oa22f80 g546880 ( .a(n_20811), .b(FE_OFN299_n_3069), .c(n_904), .d(FE_OFN135_n_27449), .o(n_21905) );
oa22f80 g546881 ( .a(n_22334), .b(FE_OFN312_n_3069), .c(n_1122), .d(FE_OFN357_n_4860), .o(n_23306) );
oa22f80 g546882 ( .a(n_22079), .b(FE_OFN239_n_4162), .c(n_515), .d(FE_OFN360_n_4860), .o(n_23051) );
oa22f80 g546883 ( .a(n_21544), .b(x_in_52_7), .c(n_21122), .d(n_22222), .o(n_23985) );
oa22f80 g546884 ( .a(n_22122), .b(FE_OFN244_n_4162), .c(n_1581), .d(FE_OFN139_n_27449), .o(n_22429) );
oa22f80 g546885 ( .a(FE_OFN734_n_22952), .b(n_21076), .c(n_534), .d(FE_OFN96_n_27449), .o(n_23921) );
oa22f80 g546886 ( .a(n_22078), .b(FE_OFN253_n_4280), .c(n_292), .d(FE_OFN136_n_27449), .o(n_23050) );
oa22f80 g546887 ( .a(FE_OFN698_n_22333), .b(n_21076), .c(n_1235), .d(FE_OFN96_n_27449), .o(n_23305) );
oa22f80 g546888 ( .a(n_22332), .b(n_23291), .c(n_1866), .d(n_27449), .o(n_23302) );
oa22f80 g546889 ( .a(FE_OFN604_n_21535), .b(n_23291), .c(n_1862), .d(FE_OFN1117_rst), .o(n_21904) );
oa22f80 g546890 ( .a(n_22076), .b(FE_OFN254_n_4280), .c(n_4), .d(FE_OFN361_n_4860), .o(n_23049) );
oa22f80 g546891 ( .a(FE_OFN720_n_20807), .b(n_23291), .c(n_823), .d(FE_OFN63_n_27012), .o(n_21903) );
oa22f80 g546892 ( .a(n_22625), .b(FE_OFN254_n_4280), .c(n_89), .d(FE_OFN142_n_27449), .o(n_23611) );
oa22f80 g546893 ( .a(n_22331), .b(FE_OFN253_n_4280), .c(n_323), .d(FE_OFN136_n_27449), .o(n_23301) );
oa22f80 g546894 ( .a(n_22330), .b(FE_OFN265_n_4280), .c(n_1559), .d(FE_OFN1143_n_27012), .o(n_23300) );
oa22f80 g546895 ( .a(FE_OFN893_n_20806), .b(n_21076), .c(n_725), .d(FE_OFN68_n_27012), .o(n_21902) );
oa22f80 g546896 ( .a(FE_OFN877_n_22329), .b(n_21076), .c(n_354), .d(FE_OFN336_n_4860), .o(n_23299) );
oa22f80 g546897 ( .a(n_21478), .b(FE_OFN269_n_4280), .c(n_1197), .d(FE_OFN116_n_27449), .o(n_21901) );
oa22f80 g546898 ( .a(n_22328), .b(FE_OFN266_n_4280), .c(n_1873), .d(FE_OFN114_n_27449), .o(n_23298) );
oa22f80 g546899 ( .a(n_22624), .b(FE_OFN260_n_4280), .c(n_1890), .d(FE_OFN76_n_27012), .o(n_23610) );
oa22f80 g546900 ( .a(n_22075), .b(FE_OFN264_n_4280), .c(n_1479), .d(FE_OFN65_n_27012), .o(n_23048) );
oa22f80 g546901 ( .a(n_20444), .b(FE_OFN258_n_4280), .c(n_722), .d(FE_OFN358_n_4860), .o(n_21539) );
oa22f80 g546902 ( .a(n_22074), .b(FE_OFN313_n_3069), .c(n_177), .d(FE_OFN142_n_27449), .o(n_23047) );
oa22f80 g546903 ( .a(n_21900), .b(x_in_32_7), .c(n_21474), .d(n_22508), .o(n_23969) );
oa22f80 g546904 ( .a(n_21087), .b(FE_OFN166_n_29269), .c(n_49), .d(FE_OFN12_n_29204), .o(n_22158) );
oa22f80 g546905 ( .a(FE_OFN995_n_22325), .b(FE_OFN166_n_29269), .c(n_297), .d(FE_OFN12_n_29204), .o(n_23297) );
oa22f80 g546906 ( .a(n_22323), .b(FE_OFN410_n_28303), .c(n_1620), .d(FE_OFN74_n_27012), .o(n_23296) );
oa22f80 g546907 ( .a(n_21128), .b(FE_OFN240_n_4162), .c(n_470), .d(FE_OFN78_n_27012), .o(n_21538) );
oa22f80 g546908 ( .a(n_22322), .b(FE_OFN413_n_28303), .c(n_1159), .d(FE_OFN77_n_27012), .o(n_23295) );
oa22f80 g546909 ( .a(n_20804), .b(FE_OFN400_n_28303), .c(n_977), .d(FE_OFN92_n_27449), .o(n_21899) );
oa22f80 g546910 ( .a(n_21489), .b(FE_OFN416_n_28303), .c(n_1432), .d(FE_OFN108_n_27449), .o(n_21898) );
oa22f80 g546911 ( .a(n_22320), .b(FE_OFN269_n_4280), .c(n_1070), .d(FE_OFN90_n_27449), .o(n_23294) );
oa22f80 g546912 ( .a(n_21086), .b(FE_OFN406_n_28303), .c(n_114), .d(FE_OFN99_n_27449), .o(n_22157) );
oa22f80 g546913 ( .a(n_22951), .b(FE_OFN293_n_3069), .c(n_90), .d(FE_OFN357_n_4860), .o(n_23920) );
oa22f80 g546914 ( .a(n_21085), .b(FE_OFN311_n_3069), .c(n_1818), .d(FE_OFN1174_n_4860), .o(n_22156) );
oa22f80 g546915 ( .a(n_22622), .b(FE_OFN416_n_28303), .c(n_690), .d(FE_OFN134_n_27449), .o(n_23609) );
oa22f80 g546916 ( .a(n_22351), .b(FE_OFN405_n_28303), .c(n_614), .d(FE_OFN98_n_27449), .o(n_23293) );
oa22f80 g546917 ( .a(FE_OFN939_n_21084), .b(n_23291), .c(n_69), .d(FE_OFN105_n_27449), .o(n_22155) );
oa22f80 g546918 ( .a(FE_OFN935_n_22317), .b(n_23291), .c(n_1215), .d(FE_OFN105_n_27449), .o(n_23292) );
oa22f80 g546919 ( .a(n_22316), .b(n_28303), .c(n_1007), .d(n_25680), .o(n_23290) );
oa22f80 g546920 ( .a(FE_OFN520_n_22315), .b(FE_OFN165_n_29269), .c(n_1783), .d(n_25680), .o(n_23289) );
oa22f80 g546921 ( .a(n_21408), .b(FE_OFN166_n_29269), .c(n_248), .d(FE_OFN1123_rst), .o(n_22428) );
oa22f80 g546922 ( .a(n_22433), .b(x_in_6_7), .c(n_21477), .d(n_467), .o(n_24268) );
in01f80 g546999 ( .a(n_22729), .o(n_22730) );
no02f80 g547000 ( .a(n_22427), .b(x_in_8_10), .o(n_22729) );
na02f80 g547001 ( .a(n_22427), .b(x_in_8_10), .o(n_23362) );
oa12f80 g547002 ( .a(n_21416), .b(n_8786), .c(n_9934), .o(n_23083) );
na02f80 g547003 ( .a(n_21181), .b(n_20870), .o(n_20871) );
no02f80 g547004 ( .a(n_23044), .b(n_23043), .o(n_23045) );
na02f80 g547005 ( .a(n_21897), .b(x_in_2_7), .o(n_22750) );
in01f80 g547006 ( .a(n_22153), .o(n_22154) );
no02f80 g547007 ( .a(n_21897), .b(x_in_2_7), .o(n_22153) );
in01f80 g547008 ( .a(n_22151), .o(n_22152) );
no02f80 g547009 ( .a(n_21880), .b(x_in_40_7), .o(n_22151) );
no02f80 g547010 ( .a(n_23041), .b(n_23040), .o(n_23042) );
na02f80 g547011 ( .a(n_22150), .b(x_in_34_7), .o(n_23065) );
in01f80 g547012 ( .a(n_22425), .o(n_22426) );
no02f80 g547013 ( .a(n_22150), .b(x_in_34_7), .o(n_22425) );
na02f80 g547014 ( .a(n_21529), .b(x_in_62_7), .o(n_22458) );
no02f80 g547015 ( .a(n_23038), .b(n_23037), .o(n_23039) );
no02f80 g547016 ( .a(n_22727), .b(n_22726), .o(n_22728) );
na02f80 g547017 ( .a(n_21537), .b(x_in_18_7), .o(n_22465) );
in01f80 g547018 ( .a(n_21895), .o(n_21896) );
no02f80 g547019 ( .a(n_21537), .b(x_in_18_7), .o(n_21895) );
no02f80 g547020 ( .a(n_21893), .b(n_21892), .o(n_21894) );
no02f80 g547021 ( .a(n_23035), .b(n_23034), .o(n_23036) );
na02f80 g547022 ( .a(n_21536), .b(x_in_50_7), .o(n_22456) );
in01f80 g547023 ( .a(n_21890), .o(n_21891) );
no02f80 g547024 ( .a(n_21536), .b(x_in_50_7), .o(n_21890) );
no02f80 g547025 ( .a(n_21552), .b(n_21167), .o(n_21168) );
no02f80 g547026 ( .a(n_23032), .b(n_23031), .o(n_23033) );
na02f80 g547027 ( .a(n_21889), .b(x_in_10_7), .o(n_22748) );
in01f80 g547028 ( .a(n_22148), .o(n_22149) );
no02f80 g547029 ( .a(n_21889), .b(x_in_10_7), .o(n_22148) );
na02f80 g547030 ( .a(FE_OFN604_n_21535), .b(n_21892), .o(n_22840) );
na02f80 g547031 ( .a(n_22696), .b(x_in_56_9), .o(n_23651) );
na02f80 g547032 ( .a(n_21888), .b(x_in_42_7), .o(n_22747) );
in01f80 g547033 ( .a(n_22146), .o(n_22147) );
no02f80 g547034 ( .a(n_21888), .b(x_in_42_7), .o(n_22146) );
no02f80 g547035 ( .a(n_21551), .b(n_21165), .o(n_21166) );
na02f80 g547036 ( .a(n_21887), .b(x_in_26_7), .o(n_22737) );
in01f80 g547037 ( .a(n_22144), .o(n_22145) );
no02f80 g547038 ( .a(n_21887), .b(x_in_26_7), .o(n_22144) );
in01f80 g547039 ( .a(n_22142), .o(n_22143) );
na02f80 g547040 ( .a(n_21886), .b(n_21112), .o(n_22142) );
no02f80 g547041 ( .a(n_22724), .b(n_22723), .o(n_22725) );
no02f80 g547042 ( .a(n_23029), .b(n_23028), .o(n_23030) );
na02f80 g547043 ( .a(n_21528), .b(x_in_58_7), .o(n_22464) );
in01f80 g547044 ( .a(n_24570), .o(n_22141) );
no02f80 g547045 ( .a(n_21851), .b(x_in_6_6), .o(n_24570) );
no02f80 g547046 ( .a(n_22721), .b(n_22720), .o(n_22722) );
no02f80 g547047 ( .a(n_22718), .b(n_22717), .o(n_22719) );
na02f80 g547048 ( .a(n_21885), .b(x_in_22_7), .o(n_22745) );
in01f80 g547049 ( .a(n_22139), .o(n_22140) );
no02f80 g547050 ( .a(n_21885), .b(x_in_22_7), .o(n_22139) );
no02f80 g547051 ( .a(n_23287), .b(n_23286), .o(n_23288) );
no02f80 g547052 ( .a(n_20874), .b(n_20470), .o(n_20471) );
na02f80 g547053 ( .a(n_21505), .b(x_in_2_8), .o(n_22457) );
no02f80 g547054 ( .a(n_22715), .b(n_22714), .o(n_22716) );
na02f80 g547055 ( .a(n_21534), .b(x_in_54_7), .o(n_22453) );
in01f80 g547056 ( .a(n_21883), .o(n_21884) );
no02f80 g547057 ( .a(n_21534), .b(x_in_54_7), .o(n_21883) );
no02f80 g547058 ( .a(n_21550), .b(n_21163), .o(n_21164) );
na02f80 g547059 ( .a(n_21533), .b(x_in_22_8), .o(n_22460) );
in01f80 g547060 ( .a(n_21881), .o(n_21882) );
no02f80 g547061 ( .a(n_21533), .b(x_in_22_8), .o(n_21881) );
no02f80 g547062 ( .a(n_22712), .b(n_22711), .o(n_22713) );
na02f80 g547063 ( .a(n_21880), .b(x_in_40_7), .o(n_22736) );
no02f80 g547064 ( .a(n_23026), .b(n_23025), .o(n_23027) );
no02f80 g547065 ( .a(n_23023), .b(n_23022), .o(n_23024) );
na02f80 g547066 ( .a(n_21504), .b(x_in_46_7), .o(n_22461) );
no02f80 g547067 ( .a(n_22709), .b(n_22708), .o(n_22710) );
no02f80 g547068 ( .a(n_22706), .b(n_22705), .o(n_22707) );
no02f80 g547069 ( .a(n_22703), .b(n_22702), .o(n_22704) );
na02f80 g547070 ( .a(n_21532), .b(x_in_30_7), .o(n_22459) );
in01f80 g547071 ( .a(n_21878), .o(n_21879) );
no02f80 g547072 ( .a(n_21532), .b(x_in_30_7), .o(n_21878) );
no02f80 g547073 ( .a(n_22700), .b(n_22699), .o(n_22701) );
na02f80 g547074 ( .a(n_21162), .b(x_in_54_8), .o(n_22190) );
in01f80 g547075 ( .a(n_21530), .o(n_21531) );
no02f80 g547076 ( .a(n_21162), .b(x_in_54_8), .o(n_21530) );
in01f80 g547077 ( .a(n_21876), .o(n_21877) );
no02f80 g547078 ( .a(n_21529), .b(x_in_62_7), .o(n_21876) );
in01f80 g547079 ( .a(n_21874), .o(n_21875) );
no02f80 g547080 ( .a(n_21528), .b(x_in_58_7), .o(n_21874) );
no02f80 g547081 ( .a(n_21187), .b(n_20868), .o(n_20869) );
in01f80 g547082 ( .a(n_23020), .o(n_23021) );
na02f80 g547083 ( .a(n_22698), .b(n_22102), .o(n_23020) );
in01f80 g547084 ( .a(n_23018), .o(n_23019) );
na02f80 g547085 ( .a(n_22697), .b(n_22104), .o(n_23018) );
in01f80 g547086 ( .a(n_23016), .o(n_23017) );
no02f80 g547087 ( .a(n_22696), .b(x_in_56_9), .o(n_23016) );
no02f80 g547088 ( .a(n_23014), .b(n_23013), .o(n_23015) );
no02f80 g547089 ( .a(n_23284), .b(n_23283), .o(n_23285) );
no02f80 g547090 ( .a(n_21186), .b(n_20866), .o(n_20867) );
in01f80 g547091 ( .a(n_21526), .o(n_21527) );
na02f80 g547092 ( .a(n_21161), .b(x_in_14_8), .o(n_21526) );
no02f80 g547093 ( .a(n_21161), .b(x_in_14_8), .o(n_22189) );
no02f80 g547094 ( .a(n_23011), .b(n_23266), .o(n_23012) );
na02f80 g547095 ( .a(n_21873), .b(x_in_34_8), .o(n_22744) );
in01f80 g547096 ( .a(n_22137), .o(n_22138) );
no02f80 g547097 ( .a(n_21873), .b(x_in_34_8), .o(n_22137) );
no02f80 g547098 ( .a(n_21185), .b(n_20864), .o(n_20865) );
na02f80 g547099 ( .a(n_21160), .b(x_in_46_8), .o(n_22187) );
in01f80 g547100 ( .a(n_21524), .o(n_21525) );
no02f80 g547101 ( .a(n_21160), .b(x_in_46_8), .o(n_21524) );
no02f80 g547102 ( .a(n_23009), .b(n_23008), .o(n_23010) );
no02f80 g547103 ( .a(n_21184), .b(n_20862), .o(n_20863) );
na02f80 g547104 ( .a(n_21523), .b(x_in_16_8), .o(n_22452) );
in01f80 g547105 ( .a(n_21871), .o(n_21872) );
no02f80 g547106 ( .a(n_21523), .b(x_in_16_8), .o(n_21871) );
no02f80 g547107 ( .a(n_22694), .b(n_22693), .o(n_22695) );
no02f80 g547108 ( .a(n_23606), .b(n_23605), .o(n_23607) );
no02f80 g547109 ( .a(n_22691), .b(n_22690), .o(n_22692) );
no02f80 g547110 ( .a(n_21183), .b(n_20860), .o(n_20861) );
na02f80 g547111 ( .a(n_21159), .b(x_in_30_8), .o(n_22186) );
in01f80 g547112 ( .a(n_21521), .o(n_21522) );
no02f80 g547113 ( .a(n_21159), .b(x_in_30_8), .o(n_21521) );
na02f80 g547114 ( .a(n_21520), .b(x_in_18_8), .o(n_22451) );
in01f80 g547115 ( .a(n_21869), .o(n_21870) );
no02f80 g547116 ( .a(n_21520), .b(x_in_18_8), .o(n_21869) );
no02f80 g547117 ( .a(n_23006), .b(n_23005), .o(n_23007) );
in01f80 g547118 ( .a(n_21867), .o(n_21868) );
na02f80 g547119 ( .a(n_21519), .b(x_in_12_8), .o(n_21867) );
no02f80 g547120 ( .a(n_21519), .b(x_in_12_8), .o(n_22446) );
no02f80 g547121 ( .a(n_21182), .b(n_20858), .o(n_20859) );
na02f80 g547122 ( .a(n_21158), .b(x_in_62_8), .o(n_22185) );
in01f80 g547123 ( .a(n_21517), .o(n_21518) );
no02f80 g547124 ( .a(n_21158), .b(x_in_62_8), .o(n_21517) );
no02f80 g547125 ( .a(n_22688), .b(n_22687), .o(n_22689) );
no02f80 g547126 ( .a(n_23003), .b(n_23002), .o(n_23004) );
na02f80 g547127 ( .a(n_21866), .b(x_in_32_6), .o(n_22743) );
no02f80 g547128 ( .a(n_22685), .b(n_22684), .o(n_22686) );
in01f80 g547129 ( .a(n_22135), .o(n_22136) );
no02f80 g547130 ( .a(n_21866), .b(x_in_32_6), .o(n_22135) );
no02f80 g547131 ( .a(n_23000), .b(n_22999), .o(n_23001) );
na02f80 g547132 ( .a(n_21516), .b(x_in_16_7), .o(n_22447) );
in01f80 g547133 ( .a(n_21864), .o(n_21865) );
no02f80 g547134 ( .a(n_21516), .b(x_in_16_7), .o(n_21864) );
no02f80 g547135 ( .a(n_22682), .b(n_22681), .o(n_22683) );
na02f80 g547136 ( .a(n_21515), .b(x_in_50_8), .o(n_22445) );
in01f80 g547137 ( .a(n_21862), .o(n_21863) );
no02f80 g547138 ( .a(n_21515), .b(x_in_50_8), .o(n_21862) );
in01f80 g547139 ( .a(n_22423), .o(n_22424) );
no02f80 g547140 ( .a(n_22134), .b(x_in_48_6), .o(n_22423) );
na02f80 g547141 ( .a(n_22134), .b(x_in_48_6), .o(n_23071) );
no02f80 g547142 ( .a(n_22997), .b(n_23265), .o(n_22998) );
na02f80 g547143 ( .a(n_22422), .b(x_in_8_9), .o(n_23359) );
in01f80 g547144 ( .a(n_22679), .o(n_22680) );
no02f80 g547145 ( .a(n_22422), .b(x_in_8_9), .o(n_22679) );
na02f80 g547146 ( .a(n_21549), .b(n_21156), .o(n_21157) );
no02f80 g547147 ( .a(n_22995), .b(n_22994), .o(n_22996) );
in01f80 g547148 ( .a(n_22132), .o(n_22133) );
no02f80 g547149 ( .a(n_21861), .b(x_in_40_6), .o(n_22132) );
na02f80 g547150 ( .a(n_21861), .b(x_in_40_6), .o(n_22740) );
no02f80 g547151 ( .a(n_22677), .b(n_22676), .o(n_22678) );
no02f80 g547152 ( .a(n_22732), .b(n_22420), .o(n_22421) );
na02f80 g547153 ( .a(n_21860), .b(x_in_24_10), .o(n_22739) );
in01f80 g547154 ( .a(n_22130), .o(n_22131) );
no02f80 g547155 ( .a(n_21860), .b(x_in_24_10), .o(n_22130) );
no02f80 g547156 ( .a(n_22674), .b(n_22673), .o(n_22675) );
in01f80 g547157 ( .a(n_23603), .o(n_23604) );
na02f80 g547158 ( .a(n_23282), .b(n_22637), .o(n_23603) );
in01f80 g547159 ( .a(n_22418), .o(n_22419) );
na02f80 g547160 ( .a(n_22129), .b(n_21433), .o(n_22418) );
in01f80 g547161 ( .a(n_22416), .o(n_22417) );
na02f80 g547162 ( .a(n_22128), .b(n_21429), .o(n_22416) );
na02f80 g547163 ( .a(n_22415), .b(x_in_56_8), .o(n_23356) );
in01f80 g547164 ( .a(n_22671), .o(n_22672) );
no02f80 g547165 ( .a(n_22415), .b(x_in_56_8), .o(n_22671) );
na02f80 g547166 ( .a(n_21514), .b(x_in_10_8), .o(n_22444) );
in01f80 g547167 ( .a(n_21858), .o(n_21859) );
no02f80 g547168 ( .a(n_21514), .b(x_in_10_8), .o(n_21858) );
no02f80 g547169 ( .a(n_22170), .b(n_21856), .o(n_21857) );
na02f80 g547170 ( .a(n_22412), .b(x_in_20_7), .o(n_23363) );
na02f80 g547171 ( .a(n_22127), .b(x_in_48_7), .o(n_23064) );
in01f80 g547172 ( .a(n_22413), .o(n_22414) );
no02f80 g547173 ( .a(n_22127), .b(x_in_48_7), .o(n_22413) );
in01f80 g547174 ( .a(n_22669), .o(n_22670) );
no02f80 g547175 ( .a(n_22412), .b(x_in_20_7), .o(n_22669) );
no02f80 g547176 ( .a(n_22992), .b(n_22991), .o(n_22993) );
no02f80 g547177 ( .a(n_22989), .b(n_22988), .o(n_22990) );
no02f80 g547178 ( .a(n_22986), .b(n_22985), .o(n_22987) );
na02f80 g547179 ( .a(n_21513), .b(x_in_42_8), .o(n_22443) );
in01f80 g547180 ( .a(n_21854), .o(n_21855) );
no02f80 g547181 ( .a(n_21513), .b(x_in_42_8), .o(n_21854) );
no02f80 g547182 ( .a(n_22169), .b(n_21852), .o(n_21853) );
in01f80 g547183 ( .a(n_23643), .o(n_22984) );
na02f80 g547184 ( .a(n_22668), .b(x_in_36_6), .o(n_23643) );
in01f80 g547185 ( .a(n_25230), .o(n_22983) );
no02f80 g547186 ( .a(n_22668), .b(x_in_36_6), .o(n_25230) );
in01f80 g547187 ( .a(n_22749), .o(n_22126) );
na02f80 g547188 ( .a(n_21851), .b(x_in_6_6), .o(n_22749) );
no02f80 g547189 ( .a(n_22981), .b(n_22980), .o(n_22982) );
no02f80 g547190 ( .a(n_21511), .b(n_21510), .o(n_21512) );
na02f80 g547191 ( .a(n_21180), .b(n_20856), .o(n_20857) );
na02f80 g547192 ( .a(n_21155), .b(n_21510), .o(n_22527) );
no02f80 g547193 ( .a(n_22666), .b(n_22665), .o(n_22667) );
no02f80 g547194 ( .a(n_23279), .b(n_23278), .o(n_23280) );
in01f80 g547195 ( .a(n_22663), .o(n_22664) );
no02f80 g547196 ( .a(n_22411), .b(x_in_20_6), .o(n_22663) );
na02f80 g547197 ( .a(n_22411), .b(x_in_20_6), .o(n_23353) );
na02f80 g547198 ( .a(n_21509), .b(x_in_26_8), .o(n_22441) );
in01f80 g547199 ( .a(n_21849), .o(n_21850) );
no02f80 g547200 ( .a(n_21509), .b(x_in_26_8), .o(n_21849) );
no02f80 g547201 ( .a(n_21507), .b(n_21506), .o(n_21508) );
na02f80 g547202 ( .a(FE_OFN632_n_21154), .b(n_21506), .o(n_22524) );
no02f80 g547203 ( .a(n_23276), .b(n_23275), .o(n_23277) );
in01f80 g547204 ( .a(n_21847), .o(n_21848) );
no02f80 g547205 ( .a(n_21505), .b(x_in_2_8), .o(n_21847) );
in01f80 g547206 ( .a(n_21845), .o(n_21846) );
no02f80 g547207 ( .a(n_21504), .b(x_in_46_7), .o(n_21845) );
in01f80 g547208 ( .a(n_21843), .o(n_21844) );
no02f80 g547209 ( .a(n_21503), .b(x_in_52_6), .o(n_21843) );
na02f80 g547210 ( .a(n_21503), .b(x_in_52_6), .o(n_22442) );
no02f80 g547211 ( .a(n_22661), .b(n_22660), .o(n_22662) );
in01f80 g547212 ( .a(n_22409), .o(n_22410) );
na02f80 g547213 ( .a(n_22125), .b(n_21447), .o(n_22409) );
no02f80 g547214 ( .a(n_22978), .b(n_22977), .o(n_22979) );
no02f80 g547215 ( .a(n_22658), .b(n_22657), .o(n_22659) );
in01f80 g547216 ( .a(n_23601), .o(n_23602) );
na02f80 g547217 ( .a(n_23274), .b(n_22634), .o(n_23601) );
no02f80 g547218 ( .a(n_21179), .b(n_20854), .o(n_20855) );
na02f80 g547219 ( .a(n_21502), .b(x_in_58_8), .o(n_22466) );
in01f80 g547220 ( .a(n_21841), .o(n_21842) );
no02f80 g547221 ( .a(n_21502), .b(x_in_58_8), .o(n_21841) );
na02f80 g547222 ( .a(n_22124), .b(x_in_60_7), .o(n_23074) );
in01f80 g547223 ( .a(n_22407), .o(n_22408) );
no02f80 g547224 ( .a(n_22124), .b(x_in_60_7), .o(n_22407) );
in01f80 g547225 ( .a(n_22405), .o(n_22406) );
na02f80 g547226 ( .a(n_22123), .b(n_21424), .o(n_22405) );
in01f80 g547227 ( .a(n_22655), .o(n_22656) );
no02f80 g547228 ( .a(n_22404), .b(x_in_60_6), .o(n_22655) );
na02f80 g547229 ( .a(n_22404), .b(x_in_60_6), .o(n_23364) );
no02f80 g547230 ( .a(n_21548), .b(n_21152), .o(n_21153) );
no02f80 g547231 ( .a(n_20873), .b(n_20468), .o(n_20469) );
no02f80 g547232 ( .a(n_21178), .b(n_20852), .o(n_20853) );
no02f80 g547233 ( .a(n_21914), .b(n_21500), .o(n_21501) );
na02f80 g547234 ( .a(n_22427), .b(n_22654), .o(n_22403) );
no02f80 g547235 ( .a(n_21547), .b(n_21150), .o(n_21151) );
no02f80 g547236 ( .a(n_21177), .b(n_20850), .o(n_20851) );
na02f80 g547237 ( .a(n_22168), .b(n_21839), .o(n_21840) );
no02f80 g547238 ( .a(n_21176), .b(n_20848), .o(n_20849) );
na02f80 g547239 ( .a(n_21553), .b(n_21148), .o(n_21149) );
no02f80 g547240 ( .a(n_21546), .b(n_21146), .o(n_21147) );
no02f80 g547241 ( .a(n_20872), .b(n_20466), .o(n_20467) );
na02f80 g547242 ( .a(n_21161), .b(n_21498), .o(n_21145) );
na02f80 g547243 ( .a(n_21089), .b(n_21838), .o(n_22778) );
na02f80 g547244 ( .a(n_21162), .b(n_21499), .o(n_21144) );
na02f80 g547245 ( .a(n_20813), .b(n_21499), .o(n_22518) );
na02f80 g547246 ( .a(n_20812), .b(n_21498), .o(n_22514) );
na02f80 g547247 ( .a(n_21160), .b(n_21497), .o(n_21143) );
na02f80 g547248 ( .a(n_20810), .b(n_21497), .o(n_22515) );
na02f80 g547249 ( .a(n_21159), .b(n_21495), .o(n_21142) );
na02f80 g547250 ( .a(n_20808), .b(n_21496), .o(n_22516) );
na02f80 g547251 ( .a(n_21158), .b(n_21496), .o(n_21141) );
na02f80 g547252 ( .a(n_20809), .b(n_21495), .o(n_22517) );
na02f80 g547253 ( .a(n_22087), .b(n_22654), .o(n_23953) );
na02f80 g547254 ( .a(n_22401), .b(n_22400), .o(n_22402) );
na02f80 g547255 ( .a(n_22401), .b(n_21647), .o(n_23374) );
na02f80 g547256 ( .a(n_21533), .b(n_21838), .o(n_21494) );
na02f80 g547257 ( .a(n_21088), .b(n_21837), .o(n_22777) );
na02f80 g547258 ( .a(n_21519), .b(n_21837), .o(n_21493) );
in01f80 g547259 ( .a(n_23075), .o(n_23350) );
na02f80 g547260 ( .a(n_21778), .b(n_4846), .o(n_23075) );
no02f80 g547261 ( .a(n_21913), .b(n_21491), .o(n_21492) );
no02f80 g547262 ( .a(n_21175), .b(n_20846), .o(n_20847) );
no02f80 g547263 ( .a(n_21174), .b(n_20844), .o(n_20845) );
no02f80 g547264 ( .a(n_22398), .b(n_22397), .o(n_22399) );
na02f80 g547265 ( .a(n_22122), .b(n_22397), .o(n_23380) );
na02f80 g547266 ( .a(n_22591), .b(x_in_14_7), .o(n_21836) );
na02f80 g547267 ( .a(n_22396), .b(n_22395), .o(n_23349) );
in01f80 g547268 ( .a(n_22652), .o(n_22653) );
no02f80 g547269 ( .a(n_22396), .b(n_22395), .o(n_22652) );
na02f80 g547270 ( .a(n_22731), .b(x_in_12_7), .o(n_22121) );
na02f80 g547271 ( .a(n_21545), .b(n_21139), .o(n_21140) );
no02f80 g547272 ( .a(n_21173), .b(n_20842), .o(n_20843) );
no02f80 g547273 ( .a(n_21172), .b(n_20840), .o(n_20841) );
no02f80 g547274 ( .a(n_21171), .b(n_20838), .o(n_20839) );
no02f80 g547275 ( .a(n_21834), .b(n_21833), .o(n_21835) );
na02f80 g547276 ( .a(n_21489), .b(n_21833), .o(n_22773) );
no02f80 g547277 ( .a(n_21169), .b(n_20836), .o(n_20837) );
no02f80 g547278 ( .a(n_21541), .b(n_21137), .o(n_21138) );
no02f80 g547279 ( .a(n_20443), .b(n_21137), .o(n_22217) );
na02f80 g547280 ( .a(n_21170), .b(n_20834), .o(n_20835) );
no02f80 g547281 ( .a(n_21487), .b(n_21486), .o(n_21488) );
no02f80 g547282 ( .a(n_21487), .b(n_20707), .o(n_22770) );
in01f80 g547283 ( .a(n_21832), .o(n_22502) );
no02f80 g547284 ( .a(n_21505), .b(n_21485), .o(n_21832) );
na02f80 g547285 ( .a(n_21135), .b(n_21485), .o(n_21136) );
in01f80 g547286 ( .a(n_22120), .o(n_22766) );
no02f80 g547287 ( .a(n_21873), .b(n_21831), .o(n_22120) );
na02f80 g547288 ( .a(n_21133), .b(n_21483), .o(n_21134) );
na02f80 g547289 ( .a(n_21463), .b(n_20715), .o(n_22501) );
na02f80 g547290 ( .a(n_21459), .b(n_20714), .o(n_22500) );
in01f80 g547291 ( .a(n_21830), .o(n_22491) );
no02f80 g547292 ( .a(n_21513), .b(n_21484), .o(n_21830) );
na02f80 g547293 ( .a(n_21131), .b(n_21484), .o(n_21132) );
in01f80 g547294 ( .a(n_21829), .o(n_22494) );
no02f80 g547295 ( .a(n_21514), .b(n_21483), .o(n_21829) );
in01f80 g547296 ( .a(n_21828), .o(n_22488) );
no02f80 g547297 ( .a(n_21509), .b(n_21482), .o(n_21828) );
na02f80 g547298 ( .a(n_21480), .b(n_20713), .o(n_22487) );
na02f80 g547299 ( .a(n_21480), .b(n_21479), .o(n_21481) );
in01f80 g547300 ( .a(n_21827), .o(n_22497) );
na02f80 g547301 ( .a(n_21478), .b(n_21823), .o(n_21827) );
in01f80 g547302 ( .a(n_22484), .o(n_21826) );
na02f80 g547303 ( .a(n_21477), .b(n_21821), .o(n_22484) );
na02f80 g547304 ( .a(n_21475), .b(n_21831), .o(n_21476) );
no02f80 g547305 ( .a(n_21824), .b(n_21823), .o(n_21825) );
oa12f80 g547306 ( .a(n_12505), .b(n_21130), .c(n_11559), .o(n_22194) );
na02f80 g547307 ( .a(n_22433), .b(n_21821), .o(n_21822) );
in01f80 g547308 ( .a(n_22208), .o(n_21820) );
na02f80 g547309 ( .a(n_21474), .b(n_21473), .o(n_22208) );
no02f80 g547310 ( .a(n_21900), .b(n_21473), .o(n_21129) );
no02f80 g547311 ( .a(n_20832), .b(n_20831), .o(n_20833) );
no02f80 g547312 ( .a(n_20832), .b(n_20044), .o(n_22205) );
na02f80 g547313 ( .a(n_21471), .b(n_20712), .o(n_22482) );
na02f80 g547314 ( .a(n_21471), .b(n_21470), .o(n_21472) );
na02f80 g547315 ( .a(n_22118), .b(n_21340), .o(n_23093) );
na02f80 g547316 ( .a(n_22118), .b(n_22117), .o(n_22119) );
no02f80 g547317 ( .a(n_21468), .b(n_21467), .o(n_21469) );
in01f80 g547318 ( .a(n_21466), .o(n_22199) );
na02f80 g547319 ( .a(n_21128), .b(n_21467), .o(n_21466) );
oa12f80 g547320 ( .a(n_21415), .b(n_21465), .c(n_8785), .o(n_22182) );
na02f80 g547321 ( .a(n_21818), .b(n_21024), .o(n_22759) );
na02f80 g547322 ( .a(n_21818), .b(n_21817), .o(n_21819) );
in01f80 g547323 ( .a(n_22976), .o(n_23665) );
no02f80 g547324 ( .a(n_22696), .b(n_22651), .o(n_22976) );
na02f80 g547325 ( .a(n_22393), .b(n_22651), .o(n_22394) );
no02f80 g547326 ( .a(n_21126), .b(n_21125), .o(n_21127) );
no02f80 g547327 ( .a(n_21126), .b(n_20364), .o(n_22477) );
na02f80 g547328 ( .a(n_21463), .b(n_21462), .o(n_21464) );
in01f80 g547329 ( .a(n_22392), .o(n_23089) );
no02f80 g547330 ( .a(n_21775), .b(n_22390), .o(n_22392) );
na02f80 g547331 ( .a(n_22396), .b(n_22390), .o(n_22391) );
na02f80 g547332 ( .a(n_21123), .b(n_21482), .o(n_21124) );
na02f80 g547333 ( .a(n_22388), .b(n_21655), .o(n_23375) );
na02f80 g547334 ( .a(n_22388), .b(n_22387), .o(n_22389) );
in01f80 g547335 ( .a(n_21934), .o(n_21461) );
na02f80 g547336 ( .a(n_21122), .b(n_21121), .o(n_21934) );
no02f80 g547337 ( .a(n_21544), .b(n_21121), .o(n_20830) );
no02f80 g547338 ( .a(n_21119), .b(n_21118), .o(n_21120) );
no02f80 g547339 ( .a(n_21119), .b(n_20359), .o(n_22473) );
na02f80 g547340 ( .a(n_21459), .b(n_21458), .o(n_21460) );
in01f80 g547341 ( .a(n_22386), .o(n_23084) );
no02f80 g547342 ( .a(n_22124), .b(n_22116), .o(n_22386) );
na02f80 g547343 ( .a(n_21815), .b(n_22116), .o(n_21816) );
in01f80 g547344 ( .a(n_24281), .o(n_23919) );
oa12f80 g547345 ( .a(n_21451), .b(n_20793), .c(n_22607), .o(n_24281) );
in01f80 g547346 ( .a(n_24278), .o(n_23918) );
oa12f80 g547347 ( .a(n_21808), .b(n_21072), .c(n_22947), .o(n_24278) );
in01f80 g547348 ( .a(n_24273), .o(n_23917) );
oa12f80 g547349 ( .a(n_21798), .b(n_21070), .c(n_22946), .o(n_24273) );
in01f80 g547350 ( .a(n_24270), .o(n_23916) );
oa12f80 g547351 ( .a(n_21787), .b(n_21068), .c(n_22945), .o(n_24270) );
ao12f80 g547352 ( .a(n_23585), .b(n_21805), .c(n_23584), .o(n_24572) );
in01f80 g547353 ( .a(n_24012), .o(n_23600) );
oa12f80 g547354 ( .a(n_21450), .b(n_22606), .c(n_20785), .o(n_24012) );
in01f80 g547355 ( .a(n_23964), .o(n_23599) );
oa12f80 g547356 ( .a(n_21449), .b(n_22605), .c(n_20783), .o(n_23964) );
in01f80 g547357 ( .a(n_24009), .o(n_23598) );
oa12f80 g547358 ( .a(n_21448), .b(n_22593), .c(n_20781), .o(n_24009) );
in01f80 g547359 ( .a(n_23990), .o(n_23597) );
oa12f80 g547360 ( .a(n_21804), .b(n_22597), .c(n_21064), .o(n_23990) );
in01f80 g547361 ( .a(n_23596), .o(n_24567) );
oa12f80 g547362 ( .a(n_19973), .b(n_23260), .c(n_19313), .o(n_23596) );
in01f80 g547363 ( .a(n_24004), .o(n_24569) );
oa12f80 g547364 ( .a(n_21802), .b(n_21062), .c(n_22604), .o(n_24004) );
ao12f80 g547365 ( .a(n_13610), .b(n_20829), .c(n_14640), .o(n_21933) );
in01f80 g547366 ( .a(n_23273), .o(n_24220) );
oa12f80 g547367 ( .a(n_20943), .b(n_22971), .c(n_20218), .o(n_23273) );
in01f80 g547368 ( .a(n_23959), .o(n_23595) );
oa12f80 g547369 ( .a(n_21807), .b(n_21059), .c(n_22603), .o(n_23959) );
in01f80 g547370 ( .a(n_24252), .o(n_23915) );
oa12f80 g547371 ( .a(n_21435), .b(n_20777), .c(n_22944), .o(n_24252) );
in01f80 g547372 ( .a(n_24001), .o(n_23594) );
oa12f80 g547373 ( .a(n_21801), .b(n_21057), .c(n_22602), .o(n_24001) );
ao12f80 g547374 ( .a(n_23262), .b(n_23263), .c(n_21108), .o(n_24219) );
in01f80 g547375 ( .a(n_24255), .o(n_23914) );
oa12f80 g547376 ( .a(n_21444), .b(n_20772), .c(n_22941), .o(n_24255) );
in01f80 g547377 ( .a(n_24287), .o(n_23913) );
oa12f80 g547378 ( .a(n_21795), .b(n_21055), .c(n_22943), .o(n_24287) );
in01f80 g547379 ( .a(n_24262), .o(n_23912) );
oa12f80 g547380 ( .a(n_21786), .b(n_21053), .c(n_22942), .o(n_24262) );
ao12f80 g547381 ( .a(n_23258), .b(n_21794), .c(n_23257), .o(n_24218) );
in01f80 g547382 ( .a(n_23998), .o(n_23593) );
oa12f80 g547383 ( .a(n_21799), .b(n_21043), .c(n_22601), .o(n_23998) );
in01f80 g547384 ( .a(n_23995), .o(n_23592) );
oa12f80 g547385 ( .a(n_21800), .b(n_21045), .c(n_22600), .o(n_23995) );
in01f80 g547386 ( .a(n_23987), .o(n_23591) );
oa12f80 g547387 ( .a(n_21797), .b(n_21050), .c(n_22599), .o(n_23987) );
in01f80 g547388 ( .a(n_23272), .o(n_24216) );
oa12f80 g547389 ( .a(n_19355), .b(n_22969), .c(n_18668), .o(n_23272) );
oa12f80 g547390 ( .a(n_3249), .b(n_22383), .c(n_2261), .o(n_23373) );
oa12f80 g547391 ( .a(n_22366), .b(n_21706), .c(n_23245), .o(n_24900) );
in01f80 g547392 ( .a(n_24915), .o(n_24528) );
oa12f80 g547393 ( .a(n_21793), .b(n_21047), .c(n_23579), .o(n_24915) );
in01f80 g547394 ( .a(n_24249), .o(n_23911) );
oa12f80 g547395 ( .a(n_21443), .b(n_20768), .c(n_22940), .o(n_24249) );
in01f80 g547396 ( .a(n_23982), .o(n_23590) );
oa12f80 g547397 ( .a(n_21442), .b(n_20766), .c(n_22598), .o(n_23982) );
in01f80 g547398 ( .a(n_24246), .o(n_23910) );
oa12f80 g547399 ( .a(n_21441), .b(n_20764), .c(n_22939), .o(n_24246) );
in01f80 g547400 ( .a(n_23979), .o(n_23589) );
oa12f80 g547401 ( .a(n_21439), .b(n_20762), .c(n_22596), .o(n_23979) );
in01f80 g547402 ( .a(n_24243), .o(n_23909) );
oa12f80 g547403 ( .a(n_21440), .b(n_20759), .c(n_22938), .o(n_24243) );
in01f80 g547404 ( .a(n_22975), .o(n_23942) );
oa12f80 g547405 ( .a(n_17334), .b(n_22647), .c(n_16737), .o(n_22975) );
in01f80 g547406 ( .a(n_23687), .o(n_23271) );
oa12f80 g547407 ( .a(n_22365), .b(n_21692), .c(n_22296), .o(n_23687) );
in01f80 g547408 ( .a(n_23682), .o(n_23270) );
oa12f80 g547409 ( .a(n_22099), .b(n_21373), .c(n_22295), .o(n_23682) );
in01f80 g547410 ( .a(n_24240), .o(n_23908) );
oa12f80 g547411 ( .a(n_21436), .b(n_20753), .c(n_22937), .o(n_24240) );
in01f80 g547412 ( .a(n_22650), .o(n_23660) );
oa12f80 g547413 ( .a(n_3152), .b(n_22381), .c(n_2250), .o(n_22650) );
in01f80 g547414 ( .a(n_23588), .o(n_24565) );
oa12f80 g547415 ( .a(n_21628), .b(n_23252), .c(n_20934), .o(n_23588) );
in01f80 g547416 ( .a(n_23394), .o(n_22974) );
oa12f80 g547417 ( .a(n_22096), .b(n_21367), .c(n_22032), .o(n_23394) );
ao12f80 g547418 ( .a(n_23255), .b(n_21431), .c(n_23254), .o(n_24215) );
in01f80 g547419 ( .a(n_22649), .o(n_23658) );
oa12f80 g547420 ( .a(n_20424), .b(n_22378), .c(n_20020), .o(n_22649) );
ao12f80 g547421 ( .a(n_13624), .b(n_21117), .c(n_14271), .o(n_22195) );
in01f80 g547422 ( .a(n_24233), .o(n_23907) );
oa12f80 g547423 ( .a(n_21427), .b(n_22936), .c(n_20744), .o(n_24233) );
in01f80 g547424 ( .a(n_23269), .o(n_24213) );
oa12f80 g547425 ( .a(n_20261), .b(n_22967), .c(n_19536), .o(n_23269) );
in01f80 g547426 ( .a(n_24591), .o(n_24194) );
oa12f80 g547427 ( .a(n_22369), .b(n_21675), .c(n_23244), .o(n_24591) );
in01f80 g547428 ( .a(n_24230), .o(n_23906) );
oa12f80 g547429 ( .a(n_21426), .b(n_22935), .c(n_20740), .o(n_24230) );
in01f80 g547430 ( .a(n_24586), .o(n_25229) );
oa12f80 g547431 ( .a(n_22635), .b(n_22040), .c(n_23243), .o(n_24586) );
in01f80 g547432 ( .a(n_24583), .o(n_24193) );
oa12f80 g547433 ( .a(n_22355), .b(n_21669), .c(n_23242), .o(n_24583) );
in01f80 g547434 ( .a(n_24227), .o(n_23905) );
oa12f80 g547435 ( .a(n_21425), .b(n_22934), .c(n_20735), .o(n_24227) );
in01f80 g547436 ( .a(n_23388), .o(n_22973) );
oa12f80 g547437 ( .a(n_22090), .b(n_22031), .c(n_21350), .o(n_23388) );
ao12f80 g547438 ( .a(n_23250), .b(n_21784), .c(n_23249), .o(n_24212) );
in01f80 g547439 ( .a(n_23268), .o(n_24210) );
oa12f80 g547440 ( .a(n_22016), .b(n_22964), .c(n_21227), .o(n_23268) );
in01f80 g547441 ( .a(n_23267), .o(n_24208) );
oa12f80 g547442 ( .a(n_20923), .b(n_22962), .c(n_20203), .o(n_23267) );
in01f80 g547443 ( .a(n_24016), .o(n_23587) );
oa12f80 g547444 ( .a(n_21445), .b(n_22592), .c(n_20732), .o(n_24016) );
in01f80 g547445 ( .a(n_24265), .o(n_23904) );
oa12f80 g547446 ( .a(n_22100), .b(n_21346), .c(n_22933), .o(n_24265) );
in01f80 g547447 ( .a(n_24284), .o(n_23903) );
oa12f80 g547448 ( .a(n_22091), .b(n_21344), .c(n_22932), .o(n_24284) );
oa12f80 g547449 ( .a(n_10797), .b(n_21116), .c(n_12048), .o(n_22210) );
ao12f80 g547450 ( .a(n_10806), .b(n_20465), .c(n_12050), .o(n_21564) );
oa12f80 g547451 ( .a(n_12534), .b(n_19725), .c(n_11591), .o(n_20474) );
ao12f80 g547452 ( .a(n_20397), .b(n_23266), .c(n_21098), .o(n_24225) );
ao12f80 g547453 ( .a(n_20725), .b(n_23265), .c(n_21417), .o(n_24224) );
in01f80 g547454 ( .a(n_23377), .o(n_23656) );
ao12f80 g547455 ( .a(n_16912), .b(n_22385), .c(n_17299), .o(n_23377) );
ao12f80 g547456 ( .a(n_13616), .b(n_20828), .c(n_14646), .o(n_21931) );
ao12f80 g547457 ( .a(n_8311), .b(n_20827), .c(n_9527), .o(n_21932) );
ao12f80 g547458 ( .a(n_21422), .b(n_21421), .c(n_21420), .o(n_22115) );
in01f80 g547459 ( .a(n_21554), .o(n_21918) );
ao12f80 g547460 ( .a(n_20106), .b(n_20465), .c(n_20105), .o(n_21554) );
oa12f80 g547461 ( .a(n_21806), .b(n_23585), .c(n_23584), .o(n_23586) );
oa12f80 g547462 ( .a(n_21109), .b(n_23263), .c(n_23262), .o(n_23264) );
ao12f80 g547463 ( .a(n_20455), .b(n_20456), .c(n_20454), .o(n_21115) );
in01f80 g547464 ( .a(n_21920), .o(n_22188) );
ao12f80 g547465 ( .a(n_20462), .b(n_20829), .c(n_20461), .o(n_21920) );
oa12f80 g547466 ( .a(n_20816), .b(n_20826), .c(n_21096), .o(n_22191) );
ao22s80 g547467 ( .a(n_20305), .b(n_23260), .c(n_20304), .d(n_22595), .o(n_23261) );
ao22s80 g547468 ( .a(n_22971), .b(n_21259), .c(n_22298), .d(n_21258), .o(n_22972) );
oa12f80 g547469 ( .a(n_21803), .b(n_23258), .c(n_23257), .o(n_23259) );
ao22s80 g547470 ( .a(n_22969), .b(n_19626), .c(n_22297), .d(n_19625), .o(n_22970) );
ao22s80 g547471 ( .a(n_22383), .b(n_4119), .c(n_21654), .d(n_4118), .o(n_22384) );
in01f80 g547472 ( .a(n_22184), .o(n_22449) );
ao12f80 g547473 ( .a(n_20825), .b(n_21116), .c(n_20824), .o(n_22184) );
ao22s80 g547474 ( .a(n_22381), .b(n_4087), .c(n_21653), .d(n_4086), .o(n_22382) );
ao22s80 g547475 ( .a(n_22647), .b(n_17564), .c(n_22033), .d(n_17563), .o(n_22648) );
ao12f80 g547476 ( .a(n_21438), .b(n_21810), .c(n_21437), .o(n_22114) );
in01f80 g547477 ( .a(n_20107), .o(n_21190) );
oa22f80 g547478 ( .a(n_19725), .b(n_12948), .c(n_19064), .d(n_12949), .o(n_20107) );
ao12f80 g547479 ( .a(n_21783), .b(n_22109), .c(n_21782), .o(n_22380) );
in01f80 g547480 ( .a(n_22438), .o(n_22734) );
ao12f80 g547481 ( .a(n_21107), .b(n_21465), .c(n_21106), .o(n_22438) );
in01f80 g547482 ( .a(n_23070), .o(n_23347) );
oa12f80 g547483 ( .a(n_21792), .b(n_21791), .c(n_21790), .o(n_23070) );
oa12f80 g547484 ( .a(n_21434), .b(n_23255), .c(n_23254), .o(n_23256) );
ao12f80 g547485 ( .a(n_21102), .b(FE_OFN818_n_20821), .c(n_21100), .o(n_21814) );
in01f80 g547486 ( .a(n_21457), .o(n_22468) );
oa12f80 g547487 ( .a(n_20460), .b(n_20827), .c(n_20459), .o(n_21457) );
oa12f80 g547488 ( .a(n_21419), .b(n_21781), .c(n_21418), .o(n_22738) );
ao12f80 g547489 ( .a(n_21414), .b(n_21413), .c(n_21412), .o(n_22113) );
in01f80 g547490 ( .a(n_22172), .o(n_21813) );
oa12f80 g547491 ( .a(n_20823), .b(n_21117), .c(n_20822), .o(n_22172) );
ao22s80 g547492 ( .a(n_23252), .b(n_22015), .c(n_22594), .d(n_22014), .o(n_23253) );
in01f80 g547493 ( .a(n_21812), .o(n_22752) );
oa12f80 g547494 ( .a(n_20820), .b(n_21130), .c(n_20819), .o(n_21812) );
ao22s80 g547495 ( .a(n_20747), .b(n_22378), .c(n_20746), .d(n_21652), .o(n_22379) );
in01f80 g547496 ( .a(n_21925), .o(n_21456) );
oa12f80 g547497 ( .a(n_20458), .b(n_20828), .c(n_20457), .o(n_21925) );
ao12f80 g547498 ( .a(n_22093), .b(n_22385), .c(n_22092), .o(n_22646) );
ao22s80 g547499 ( .a(n_20577), .b(n_22967), .c(n_20576), .d(n_22294), .o(n_22968) );
oa12f80 g547500 ( .a(n_21785), .b(n_23250), .c(n_23249), .o(n_23251) );
ao12f80 g547501 ( .a(n_19723), .b(n_19722), .c(n_19721), .o(n_20464) );
in01f80 g547502 ( .a(n_23352), .o(n_22966) );
oa12f80 g547503 ( .a(n_22088), .b(n_22352), .c(n_22373), .o(n_23352) );
ao22s80 g547504 ( .a(n_22964), .b(n_22283), .c(n_22293), .d(n_22282), .o(n_22965) );
oa12f80 g547505 ( .a(n_20818), .b(n_20817), .c(n_21097), .o(n_22178) );
ao22s80 g547506 ( .a(n_22962), .b(n_21221), .c(n_22292), .d(n_21220), .o(n_22963) );
oa22f80 g547507 ( .a(n_21335), .b(n_22960), .c(n_1835), .d(FE_OFN122_n_27449), .o(n_22112) );
oa22f80 g547508 ( .a(n_20356), .b(FE_OFN412_n_28303), .c(n_1830), .d(FE_OFN329_n_4860), .o(n_21114) );
oa22f80 g547509 ( .a(n_22109), .b(n_22960), .c(n_201), .d(FE_OFN324_n_4860), .o(n_22110) );
oa22f80 g547510 ( .a(n_20705), .b(FE_OFN300_n_3069), .c(n_670), .d(n_29617), .o(n_21455) );
oa22f80 g547511 ( .a(n_22291), .b(n_22960), .c(n_1874), .d(FE_OFN63_n_27012), .o(n_22961) );
oa22f80 g547512 ( .a(n_22029), .b(FE_OFN230_n_4162), .c(n_312), .d(n_25680), .o(n_22645) );
oa22f80 g547513 ( .a(FE_OFN819_n_20821), .b(n_22960), .c(n_1778), .d(n_25680), .o(n_21113) );
oa22f80 g547514 ( .a(n_21099), .b(FE_OFN166_n_29269), .c(n_1655), .d(FE_OFN335_n_4860), .o(n_21454) );
oa22f80 g547515 ( .a(n_21095), .b(FE_OFN165_n_29269), .c(n_615), .d(FE_OFN72_n_27012), .o(n_21453) );
oa22f80 g547516 ( .a(FE_OFN664_n_22027), .b(n_22960), .c(n_1609), .d(n_25680), .o(n_22644) );
oa22f80 g547517 ( .a(FE_OFN462_n_21334), .b(n_21076), .c(n_579), .d(FE_OFN1108_rst), .o(n_22108) );
oa22f80 g547518 ( .a(n_21810), .b(n_21076), .c(n_582), .d(n_27449), .o(n_21811) );
oa22f80 g547519 ( .a(n_21651), .b(FE_OFN295_n_3069), .c(n_1937), .d(FE_OFN130_n_27449), .o(n_22377) );
oa22f80 g547520 ( .a(n_21331), .b(FE_OFN295_n_3069), .c(n_485), .d(FE_OFN76_n_27012), .o(n_22107) );
oa22f80 g547521 ( .a(n_21332), .b(FE_OFN297_n_3069), .c(n_572), .d(FE_OFN141_n_27449), .o(n_22106) );
oa22f80 g547522 ( .a(n_19396), .b(FE_OFN166_n_29269), .c(n_542), .d(FE_OFN1143_n_27012), .o(n_19724) );
oa22f80 g547523 ( .a(n_21649), .b(n_29269), .c(n_1954), .d(FE_OFN77_n_27012), .o(n_22376) );
oa22f80 g547524 ( .a(FE_OFN496_n_21648), .b(n_29046), .c(n_535), .d(n_27449), .o(n_22375) );
oa22f80 g547525 ( .a(n_20704), .b(FE_OFN312_n_3069), .c(n_1735), .d(FE_OFN92_n_27449), .o(n_21452) );
oa22f80 g547526 ( .a(n_21012), .b(FE_OFN306_n_3069), .c(n_492), .d(FE_OFN94_n_27449), .o(n_21809) );
oa22f80 g547527 ( .a(n_22373), .b(FE_OFN312_n_3069), .c(n_1638), .d(FE_OFN113_n_27449), .o(n_22374) );
oa22f80 g547528 ( .a(n_22289), .b(FE_OFN312_n_3069), .c(n_501), .d(FE_OFN330_n_4860), .o(n_22959) );
oa22f80 g547529 ( .a(n_21328), .b(FE_OFN314_n_3069), .c(n_79), .d(FE_OFN330_n_4860), .o(n_22105) );
oa22f80 g547530 ( .a(n_21646), .b(FE_OFN308_n_3069), .c(n_399), .d(FE_OFN114_n_27449), .o(n_22371) );
oa22f80 g547531 ( .a(FE_OFN684_n_22025), .b(n_23813), .c(n_202), .d(FE_OFN102_n_27449), .o(n_22643) );
oa22f80 g547532 ( .a(n_19676), .b(n_23813), .c(n_812), .d(FE_OFN1118_rst), .o(n_20463) );
oa22f80 g547533 ( .a(n_22287), .b(n_23813), .c(n_310), .d(n_25680), .o(n_22958) );
oa22f80 g547534 ( .a(n_22286), .b(FE_OFN219_n_23315), .c(n_1676), .d(FE_OFN1111_rst), .o(n_22957) );
oa22f80 g547535 ( .a(n_22023), .b(FE_OFN221_n_23315), .c(n_1686), .d(FE_OFN1123_rst), .o(n_22642) );
na02f80 g547565 ( .a(n_21808), .b(n_21073), .o(n_23038) );
na02f80 g547566 ( .a(n_21451), .b(n_20794), .o(n_23041) );
na02f80 g547567 ( .a(n_22369), .b(n_21676), .o(n_23284) );
na02f80 g547568 ( .a(n_21807), .b(n_21060), .o(n_22715) );
in01f80 g547569 ( .a(n_22640), .o(n_22641) );
na02f80 g547570 ( .a(n_22368), .b(n_21755), .o(n_22640) );
no02f80 g547571 ( .a(n_21066), .b(x_in_6_7), .o(n_21806) );
na02f80 g547572 ( .a(n_21450), .b(n_20786), .o(n_22718) );
in01f80 g547573 ( .a(n_22103), .o(n_22104) );
no02f80 g547574 ( .a(n_22400), .b(x_in_24_12), .o(n_22103) );
na02f80 g547575 ( .a(n_21449), .b(n_20784), .o(n_22666) );
na02f80 g547576 ( .a(n_21805), .b(n_21067), .o(n_22986) );
na02f80 g547577 ( .a(n_20826), .b(x_in_38_10), .o(n_21886) );
na02f80 g547578 ( .a(n_21448), .b(n_20782), .o(n_22724) );
in01f80 g547579 ( .a(n_21111), .o(n_21112) );
no02f80 g547580 ( .a(n_20826), .b(x_in_38_10), .o(n_21111) );
na02f80 g547581 ( .a(n_21804), .b(n_21065), .o(n_22709) );
na02f80 g547582 ( .a(n_21110), .b(x_in_38_9), .o(n_22125) );
in01f80 g547583 ( .a(n_21446), .o(n_21447) );
no02f80 g547584 ( .a(n_21110), .b(x_in_38_9), .o(n_21446) );
in01f80 g547585 ( .a(n_22101), .o(n_22102) );
no02f80 g547586 ( .a(n_21796), .b(x_in_24_11), .o(n_22101) );
no02f80 g547587 ( .a(n_20435), .b(x_in_52_7), .o(n_21109) );
na02f80 g547588 ( .a(n_21445), .b(n_20733), .o(n_22727) );
no02f80 g547589 ( .a(n_21052), .b(x_in_14_7), .o(n_21803) );
na02f80 g547590 ( .a(n_21802), .b(n_21063), .o(n_22721) );
na02f80 g547591 ( .a(n_21801), .b(n_21058), .o(n_22712) );
na02f80 g547592 ( .a(n_21800), .b(n_21046), .o(n_22700) );
na02f80 g547593 ( .a(n_21799), .b(n_21044), .o(n_22703) );
na02f80 g547594 ( .a(n_21798), .b(n_21071), .o(n_23035) );
na02f80 g547595 ( .a(n_21797), .b(n_21051), .o(n_22688) );
na02f80 g547596 ( .a(n_21796), .b(x_in_24_11), .o(n_22698) );
na02f80 g547597 ( .a(n_22400), .b(x_in_24_12), .o(n_22697) );
na02f80 g547598 ( .a(n_21444), .b(n_20773), .o(n_22992) );
in01f80 g547599 ( .a(n_22638), .o(n_22639) );
na02f80 g547600 ( .a(n_22367), .b(n_21712), .o(n_22638) );
na02f80 g547601 ( .a(n_21795), .b(n_21056), .o(n_23023) );
na02f80 g547602 ( .a(n_21794), .b(n_21037), .o(n_22706) );
na02f80 g547603 ( .a(n_22366), .b(n_21707), .o(n_23287) );
na02f80 g547604 ( .a(n_21443), .b(n_20769), .o(n_23009) );
na02f80 g547605 ( .a(n_21108), .b(n_20422), .o(n_22694) );
no02f80 g547606 ( .a(n_20829), .b(n_20461), .o(n_20462) );
na02f80 g547607 ( .a(n_21793), .b(n_21048), .o(n_23606) );
no02f80 g547608 ( .a(n_21116), .b(n_20824), .o(n_20825) );
na02f80 g547609 ( .a(n_21442), .b(n_20767), .o(n_22691) );
na02f80 g547610 ( .a(n_21441), .b(n_20765), .o(n_23006) );
na02f80 g547611 ( .a(n_22100), .b(n_21347), .o(n_23029) );
na02f80 g547612 ( .a(n_21440), .b(n_20760), .o(n_23003) );
na02f80 g547613 ( .a(n_21439), .b(n_20763), .o(n_22685) );
na02f80 g547614 ( .a(n_22365), .b(n_21693), .o(n_23000) );
no02f80 g547615 ( .a(n_21810), .b(n_21437), .o(n_21438) );
no02f80 g547616 ( .a(n_21013), .b(n_21437), .o(n_22448) );
na02f80 g547617 ( .a(n_22099), .b(n_21374), .o(n_22682) );
na02f80 g547618 ( .a(n_22362), .b(x_in_44_9), .o(n_23282) );
in01f80 g547619 ( .a(n_22363), .o(n_22364) );
na02f80 g547620 ( .a(n_22098), .b(n_21372), .o(n_22363) );
in01f80 g547621 ( .a(n_22636), .o(n_22637) );
no02f80 g547622 ( .a(n_22362), .b(x_in_44_9), .o(n_22636) );
na02f80 g547623 ( .a(n_21436), .b(n_20754), .o(n_22995) );
no02f80 g547624 ( .a(n_21465), .b(n_21106), .o(n_21107) );
in01f80 g547625 ( .a(n_22360), .o(n_22361) );
na02f80 g547626 ( .a(n_22097), .b(n_21370), .o(n_22360) );
na02f80 g547627 ( .a(n_21435), .b(n_20778), .o(n_23014) );
no02f80 g547628 ( .a(n_20750), .b(x_in_32_7), .o(n_21434) );
na02f80 g547629 ( .a(n_21791), .b(n_21790), .o(n_21792) );
na02f80 g547630 ( .a(n_22096), .b(n_21368), .o(n_22677) );
na02f80 g547631 ( .a(n_21105), .b(x_in_24_9), .o(n_22129) );
in01f80 g547632 ( .a(n_21432), .o(n_21433) );
no02f80 g547633 ( .a(n_21105), .b(x_in_24_9), .o(n_21432) );
na02f80 g547634 ( .a(n_21117), .b(n_20822), .o(n_20823) );
na02f80 g547635 ( .a(n_21431), .b(n_20751), .o(n_22674) );
in01f80 g547636 ( .a(n_21788), .o(n_21789) );
na02f80 g547637 ( .a(n_21430), .b(n_20749), .o(n_21788) );
na02f80 g547638 ( .a(n_21104), .b(x_in_28_10), .o(n_22128) );
na02f80 g547639 ( .a(n_21787), .b(n_21069), .o(n_23032) );
in01f80 g547640 ( .a(n_21428), .o(n_21429) );
no02f80 g547641 ( .a(n_21104), .b(x_in_28_10), .o(n_21428) );
in01f80 g547642 ( .a(n_22358), .o(n_22359) );
na02f80 g547643 ( .a(n_22095), .b(n_21360), .o(n_22358) );
na02f80 g547644 ( .a(n_21427), .b(n_20745), .o(n_22989) );
in01f80 g547645 ( .a(n_22356), .o(n_22357) );
na02f80 g547646 ( .a(n_22094), .b(n_21358), .o(n_22356) );
no02f80 g547647 ( .a(n_22385), .b(n_22092), .o(n_22093) );
na02f80 g547648 ( .a(n_21426), .b(n_20741), .o(n_22981) );
na02f80 g547649 ( .a(n_22635), .b(n_22041), .o(n_23279) );
na02f80 g547650 ( .a(n_22091), .b(n_21345), .o(n_23044) );
na02f80 g547651 ( .a(n_22355), .b(n_21670), .o(n_23276) );
na02f80 g547652 ( .a(n_21786), .b(n_21054), .o(n_23026) );
na02f80 g547653 ( .a(n_22090), .b(n_21351), .o(n_22661) );
no02f80 g547654 ( .a(n_21030), .b(x_in_12_7), .o(n_21785) );
na02f80 g547655 ( .a(n_21425), .b(n_20736), .o(n_22978) );
no02f80 g547656 ( .a(n_19722), .b(n_19721), .o(n_19723) );
na02f80 g547657 ( .a(n_19396), .b(n_19721), .o(n_20876) );
na02f80 g547658 ( .a(n_21784), .b(n_21031), .o(n_22658) );
na02f80 g547659 ( .a(n_22354), .b(x_in_44_8), .o(n_23274) );
in01f80 g547660 ( .a(n_22633), .o(n_22634) );
no02f80 g547661 ( .a(n_22354), .b(x_in_44_8), .o(n_22633) );
in01f80 g547662 ( .a(n_22631), .o(n_22632) );
na02f80 g547663 ( .a(n_22353), .b(n_21659), .o(n_22631) );
na02f80 g547664 ( .a(n_21103), .b(x_in_28_9), .o(n_22123) );
in01f80 g547665 ( .a(n_21423), .o(n_21424) );
no02f80 g547666 ( .a(n_21103), .b(x_in_28_9), .o(n_21423) );
no02f80 g547667 ( .a(n_20465), .b(n_20105), .o(n_20106) );
no02f80 g547668 ( .a(n_22109), .b(n_21782), .o(n_21783) );
no02f80 g547669 ( .a(n_21329), .b(n_21782), .o(n_22733) );
no02f80 g547670 ( .a(FE_OFN818_n_20821), .b(n_21100), .o(n_21102) );
na02f80 g547671 ( .a(n_20821), .b(n_21100), .o(n_22176) );
na02f80 g547672 ( .a(n_21130), .b(n_20819), .o(n_20820) );
in01f80 g547673 ( .a(n_22089), .o(n_23059) );
na02f80 g547674 ( .a(n_21780), .b(n_11463), .o(n_22089) );
na02f80 g547675 ( .a(n_21099), .b(n_21420), .o(n_22436) );
no02f80 g547676 ( .a(n_21421), .b(n_21420), .o(n_21422) );
na02f80 g547677 ( .a(n_21781), .b(n_21418), .o(n_21419) );
no02f80 g547678 ( .a(n_21781), .b(n_21796), .o(n_22401) );
na02f80 g547679 ( .a(n_20396), .b(n_21098), .o(n_23011) );
na02f80 g547680 ( .a(n_20724), .b(n_21417), .o(n_22997) );
no02f80 g547681 ( .a(n_22352), .b(n_22362), .o(n_23348) );
na02f80 g547682 ( .a(n_22352), .b(n_22373), .o(n_22088) );
na02f80 g547683 ( .a(n_20817), .b(n_21097), .o(n_20818) );
no02f80 g547684 ( .a(n_21104), .b(n_21097), .o(n_22175) );
na02f80 g547685 ( .a(n_20827), .b(n_20459), .o(n_20460) );
na02f80 g547686 ( .a(n_20828), .b(n_20457), .o(n_20458) );
na02f80 g547687 ( .a(n_20706), .b(n_21096), .o(n_22174) );
na02f80 g547688 ( .a(n_20826), .b(n_21096), .o(n_20816) );
no02f80 g547689 ( .a(n_20456), .b(n_20008), .o(n_21917) );
no02f80 g547690 ( .a(n_20456), .b(n_20454), .o(n_20455) );
in01f80 g547691 ( .a(n_22427), .o(n_22087) );
oa12f80 g547692 ( .a(n_21780), .b(n_21039), .c(n_12547), .o(n_22427) );
na03f80 g547693 ( .a(n_10833), .b(n_21465), .c(n_21415), .o(n_21416) );
oa12f80 g547694 ( .a(n_21023), .b(n_8014), .c(n_8013), .o(n_22732) );
no02f80 g547695 ( .a(n_21413), .b(n_21412), .o(n_21414) );
in01f80 g547696 ( .a(n_21411), .o(n_22171) );
na02f80 g547697 ( .a(n_21095), .b(n_21412), .o(n_21411) );
in01f80 g547698 ( .a(n_23247), .o(n_24203) );
oa12f80 g547699 ( .a(n_21005), .b(n_22953), .c(n_20273), .o(n_23247) );
oa12f80 g547700 ( .a(n_13216), .b(n_20453), .c(n_14249), .o(n_21551) );
oa12f80 g547701 ( .a(n_16126), .b(n_20452), .c(n_16690), .o(n_21552) );
ao12f80 g547702 ( .a(n_15559), .b(n_19720), .c(n_16263), .o(n_20874) );
oa12f80 g547703 ( .a(n_15415), .b(n_20451), .c(n_14636), .o(n_21550) );
oa12f80 g547704 ( .a(n_15412), .b(n_20104), .c(n_14765), .o(n_21187) );
in01f80 g547705 ( .a(n_22630), .o(n_23623) );
oa12f80 g547706 ( .a(n_21311), .b(n_20622), .c(n_22318), .o(n_22630) );
oa12f80 g547707 ( .a(n_15398), .b(n_20103), .c(n_14742), .o(n_21185) );
oa12f80 g547708 ( .a(n_14382), .b(n_20102), .c(n_15143), .o(n_21184) );
ao12f80 g547709 ( .a(n_14715), .b(n_20101), .c(n_15386), .o(n_21183) );
oa12f80 g547710 ( .a(n_15368), .b(n_20100), .c(n_14688), .o(n_21182) );
in01f80 g547711 ( .a(n_22086), .o(n_23061) );
oa12f80 g547712 ( .a(n_21308), .b(n_21779), .c(n_20602), .o(n_22086) );
oa12f80 g547713 ( .a(n_13154), .b(n_20450), .c(n_14316), .o(n_21549) );
in01f80 g547714 ( .a(n_22955), .o(n_23925) );
oa12f80 g547715 ( .a(n_20996), .b(n_22623), .c(n_20275), .o(n_22955) );
ao12f80 g547716 ( .a(n_16102), .b(n_21094), .c(n_16681), .o(n_22170) );
oa12f80 g547717 ( .a(n_15408), .b(n_20099), .c(n_14797), .o(n_21186) );
in01f80 g547718 ( .a(n_22085), .o(n_23058) );
ao12f80 g547719 ( .a(n_11020), .b(n_21776), .c(n_12122), .o(n_22085) );
in01f80 g547720 ( .a(n_22629), .o(n_23621) );
oa12f80 g547721 ( .a(n_20994), .b(n_20265), .c(n_22324), .o(n_22629) );
in01f80 g547722 ( .a(n_22628), .o(n_23618) );
oa12f80 g547723 ( .a(n_21300), .b(n_22321), .c(n_20585), .o(n_22628) );
ao12f80 g547724 ( .a(n_15503), .b(n_21093), .c(n_16251), .o(n_22169) );
oa12f80 g547725 ( .a(n_10643), .b(n_20098), .c(n_11781), .o(n_21180) );
oa12f80 g547726 ( .a(n_11425), .b(n_20097), .c(n_12478), .o(n_21181) );
oa12f80 g547727 ( .a(n_14288), .b(n_20096), .c(n_15084), .o(n_21179) );
ao12f80 g547728 ( .a(n_15373), .b(n_20449), .c(n_14702), .o(n_21548) );
ao12f80 g547729 ( .a(n_12276), .b(n_19719), .c(n_12491), .o(n_20873) );
oa12f80 g547730 ( .a(n_14351), .b(n_20095), .c(n_15132), .o(n_21178) );
oa12f80 g547731 ( .a(n_16087), .b(n_20815), .c(n_16688), .o(n_21914) );
oa12f80 g547732 ( .a(n_14307), .b(n_20448), .c(n_15114), .o(n_21547) );
ao12f80 g547733 ( .a(n_13651), .b(n_20094), .c(n_14402), .o(n_21177) );
ao12f80 g547734 ( .a(n_8327), .b(n_20447), .c(n_8954), .o(n_21553) );
oa12f80 g547735 ( .a(n_13185), .b(n_21092), .c(n_14366), .o(n_22168) );
ao12f80 g547736 ( .a(n_13997), .b(n_20093), .c(n_14961), .o(n_21176) );
ao12f80 g547737 ( .a(n_14419), .b(n_20446), .c(n_15156), .o(n_21546) );
ao12f80 g547738 ( .a(n_11446), .b(n_19718), .c(n_11789), .o(n_20872) );
oa12f80 g547739 ( .a(n_13164), .b(n_20814), .c(n_14328), .o(n_21913) );
oa12f80 g547740 ( .a(n_13923), .b(n_20092), .c(n_14915), .o(n_21175) );
oa12f80 g547741 ( .a(n_13901), .b(n_20091), .c(n_14911), .o(n_21174) );
oa12f80 g547742 ( .a(n_11479), .b(n_20445), .c(n_12458), .o(n_21545) );
oa22f80 g547743 ( .a(n_20985), .b(n_7110), .c(n_3600), .d(n_21777), .o(n_21778) );
oa12f80 g547744 ( .a(n_15524), .b(n_20090), .c(n_16255), .o(n_21173) );
oa12f80 g547745 ( .a(n_13974), .b(n_20089), .c(n_14906), .o(n_21172) );
ao12f80 g547746 ( .a(n_13959), .b(n_20088), .c(n_14933), .o(n_21171) );
oa12f80 g547747 ( .a(n_10683), .b(n_20087), .c(n_11800), .o(n_21169) );
ao12f80 g547748 ( .a(n_8319), .b(n_20086), .c(n_8950), .o(n_21170) );
ao12f80 g547749 ( .a(n_21727), .b(n_21726), .c(n_21725), .o(n_22351) );
ao12f80 g547750 ( .a(n_20721), .b(n_20720), .c(n_20719), .o(n_21410) );
in01f80 g547751 ( .a(FE_OFN632_n_21154), .o(n_21507) );
ao12f80 g547752 ( .a(n_19717), .b(n_20097), .c(n_19716), .o(n_21154) );
ao12f80 g547753 ( .a(n_21764), .b(n_21763), .c(n_21762), .o(n_22350) );
oa12f80 g547754 ( .a(n_20373), .b(n_20372), .c(n_20371), .o(n_21897) );
ao12f80 g547755 ( .a(n_21761), .b(n_21760), .c(n_21759), .o(n_22349) );
oa12f80 g547756 ( .a(n_20718), .b(n_20717), .c(n_20716), .o(n_22150) );
ao12f80 g547757 ( .a(n_22048), .b(n_22047), .c(n_22046), .o(n_22627) );
ao12f80 g547758 ( .a(n_21342), .b(n_21768), .c(n_21341), .o(n_22084) );
ao12f80 g547759 ( .a(n_21758), .b(n_21757), .c(n_21756), .o(n_22348) );
ao22s80 g547760 ( .a(n_21319), .b(n_22953), .c(n_21318), .d(n_22281), .o(n_22954) );
oa12f80 g547761 ( .a(n_20052), .b(n_20051), .c(n_20394), .o(n_21537) );
ao12f80 g547762 ( .a(n_20790), .b(n_21081), .c(n_20789), .o(n_21409) );
ao12f80 g547763 ( .a(n_21753), .b(n_21752), .c(n_21751), .o(n_22347) );
oa12f80 g547764 ( .a(n_20033), .b(n_20032), .c(n_20393), .o(n_21536) );
ao12f80 g547765 ( .a(n_20383), .b(n_20392), .c(n_20382), .o(n_21091) );
in01f80 g547766 ( .a(n_21477), .o(n_22433) );
ao12f80 g547767 ( .a(n_20083), .b(n_20452), .c(n_20082), .o(n_21477) );
ao12f80 g547768 ( .a(n_21747), .b(n_21746), .c(n_21745), .o(n_22346) );
oa12f80 g547769 ( .a(n_20376), .b(n_20375), .c(n_20374), .o(n_21889) );
ao12f80 g547770 ( .a(n_21397), .b(n_21396), .c(n_21395), .o(n_22083) );
oa12f80 g547771 ( .a(n_20391), .b(n_20390), .c(n_20389), .o(n_21888) );
ao12f80 g547772 ( .a(n_21355), .b(n_21354), .c(n_21353), .o(n_22082) );
in01f80 g547773 ( .a(n_21487), .o(n_21090) );
oa12f80 g547774 ( .a(n_20081), .b(n_20453), .c(n_20080), .o(n_21487) );
oa12f80 g547775 ( .a(n_20388), .b(n_20387), .c(n_20386), .o(n_21887) );
ao12f80 g547776 ( .a(n_21744), .b(n_21743), .c(n_21742), .o(n_22345) );
ao12f80 g547777 ( .a(n_21741), .b(n_21740), .c(n_21739), .o(n_22344) );
in01f80 g547778 ( .a(n_21815), .o(n_22124) );
ao12f80 g547779 ( .a(n_20413), .b(n_20815), .c(n_20412), .o(n_21815) );
oa12f80 g547780 ( .a(n_20049), .b(n_20048), .c(n_20378), .o(n_21528) );
ao12f80 g547781 ( .a(n_21377), .b(n_21376), .c(n_21375), .o(n_22081) );
oa12f80 g547782 ( .a(n_20385), .b(n_20384), .c(n_20708), .o(n_21851) );
ao12f80 g547783 ( .a(n_21403), .b(n_21402), .c(n_21401), .o(n_22080) );
ao12f80 g547784 ( .a(n_21750), .b(n_21749), .c(n_21748), .o(n_22343) );
in01f80 g547785 ( .a(n_21135), .o(n_21505) );
ao12f80 g547786 ( .a(n_19695), .b(n_20093), .c(n_19694), .o(n_21135) );
oa12f80 g547787 ( .a(n_20066), .b(n_20065), .c(n_20410), .o(n_21534) );
in01f80 g547788 ( .a(n_21533), .o(n_21089) );
oa12f80 g547789 ( .a(n_20079), .b(n_20451), .c(n_20078), .o(n_21533) );
ao12f80 g547790 ( .a(n_21730), .b(n_21729), .c(n_21728), .o(n_22342) );
oa12f80 g547791 ( .a(n_20402), .b(n_20401), .c(n_20400), .o(n_22591) );
ao12f80 g547792 ( .a(n_21724), .b(n_21723), .c(n_21722), .o(n_22341) );
ao12f80 g547793 ( .a(n_21721), .b(n_21720), .c(n_21719), .o(n_22340) );
oa12f80 g547794 ( .a(n_20064), .b(n_20063), .c(n_20408), .o(n_21532) );
in01f80 g547795 ( .a(n_21162), .o(n_20813) );
oa12f80 g547796 ( .a(n_19715), .b(n_20104), .c(n_19714), .o(n_21162) );
oa12f80 g547797 ( .a(n_20062), .b(n_20061), .c(n_20411), .o(n_21529) );
ao12f80 g547798 ( .a(n_21733), .b(n_21732), .c(n_21731), .o(n_22339) );
ao12f80 g547799 ( .a(n_21718), .b(n_21717), .c(n_21716), .o(n_22338) );
ao12f80 g547800 ( .a(n_21710), .b(n_21709), .c(n_21708), .o(n_22337) );
ao12f80 g547801 ( .a(n_22036), .b(n_22035), .c(n_22034), .o(n_22626) );
in01f80 g547802 ( .a(n_21161), .o(n_20812) );
oa12f80 g547803 ( .a(n_19713), .b(n_20099), .c(n_19712), .o(n_21161) );
ao12f80 g547804 ( .a(n_21705), .b(n_21704), .c(n_21703), .o(n_22336) );
in01f80 g547805 ( .a(n_21119), .o(n_20811) );
oa12f80 g547806 ( .a(n_19697), .b(n_20094), .c(n_19696), .o(n_21119) );
in01f80 g547807 ( .a(n_21475), .o(n_21873) );
ao12f80 g547808 ( .a(n_20068), .b(n_20446), .c(n_20067), .o(n_21475) );
in01f80 g547809 ( .a(n_21160), .o(n_20810) );
oa12f80 g547810 ( .a(n_19711), .b(n_20103), .c(n_19710), .o(n_21160) );
ao12f80 g547811 ( .a(n_21715), .b(n_21714), .c(n_21713), .o(n_22335) );
ao12f80 g547812 ( .a(n_21702), .b(n_21701), .c(n_21700), .o(n_22334) );
in01f80 g547813 ( .a(n_21471), .o(n_21523) );
ao12f80 g547814 ( .a(n_19709), .b(n_20102), .c(n_19708), .o(n_21471) );
ao12f80 g547815 ( .a(n_21387), .b(n_21386), .c(n_21385), .o(n_22079) );
in01f80 g547816 ( .a(n_22122), .o(n_22398) );
ao12f80 g547817 ( .a(n_20731), .b(n_21092), .c(n_20730), .o(n_22122) );
ao12f80 g547818 ( .a(n_22306), .b(n_22305), .c(n_22304), .o(n_22952) );
ao12f80 g547819 ( .a(n_21384), .b(n_21383), .c(n_21382), .o(n_22078) );
in01f80 g547820 ( .a(n_21159), .o(n_20809) );
oa12f80 g547821 ( .a(n_19707), .b(n_20101), .c(n_19706), .o(n_21159) );
in01f80 g547822 ( .a(n_21463), .o(n_21520) );
ao12f80 g547823 ( .a(n_19699), .b(n_20095), .c(n_19698), .o(n_21463) );
ao12f80 g547824 ( .a(n_21699), .b(n_21698), .c(n_21697), .o(n_22333) );
in01f80 g547825 ( .a(n_21519), .o(n_21088) );
oa12f80 g547826 ( .a(n_20074), .b(n_20449), .c(n_20073), .o(n_21519) );
ao12f80 g547827 ( .a(n_21391), .b(n_21390), .c(n_21389), .o(n_22077) );
in01f80 g547828 ( .a(n_21158), .o(n_20808) );
oa12f80 g547829 ( .a(n_19705), .b(n_20100), .c(n_19704), .o(n_21158) );
ao12f80 g547830 ( .a(n_21696), .b(n_21695), .c(n_21694), .o(n_22332) );
in01f80 g547831 ( .a(FE_OFN604_n_21535), .o(n_21893) );
ao12f80 g547832 ( .a(n_20057), .b(n_20445), .c(n_20056), .o(n_21535) );
oa12f80 g547833 ( .a(n_20060), .b(n_20059), .c(n_20409), .o(n_21504) );
ao12f80 g547834 ( .a(n_21381), .b(n_21380), .c(n_21379), .o(n_22076) );
oa12f80 g547835 ( .a(n_20380), .b(n_20379), .c(n_20381), .o(n_21866) );
ao12f80 g547836 ( .a(n_20047), .b(n_20046), .c(n_20045), .o(n_20807) );
ao12f80 g547837 ( .a(n_22045), .b(n_22044), .c(n_22043), .o(n_22625) );
oa12f80 g547838 ( .a(n_20043), .b(n_20042), .c(n_20377), .o(n_21516) );
ao12f80 g547839 ( .a(n_21691), .b(n_21690), .c(n_21689), .o(n_22331) );
in01f80 g547840 ( .a(n_21459), .o(n_21515) );
ao12f80 g547841 ( .a(n_19685), .b(n_20088), .c(n_19684), .o(n_21459) );
in01f80 g547842 ( .a(n_22118), .o(n_22127) );
ao12f80 g547843 ( .a(n_20399), .b(n_20814), .c(n_20398), .o(n_22118) );
oa12f80 g547844 ( .a(n_20711), .b(n_20710), .c(n_21025), .o(n_22134) );
ao12f80 g547845 ( .a(n_21688), .b(n_21687), .c(n_21686), .o(n_22330) );
ao12f80 g547846 ( .a(n_20041), .b(n_20040), .c(n_20039), .o(n_20806) );
in01f80 g547847 ( .a(n_21128), .o(n_21468) );
ao12f80 g547848 ( .a(n_19680), .b(n_20086), .c(n_19679), .o(n_21128) );
ao22s80 g547849 ( .a(n_21632), .b(n_21779), .c(n_21631), .d(n_20984), .o(n_22329) );
oa12f80 g547850 ( .a(n_21027), .b(n_21026), .c(n_21343), .o(n_22422) );
in01f80 g547851 ( .a(n_21478), .o(n_21824) );
ao12f80 g547852 ( .a(n_20077), .b(n_20450), .c(n_20076), .o(n_21478) );
ao12f80 g547853 ( .a(n_21685), .b(n_21684), .c(n_21683), .o(n_22328) );
ao22s80 g547854 ( .a(n_21306), .b(n_22623), .c(n_21305), .d(n_22012), .o(n_22624) );
in01f80 g547855 ( .a(n_21818), .o(n_21880) );
ao12f80 g547856 ( .a(n_20070), .b(n_20448), .c(n_20069), .o(n_21818) );
oa12f80 g547857 ( .a(n_20369), .b(n_20368), .c(n_20709), .o(n_21861) );
in01f80 g547858 ( .a(n_21900), .o(n_21474) );
oa12f80 g547859 ( .a(n_19689), .b(n_20090), .c(n_19688), .o(n_21900) );
ao12f80 g547860 ( .a(n_21738), .b(n_21737), .c(n_21736), .o(n_22327) );
ao12f80 g547861 ( .a(n_21366), .b(n_21365), .c(n_21364), .o(n_22075) );
oa12f80 g547862 ( .a(n_20407), .b(n_20406), .c(n_20405), .o(n_21860) );
in01f80 g547863 ( .a(n_20832), .o(n_20444) );
oa12f80 g547864 ( .a(n_19393), .b(n_19719), .c(n_19392), .o(n_20832) );
ao12f80 g547865 ( .a(n_21363), .b(n_21362), .c(n_21361), .o(n_22074) );
in01f80 g547866 ( .a(n_22393), .o(n_22696) );
ao22s80 g547867 ( .a(n_20983), .b(n_12546), .c(n_21776), .d(n_12545), .o(n_22393) );
oa12f80 g547868 ( .a(n_21020), .b(n_21021), .c(n_21019), .o(n_22415) );
in01f80 g547869 ( .a(n_21133), .o(n_21514) );
ao12f80 g547870 ( .a(n_19693), .b(n_20092), .c(n_19692), .o(n_21133) );
ao12f80 g547871 ( .a(n_20367), .b(n_20366), .c(n_20365), .o(n_21087) );
in01f80 g547872 ( .a(n_21126), .o(n_20805) );
oa12f80 g547873 ( .a(n_19683), .b(n_20087), .c(n_19682), .o(n_21126) );
ao12f80 g547874 ( .a(n_21682), .b(n_21681), .c(n_21680), .o(n_22326) );
ao22s80 g547875 ( .a(n_21302), .b(n_22324), .c(n_21301), .d(n_21621), .o(n_22325) );
in01f80 g547876 ( .a(n_22388), .o(n_22412) );
ao12f80 g547877 ( .a(n_20743), .b(n_21094), .c(n_20742), .o(n_22388) );
ao12f80 g547878 ( .a(n_21679), .b(n_21678), .c(n_21677), .o(n_22323) );
ao22s80 g547879 ( .a(n_21627), .b(n_22321), .c(n_21626), .d(n_21620), .o(n_22322) );
ao12f80 g547880 ( .a(n_20055), .b(n_20054), .c(n_20053), .o(n_20804) );
in01f80 g547881 ( .a(n_20443), .o(n_21541) );
oa12f80 g547882 ( .a(n_19391), .b(n_19718), .c(n_19390), .o(n_20443) );
in01f80 g547883 ( .a(n_21131), .o(n_21513) );
ao12f80 g547884 ( .a(n_19691), .b(n_20091), .c(n_19690), .o(n_21131) );
oa12f80 g547885 ( .a(n_20404), .b(n_20403), .c(n_20729), .o(n_21885) );
in01f80 g547886 ( .a(n_21544), .o(n_21122) );
oa12f80 g547887 ( .a(n_19395), .b(n_19720), .c(n_19394), .o(n_21544) );
in01f80 g547888 ( .a(n_21775), .o(n_22396) );
oa12f80 g547889 ( .a(n_20739), .b(n_21093), .c(n_20738), .o(n_21775) );
oa12f80 g547890 ( .a(n_21339), .b(n_21338), .c(n_21337), .o(n_22668) );
in01f80 g547891 ( .a(n_21489), .o(n_21834) );
ao12f80 g547892 ( .a(n_20072), .b(n_20447), .c(n_20071), .o(n_21489) );
ao12f80 g547893 ( .a(n_21673), .b(n_21672), .c(n_21671), .o(n_22320) );
ao12f80 g547894 ( .a(n_20419), .b(n_20801), .c(n_20418), .o(n_21086) );
in01f80 g547895 ( .a(n_21155), .o(n_21511) );
ao12f80 g547896 ( .a(n_19703), .b(n_20098), .c(n_19702), .o(n_21155) );
ao12f80 g547897 ( .a(n_22301), .b(n_22300), .c(n_22299), .o(n_22951) );
oa12f80 g547898 ( .a(n_21018), .b(n_21017), .c(n_21336), .o(n_22411) );
in01f80 g547899 ( .a(n_21123), .o(n_21509) );
ao12f80 g547900 ( .a(n_19687), .b(n_20089), .c(n_19686), .o(n_21123) );
ao12f80 g547901 ( .a(n_20416), .b(n_20795), .c(n_20415), .o(n_21085) );
ao12f80 g547902 ( .a(n_22039), .b(n_22038), .c(n_22037), .o(n_22622) );
oa12f80 g547903 ( .a(n_20036), .b(n_20035), .c(n_20037), .o(n_21503) );
ao12f80 g547904 ( .a(n_20362), .b(n_20361), .c(n_20360), .o(n_21084) );
ao22s80 g547905 ( .a(n_21635), .b(n_21622), .c(n_21636), .d(n_22318), .o(n_22319) );
ao12f80 g547906 ( .a(n_21668), .b(n_21667), .c(n_21666), .o(n_22317) );
oa12f80 g547907 ( .a(n_20728), .b(n_20727), .c(n_20726), .o(n_22731) );
ao12f80 g547908 ( .a(n_21665), .b(n_21664), .c(n_21663), .o(n_22316) );
ao12f80 g547909 ( .a(n_21662), .b(n_21661), .c(n_21660), .o(n_22315) );
in01f80 g547910 ( .a(n_21480), .o(n_21502) );
ao12f80 g547911 ( .a(n_19701), .b(n_20096), .c(n_19700), .o(n_21480) );
ao12f80 g547912 ( .a(n_20723), .b(n_21077), .c(n_20722), .o(n_21408) );
oa12f80 g547913 ( .a(n_21016), .b(n_21015), .c(n_21014), .o(n_22404) );
oa22f80 g547914 ( .a(n_20328), .b(FE_OFN264_n_4280), .c(n_1823), .d(n_28607), .o(n_21083) );
oa22f80 g547915 ( .a(n_22280), .b(FE_OFN219_n_23315), .c(n_1494), .d(n_28607), .o(n_22950) );
oa22f80 g547916 ( .a(n_21619), .b(FE_OFN221_n_23315), .c(n_1090), .d(FE_OFN128_n_27449), .o(n_22314) );
oa22f80 g547917 ( .a(n_21618), .b(FE_OFN206_n_28771), .c(n_288), .d(n_27452), .o(n_22313) );
oa22f80 g547918 ( .a(n_21295), .b(FE_OFN313_n_3069), .c(n_1287), .d(FE_OFN139_n_27449), .o(n_22073) );
oa22f80 g547919 ( .a(n_20975), .b(FE_OFN204_n_28771), .c(n_1079), .d(FE_OFN92_n_27449), .o(n_21774) );
oa22f80 g547920 ( .a(n_21617), .b(n_23315), .c(n_1657), .d(FE_OFN77_n_27012), .o(n_22312) );
oa22f80 g547921 ( .a(n_22011), .b(FE_OFN406_n_28303), .c(n_423), .d(FE_OFN76_n_27012), .o(n_22621) );
oa22f80 g547922 ( .a(n_20671), .b(FE_OFN256_n_4280), .c(n_529), .d(FE_OFN1174_n_4860), .o(n_21407) );
oa22f80 g547923 ( .a(n_21294), .b(FE_OFN417_n_28303), .c(n_1091), .d(n_27452), .o(n_22072) );
oa22f80 g547924 ( .a(n_20670), .b(FE_OFN310_n_3069), .c(n_1910), .d(FE_OFN20_n_27452), .o(n_21406) );
oa22f80 g547925 ( .a(n_21292), .b(FE_OFN308_n_3069), .c(n_1340), .d(n_27012), .o(n_22070) );
oa22f80 g547926 ( .a(n_21287), .b(FE_OFN309_n_3069), .c(n_1190), .d(n_27452), .o(n_22069) );
oa22f80 g547927 ( .a(n_20982), .b(FE_OFN299_n_3069), .c(n_1291), .d(FE_OFN21_n_27452), .o(n_21773) );
oa22f80 g547928 ( .a(n_20363), .b(FE_OFN314_n_3069), .c(n_1452), .d(FE_OFN17_n_29617), .o(n_20803) );
oa22f80 g547929 ( .a(n_20981), .b(FE_OFN308_n_3069), .c(n_1242), .d(n_29617), .o(n_21772) );
oa22f80 g547930 ( .a(n_21291), .b(n_28608), .c(n_731), .d(n_27452), .o(n_22068) );
oa22f80 g547931 ( .a(n_21616), .b(FE_OFN293_n_3069), .c(n_1379), .d(FE_OFN21_n_27452), .o(n_22311) );
oa22f80 g547932 ( .a(n_21290), .b(n_26454), .c(n_1566), .d(FE_OFN14_n_29068), .o(n_22067) );
oa22f80 g547933 ( .a(n_20980), .b(n_26454), .c(n_963), .d(FE_OFN14_n_29068), .o(n_21771) );
oa22f80 g547934 ( .a(n_22009), .b(n_28608), .c(n_111), .d(FE_OFN122_n_27449), .o(n_22620) );
oa22f80 g547935 ( .a(FE_OFN648_n_22008), .b(n_23813), .c(n_712), .d(FE_OFN105_n_27449), .o(n_22619) );
oa22f80 g547936 ( .a(n_22007), .b(FE_OFN162_n_26454), .c(n_94), .d(FE_OFN95_n_27449), .o(n_22618) );
oa22f80 g547937 ( .a(n_21293), .b(n_26454), .c(n_1338), .d(FE_OFN98_n_27449), .o(n_22066) );
oa22f80 g547938 ( .a(n_21289), .b(FE_OFN253_n_4280), .c(n_1257), .d(FE_OFN350_n_4860), .o(n_22065) );
oa22f80 g547939 ( .a(n_22002), .b(FE_OFN154_n_22615), .c(n_347), .d(FE_OFN17_n_29617), .o(n_22617) );
oa22f80 g547940 ( .a(n_22006), .b(n_22615), .c(n_1668), .d(FE_OFN98_n_27449), .o(n_22616) );
oa22f80 g547941 ( .a(n_22005), .b(FE_OFN235_n_4162), .c(n_77), .d(FE_OFN129_n_27449), .o(n_22614) );
oa22f80 g547942 ( .a(n_21999), .b(FE_OFN293_n_3069), .c(n_1000), .d(FE_OFN324_n_4860), .o(n_22613) );
oa22f80 g547943 ( .a(n_20038), .b(n_4162), .c(n_571), .d(FE_OFN353_n_4860), .o(n_20442) );
oa22f80 g547944 ( .a(n_21281), .b(n_4162), .c(n_91), .d(FE_OFN115_n_27449), .o(n_22064) );
oa22f80 g547945 ( .a(n_20801), .b(FE_OFN234_n_4162), .c(n_1523), .d(FE_OFN99_n_27449), .o(n_20802) );
oa22f80 g547946 ( .a(n_22004), .b(n_22960), .c(n_1688), .d(FE_OFN324_n_4860), .o(n_22612) );
oa22f80 g547947 ( .a(n_21286), .b(FE_OFN236_n_4162), .c(n_1500), .d(FE_OFN72_n_27012), .o(n_22063) );
oa22f80 g547948 ( .a(n_20034), .b(FE_OFN239_n_4162), .c(n_1179), .d(FE_OFN135_n_27449), .o(n_20441) );
oa22f80 g547949 ( .a(n_21285), .b(FE_OFN251_n_4162), .c(n_193), .d(rst), .o(n_22062) );
oa22f80 g547950 ( .a(n_20979), .b(FE_OFN295_n_3069), .c(n_384), .d(FE_OFN130_n_27449), .o(n_21770) );
oa22f80 g547951 ( .a(n_21768), .b(FE_OFN244_n_4162), .c(n_1748), .d(FE_OFN139_n_27449), .o(n_21769) );
oa22f80 g547952 ( .a(n_22003), .b(FE_OFN313_n_3069), .c(n_513), .d(FE_OFN1124_rst), .o(n_22611) );
oa22f80 g547953 ( .a(n_20977), .b(FE_OFN299_n_3069), .c(n_912), .d(FE_OFN1119_rst), .o(n_21767) );
oa22f80 g547954 ( .a(n_21284), .b(FE_OFN266_n_4280), .c(n_1294), .d(FE_OFN129_n_27449), .o(n_22061) );
oa22f80 g547955 ( .a(n_21283), .b(FE_OFN405_n_28303), .c(n_1040), .d(FE_OFN89_n_27449), .o(n_22060) );
oa22f80 g547956 ( .a(n_21081), .b(FE_OFN416_n_28303), .c(n_1847), .d(FE_OFN134_n_27449), .o(n_21082) );
oa22f80 g547957 ( .a(n_20976), .b(FE_OFN152_n_22615), .c(n_766), .d(FE_OFN361_n_4860), .o(n_21766) );
oa22f80 g547958 ( .a(n_21288), .b(FE_OFN152_n_22615), .c(n_1641), .d(FE_OFN349_n_4860), .o(n_22059) );
oa22f80 g547959 ( .a(n_19656), .b(FE_OFN240_n_4162), .c(n_1085), .d(FE_OFN142_n_27449), .o(n_20440) );
oa22f80 g547960 ( .a(n_22001), .b(FE_OFN152_n_22615), .c(n_811), .d(FE_OFN358_n_4860), .o(n_22610) );
oa22f80 g547961 ( .a(n_21615), .b(FE_OFN152_n_22615), .c(n_1507), .d(FE_OFN74_n_27012), .o(n_22309) );
oa22f80 g547962 ( .a(FE_OFN524_n_21282), .b(n_23291), .c(n_1750), .d(n_27449), .o(n_22058) );
oa22f80 g547963 ( .a(n_20326), .b(FE_OFN169_n_22948), .c(n_1406), .d(FE_OFN352_n_4860), .o(n_21080) );
oa22f80 g547964 ( .a(n_20325), .b(FE_OFN170_n_22948), .c(n_1697), .d(FE_OFN353_n_4860), .o(n_21079) );
oa22f80 g547965 ( .a(n_21279), .b(n_22615), .c(n_896), .d(FE_OFN335_n_4860), .o(n_22057) );
oa22f80 g547966 ( .a(n_21614), .b(FE_OFN406_n_28303), .c(n_945), .d(FE_OFN360_n_4860), .o(n_22308) );
oa22f80 g547967 ( .a(n_21278), .b(n_22615), .c(n_1590), .d(FE_OFN330_n_4860), .o(n_22056) );
oa22f80 g547968 ( .a(n_19678), .b(FE_OFN152_n_22615), .c(n_406), .d(FE_OFN104_n_27449), .o(n_20085) );
oa22f80 g547969 ( .a(n_20974), .b(FE_OFN254_n_4280), .c(n_1056), .d(FE_OFN142_n_27449), .o(n_21765) );
oa22f80 g547970 ( .a(n_20000), .b(FE_OFN269_n_4280), .c(n_1080), .d(FE_OFN1143_n_27012), .o(n_20800) );
oa22f80 g547971 ( .a(n_21277), .b(FE_OFN310_n_3069), .c(n_1635), .d(FE_OFN115_n_27449), .o(n_22055) );
oa22f80 g547972 ( .a(n_19681), .b(FE_OFN267_n_4280), .c(n_750), .d(FE_OFN92_n_27449), .o(n_20084) );
oa22f80 g547973 ( .a(n_21275), .b(FE_OFN299_n_3069), .c(n_1148), .d(FE_OFN350_n_4860), .o(n_22054) );
oa22f80 g547974 ( .a(n_20001), .b(FE_OFN297_n_3069), .c(n_1028), .d(FE_OFN138_n_27449), .o(n_20799) );
oa22f80 g547975 ( .a(n_21274), .b(FE_OFN296_n_3069), .c(n_1798), .d(FE_OFN11_n_29204), .o(n_22053) );
oa22f80 g547976 ( .a(n_19999), .b(FE_OFN300_n_3069), .c(n_1228), .d(FE_OFN326_n_4860), .o(n_20798) );
oa22f80 g547977 ( .a(n_21077), .b(n_21076), .c(n_1339), .d(n_27709), .o(n_21078) );
oa22f80 g547978 ( .a(n_21272), .b(FE_OFN269_n_4280), .c(n_1207), .d(n_29068), .o(n_22052) );
oa22f80 g547979 ( .a(FE_OFN771_n_20323), .b(n_21076), .c(n_1274), .d(n_27449), .o(n_21075) );
oa22f80 g547980 ( .a(n_22279), .b(FE_OFN171_n_22948), .c(n_1361), .d(FE_OFN1109_rst), .o(n_22949) );
oa22f80 g547981 ( .a(n_20322), .b(FE_OFN173_n_22948), .c(n_1390), .d(FE_OFN1123_rst), .o(n_21074) );
oa22f80 g547982 ( .a(n_22590), .b(FE_OFN311_n_3069), .c(n_850), .d(FE_OFN1174_n_4860), .o(n_23246) );
oa22f80 g547983 ( .a(n_19998), .b(FE_OFN169_n_22948), .c(n_854), .d(FE_OFN1120_rst), .o(n_20797) );
oa22f80 g547984 ( .a(n_21612), .b(FE_OFN410_n_28303), .c(n_1001), .d(FE_OFN130_n_27449), .o(n_22307) );
oa22f80 g547985 ( .a(n_21271), .b(n_28303), .c(n_1658), .d(FE_OFN68_n_27012), .o(n_22051) );
oa22f80 g547986 ( .a(n_22000), .b(FE_OFN265_n_4280), .c(n_1670), .d(FE_OFN134_n_27449), .o(n_22609) );
oa22f80 g547987 ( .a(n_21270), .b(n_23291), .c(n_1675), .d(n_27449), .o(n_22050) );
oa22f80 g547988 ( .a(n_20667), .b(n_23291), .c(n_1674), .d(FE_OFN95_n_27449), .o(n_21405) );
oa22f80 g547989 ( .a(n_20795), .b(FE_OFN247_n_4162), .c(n_1718), .d(FE_OFN134_n_27449), .o(n_20796) );
no02f80 g548068 ( .a(n_20097), .b(n_19716), .o(n_19717) );
no02f80 g548069 ( .a(n_21763), .b(n_21762), .o(n_21764) );
in01f80 g548070 ( .a(n_20793), .o(n_20794) );
no02f80 g548071 ( .a(n_20421), .b(x_in_2_6), .o(n_20793) );
no02f80 g548072 ( .a(n_21760), .b(n_21759), .o(n_21761) );
na02f80 g548073 ( .a(n_20792), .b(x_in_34_6), .o(n_21808) );
in01f80 g548074 ( .a(n_21072), .o(n_21073) );
no02f80 g548075 ( .a(n_20792), .b(x_in_34_6), .o(n_21072) );
no02f80 g548076 ( .a(n_22047), .b(n_22046), .o(n_22048) );
no02f80 g548077 ( .a(n_21757), .b(n_21756), .o(n_21758) );
na02f80 g548078 ( .a(n_21404), .b(x_in_8_9), .o(n_22368) );
in01f80 g548079 ( .a(n_21754), .o(n_21755) );
no02f80 g548080 ( .a(n_21404), .b(x_in_8_9), .o(n_21754) );
na02f80 g548081 ( .a(n_20791), .b(x_in_18_6), .o(n_21798) );
in01f80 g548082 ( .a(n_21070), .o(n_21071) );
no02f80 g548083 ( .a(n_20791), .b(x_in_18_6), .o(n_21070) );
na02f80 g548084 ( .a(n_21392), .b(x_in_56_8), .o(n_22367) );
na02f80 g548085 ( .a(n_21388), .b(x_in_36_6), .o(n_22366) );
no02f80 g548086 ( .a(n_21081), .b(n_20789), .o(n_20790) );
no02f80 g548087 ( .a(n_21752), .b(n_21751), .o(n_21753) );
na02f80 g548088 ( .a(n_20788), .b(x_in_50_6), .o(n_21787) );
in01f80 g548089 ( .a(n_21068), .o(n_21069) );
no02f80 g548090 ( .a(n_20788), .b(x_in_50_6), .o(n_21068) );
no02f80 g548091 ( .a(n_21749), .b(n_21748), .o(n_21750) );
in01f80 g548092 ( .a(n_23585), .o(n_21067) );
no02f80 g548093 ( .a(n_20787), .b(x_in_6_6), .o(n_23585) );
in01f80 g548094 ( .a(n_21805), .o(n_21066) );
na02f80 g548095 ( .a(n_20787), .b(x_in_6_6), .o(n_21805) );
no02f80 g548096 ( .a(n_20452), .b(n_20082), .o(n_20083) );
no02f80 g548097 ( .a(n_21746), .b(n_21745), .o(n_21747) );
na02f80 g548098 ( .a(n_20439), .b(x_in_10_6), .o(n_21450) );
in01f80 g548099 ( .a(n_20785), .o(n_20786) );
no02f80 g548100 ( .a(n_20439), .b(x_in_10_6), .o(n_20785) );
na02f80 g548101 ( .a(n_20438), .b(x_in_42_6), .o(n_21449) );
in01f80 g548102 ( .a(n_20783), .o(n_20784) );
no02f80 g548103 ( .a(n_20438), .b(x_in_42_6), .o(n_20783) );
na02f80 g548104 ( .a(n_20453), .b(n_20080), .o(n_20081) );
na02f80 g548105 ( .a(n_20437), .b(x_in_26_6), .o(n_21448) );
in01f80 g548106 ( .a(n_20781), .o(n_20782) );
no02f80 g548107 ( .a(n_20437), .b(x_in_26_6), .o(n_20781) );
no02f80 g548108 ( .a(n_21743), .b(n_21742), .o(n_21744) );
no02f80 g548109 ( .a(n_21740), .b(n_21739), .o(n_21741) );
in01f80 g548110 ( .a(n_21064), .o(n_21065) );
no02f80 g548111 ( .a(n_20761), .b(x_in_58_6), .o(n_21064) );
no02f80 g548112 ( .a(n_20327), .b(n_20789), .o(n_21892) );
in01f80 g548113 ( .a(n_21062), .o(n_21063) );
no02f80 g548114 ( .a(n_20780), .b(x_in_6_5), .o(n_21062) );
na02f80 g548115 ( .a(n_20780), .b(x_in_6_5), .o(n_21802) );
no02f80 g548116 ( .a(n_21737), .b(n_21736), .o(n_21738) );
no02f80 g548117 ( .a(n_21402), .b(n_21401), .o(n_21403) );
in01f80 g548118 ( .a(n_21399), .o(n_21400) );
na02f80 g548119 ( .a(n_21061), .b(n_20697), .o(n_21399) );
in01f80 g548120 ( .a(n_21734), .o(n_21735) );
na02f80 g548121 ( .a(n_21398), .b(n_21003), .o(n_21734) );
na02f80 g548122 ( .a(n_20779), .b(x_in_22_6), .o(n_21807) );
in01f80 g548123 ( .a(n_21059), .o(n_21060) );
no02f80 g548124 ( .a(n_20779), .b(x_in_22_6), .o(n_21059) );
no02f80 g548125 ( .a(n_21732), .b(n_21731), .o(n_21733) );
na02f80 g548126 ( .a(n_20436), .b(x_in_2_7), .o(n_21435) );
in01f80 g548127 ( .a(n_20777), .o(n_20778) );
no02f80 g548128 ( .a(n_20436), .b(x_in_2_7), .o(n_20777) );
na02f80 g548129 ( .a(n_20776), .b(x_in_54_6), .o(n_21801) );
in01f80 g548130 ( .a(n_21057), .o(n_21058) );
no02f80 g548131 ( .a(n_20776), .b(x_in_54_6), .o(n_21057) );
in01f80 g548132 ( .a(n_21108), .o(n_20435) );
na02f80 g548133 ( .a(n_20075), .b(x_in_52_6), .o(n_21108) );
na02f80 g548134 ( .a(n_20451), .b(n_20078), .o(n_20079) );
na02f80 g548135 ( .a(n_20775), .b(x_in_22_7), .o(n_21795) );
in01f80 g548136 ( .a(n_21055), .o(n_21056) );
no02f80 g548137 ( .a(n_20775), .b(x_in_22_7), .o(n_21055) );
no02f80 g548138 ( .a(n_21396), .b(n_21395), .o(n_21397) );
no02f80 g548139 ( .a(n_21729), .b(n_21728), .o(n_21730) );
na02f80 g548140 ( .a(n_20774), .b(x_in_40_6), .o(n_21786) );
in01f80 g548141 ( .a(n_21053), .o(n_21054) );
no02f80 g548142 ( .a(n_20774), .b(x_in_40_6), .o(n_21053) );
na02f80 g548143 ( .a(n_20104), .b(n_19714), .o(n_19715) );
na02f80 g548144 ( .a(n_19720), .b(n_19394), .o(n_19395) );
no02f80 g548145 ( .a(n_21726), .b(n_21725), .o(n_21727) );
in01f80 g548146 ( .a(n_21794), .o(n_21052) );
na02f80 g548147 ( .a(n_20752), .b(x_in_14_6), .o(n_21794) );
no02f80 g548148 ( .a(n_21723), .b(n_21722), .o(n_21724) );
na02f80 g548149 ( .a(n_20758), .b(x_in_46_6), .o(n_21799) );
no02f80 g548150 ( .a(n_21720), .b(n_21719), .o(n_21721) );
no02f80 g548151 ( .a(n_21717), .b(n_21716), .o(n_21718) );
na02f80 g548152 ( .a(n_20434), .b(x_in_54_7), .o(n_21444) );
in01f80 g548153 ( .a(n_20772), .o(n_20773) );
no02f80 g548154 ( .a(n_20434), .b(x_in_54_7), .o(n_20772) );
na02f80 g548155 ( .a(n_20771), .b(x_in_62_6), .o(n_21797) );
in01f80 g548156 ( .a(n_21050), .o(n_21051) );
no02f80 g548157 ( .a(n_20771), .b(x_in_62_6), .o(n_21050) );
in01f80 g548158 ( .a(n_21393), .o(n_21394) );
na02f80 g548159 ( .a(n_21049), .b(n_20702), .o(n_21393) );
no02f80 g548160 ( .a(n_21714), .b(n_21713), .o(n_21715) );
in01f80 g548161 ( .a(n_21711), .o(n_21712) );
no02f80 g548162 ( .a(n_21392), .b(x_in_56_8), .o(n_21711) );
no02f80 g548163 ( .a(n_21390), .b(n_21389), .o(n_21391) );
no02f80 g548164 ( .a(n_21709), .b(n_21708), .o(n_21710) );
in01f80 g548165 ( .a(n_21706), .o(n_21707) );
no02f80 g548166 ( .a(n_21388), .b(x_in_36_6), .o(n_21706) );
na02f80 g548167 ( .a(n_20099), .b(n_19712), .o(n_19713) );
no02f80 g548168 ( .a(n_21704), .b(n_21703), .o(n_21705) );
na02f80 g548169 ( .a(n_20770), .b(x_in_34_7), .o(n_21793) );
in01f80 g548170 ( .a(n_21047), .o(n_21048) );
no02f80 g548171 ( .a(n_20770), .b(x_in_34_7), .o(n_21047) );
na02f80 g548172 ( .a(n_20103), .b(n_19710), .o(n_19711) );
na02f80 g548173 ( .a(n_20433), .b(x_in_46_7), .o(n_21443) );
in01f80 g548174 ( .a(n_20768), .o(n_20769) );
no02f80 g548175 ( .a(n_20433), .b(x_in_46_7), .o(n_20768) );
no02f80 g548176 ( .a(n_21701), .b(n_21700), .o(n_21702) );
no02f80 g548177 ( .a(n_20102), .b(n_19708), .o(n_19709) );
na02f80 g548178 ( .a(n_20432), .b(x_in_16_7), .o(n_21442) );
in01f80 g548179 ( .a(n_20766), .o(n_20767) );
no02f80 g548180 ( .a(n_20432), .b(x_in_16_7), .o(n_20766) );
no02f80 g548181 ( .a(n_21386), .b(n_21385), .o(n_21387) );
no02f80 g548182 ( .a(n_22305), .b(n_22304), .o(n_22306) );
no02f80 g548183 ( .a(n_21383), .b(n_21382), .o(n_21384) );
na02f80 g548184 ( .a(n_20101), .b(n_19706), .o(n_19707) );
na02f80 g548185 ( .a(n_20431), .b(x_in_30_7), .o(n_21441) );
in01f80 g548186 ( .a(n_20764), .o(n_20765) );
no02f80 g548187 ( .a(n_20431), .b(x_in_30_7), .o(n_20764) );
na02f80 g548188 ( .a(n_20430), .b(x_in_18_7), .o(n_21439) );
in01f80 g548189 ( .a(n_20762), .o(n_20763) );
no02f80 g548190 ( .a(n_20430), .b(x_in_18_7), .o(n_20762) );
na02f80 g548191 ( .a(n_20761), .b(x_in_58_6), .o(n_21804) );
no02f80 g548192 ( .a(n_21698), .b(n_21697), .o(n_21699) );
na02f80 g548193 ( .a(n_20100), .b(n_19704), .o(n_19705) );
na02f80 g548194 ( .a(n_20429), .b(x_in_62_7), .o(n_21440) );
in01f80 g548195 ( .a(n_20759), .o(n_20760) );
no02f80 g548196 ( .a(n_20429), .b(x_in_62_7), .o(n_20759) );
in01f80 g548197 ( .a(n_21045), .o(n_21046) );
no02f80 g548198 ( .a(n_20757), .b(x_in_30_6), .o(n_21045) );
in01f80 g548199 ( .a(n_21043), .o(n_21044) );
no02f80 g548200 ( .a(n_20758), .b(x_in_46_6), .o(n_21043) );
no02f80 g548201 ( .a(n_21695), .b(n_21694), .o(n_21696) );
no02f80 g548202 ( .a(n_21380), .b(n_21379), .o(n_21381) );
in01f80 g548203 ( .a(n_21692), .o(n_21693) );
no02f80 g548204 ( .a(n_21378), .b(x_in_32_5), .o(n_21692) );
na02f80 g548205 ( .a(n_21378), .b(x_in_32_5), .o(n_22365) );
na02f80 g548206 ( .a(n_20757), .b(x_in_30_6), .o(n_21800) );
no02f80 g548207 ( .a(n_21376), .b(n_21375), .o(n_21377) );
no02f80 g548208 ( .a(n_22044), .b(n_22043), .o(n_22045) );
na02f80 g548209 ( .a(n_21042), .b(x_in_16_6), .o(n_22099) );
in01f80 g548210 ( .a(n_21373), .o(n_21374) );
no02f80 g548211 ( .a(n_21042), .b(x_in_16_6), .o(n_21373) );
in01f80 g548212 ( .a(n_20755), .o(n_20756) );
na02f80 g548213 ( .a(n_20428), .b(n_20027), .o(n_20755) );
no02f80 g548214 ( .a(n_21690), .b(n_21689), .o(n_21691) );
na02f80 g548215 ( .a(n_20427), .b(x_in_50_7), .o(n_21436) );
in01f80 g548216 ( .a(n_20753), .o(n_20754) );
no02f80 g548217 ( .a(n_20427), .b(x_in_50_7), .o(n_20753) );
na02f80 g548218 ( .a(n_21041), .b(x_in_48_5), .o(n_22098) );
in01f80 g548219 ( .a(n_21371), .o(n_21372) );
no02f80 g548220 ( .a(n_21041), .b(x_in_48_5), .o(n_21371) );
no02f80 g548221 ( .a(n_21687), .b(n_21686), .o(n_21688) );
na02f80 g548222 ( .a(n_21040), .b(x_in_8_8), .o(n_22097) );
in01f80 g548223 ( .a(n_21369), .o(n_21370) );
no02f80 g548224 ( .a(n_21040), .b(x_in_8_8), .o(n_21369) );
na02f80 g548225 ( .a(n_21039), .b(n_10610), .o(n_21780) );
no02f80 g548226 ( .a(n_20450), .b(n_20076), .o(n_20077) );
no02f80 g548227 ( .a(n_21684), .b(n_21683), .o(n_21685) );
na02f80 g548228 ( .a(n_21038), .b(x_in_40_5), .o(n_22096) );
in01f80 g548229 ( .a(n_21367), .o(n_21368) );
no02f80 g548230 ( .a(n_21038), .b(x_in_40_5), .o(n_21367) );
in01f80 g548231 ( .a(n_23258), .o(n_21037) );
no02f80 g548232 ( .a(n_20752), .b(x_in_14_6), .o(n_23258) );
in01f80 g548233 ( .a(n_23255), .o(n_20751) );
no02f80 g548234 ( .a(n_20426), .b(x_in_32_6), .o(n_23255) );
in01f80 g548235 ( .a(n_21431), .o(n_20750) );
na02f80 g548236 ( .a(n_20426), .b(x_in_32_6), .o(n_21431) );
no02f80 g548237 ( .a(n_21681), .b(n_21680), .o(n_21682) );
no02f80 g548238 ( .a(n_21365), .b(n_21364), .o(n_21366) );
na02f80 g548239 ( .a(n_20425), .b(x_in_24_8), .o(n_21430) );
in01f80 g548240 ( .a(n_20748), .o(n_20749) );
no02f80 g548241 ( .a(n_20425), .b(x_in_24_8), .o(n_20748) );
na02f80 g548242 ( .a(n_19719), .b(n_19392), .o(n_19393) );
no02f80 g548243 ( .a(n_21362), .b(n_21361), .o(n_21363) );
in01f80 g548244 ( .a(n_22302), .o(n_22303) );
na02f80 g548245 ( .a(n_22042), .b(n_21630), .o(n_22302) );
in01f80 g548246 ( .a(n_20746), .o(n_20747) );
na02f80 g548247 ( .a(n_20424), .b(n_20021), .o(n_20746) );
na02f80 g548248 ( .a(n_21036), .b(x_in_56_7), .o(n_22095) );
in01f80 g548249 ( .a(n_21359), .o(n_21360) );
no02f80 g548250 ( .a(n_21036), .b(x_in_56_7), .o(n_21359) );
na02f80 g548251 ( .a(n_20423), .b(x_in_10_7), .o(n_21427) );
in01f80 g548252 ( .a(n_20744), .o(n_20745) );
no02f80 g548253 ( .a(n_20423), .b(x_in_10_7), .o(n_20744) );
in01f80 g548254 ( .a(n_23262), .o(n_20422) );
no02f80 g548255 ( .a(n_20075), .b(x_in_52_6), .o(n_23262) );
na02f80 g548256 ( .a(n_21035), .b(x_in_48_6), .o(n_22094) );
in01f80 g548257 ( .a(n_21357), .o(n_21358) );
no02f80 g548258 ( .a(n_21035), .b(x_in_48_6), .o(n_21357) );
no02f80 g548259 ( .a(n_21094), .b(n_20742), .o(n_20743) );
na02f80 g548260 ( .a(n_21356), .b(x_in_20_6), .o(n_22369) );
no02f80 g548261 ( .a(n_21678), .b(n_21677), .o(n_21679) );
in01f80 g548262 ( .a(n_21675), .o(n_21676) );
no02f80 g548263 ( .a(n_21356), .b(x_in_20_6), .o(n_21675) );
no02f80 g548264 ( .a(n_21354), .b(n_21353), .o(n_21355) );
na02f80 g548265 ( .a(n_20421), .b(x_in_2_6), .o(n_21451) );
na02f80 g548266 ( .a(n_20420), .b(x_in_42_7), .o(n_21426) );
in01f80 g548267 ( .a(n_20740), .o(n_20741) );
no02f80 g548268 ( .a(n_20420), .b(x_in_42_7), .o(n_20740) );
na02f80 g548269 ( .a(n_21093), .b(n_20738), .o(n_20739) );
na02f80 g548270 ( .a(n_21674), .b(x_in_36_5), .o(n_22635) );
in01f80 g548271 ( .a(n_22040), .o(n_22041) );
no02f80 g548272 ( .a(n_21674), .b(x_in_36_5), .o(n_22040) );
no02f80 g548273 ( .a(n_21672), .b(n_21671), .o(n_21673) );
no02f80 g548274 ( .a(n_20801), .b(n_20418), .o(n_20419) );
no02f80 g548275 ( .a(n_20098), .b(n_19702), .o(n_19703) );
no02f80 g548276 ( .a(n_20002), .b(n_20418), .o(n_21510) );
no02f80 g548277 ( .a(n_22300), .b(n_22299), .o(n_22301) );
in01f80 g548278 ( .a(n_21669), .o(n_21670) );
no02f80 g548279 ( .a(n_21352), .b(x_in_20_5), .o(n_21669) );
na02f80 g548280 ( .a(n_21352), .b(x_in_20_5), .o(n_22355) );
in01f80 g548281 ( .a(n_21033), .o(n_21034) );
na02f80 g548282 ( .a(n_20737), .b(n_20341), .o(n_21033) );
na02f80 g548283 ( .a(n_20417), .b(x_in_26_7), .o(n_21425) );
in01f80 g548284 ( .a(n_20735), .o(n_20736) );
no02f80 g548285 ( .a(n_20417), .b(x_in_26_7), .o(n_20735) );
no02f80 g548286 ( .a(n_20795), .b(n_20415), .o(n_20416) );
no02f80 g548287 ( .a(n_19997), .b(n_20415), .o(n_21506) );
no02f80 g548288 ( .a(n_22038), .b(n_22037), .o(n_22039) );
in01f80 g548289 ( .a(n_21350), .o(n_21351) );
no02f80 g548290 ( .a(n_21032), .b(x_in_52_5), .o(n_21350) );
na02f80 g548291 ( .a(n_21032), .b(x_in_52_5), .o(n_22090) );
no02f80 g548292 ( .a(n_22035), .b(n_22034), .o(n_22036) );
no02f80 g548293 ( .a(n_21667), .b(n_21666), .o(n_21668) );
in01f80 g548294 ( .a(n_23250), .o(n_21031) );
no02f80 g548295 ( .a(n_20734), .b(x_in_12_6), .o(n_23250) );
in01f80 g548296 ( .a(n_21784), .o(n_21030) );
na02f80 g548297 ( .a(n_20734), .b(x_in_12_6), .o(n_21784) );
no02f80 g548298 ( .a(n_21664), .b(n_21663), .o(n_21665) );
no02f80 g548299 ( .a(n_21661), .b(n_21660), .o(n_21662) );
in01f80 g548300 ( .a(n_21658), .o(n_21659) );
no02f80 g548301 ( .a(n_21349), .b(x_in_44_7), .o(n_21658) );
na02f80 g548302 ( .a(n_21349), .b(x_in_44_7), .o(n_22353) );
no02f80 g548303 ( .a(n_20096), .b(n_19700), .o(n_19701) );
na02f80 g548304 ( .a(n_20414), .b(x_in_58_7), .o(n_21445) );
in01f80 g548305 ( .a(n_20732), .o(n_20733) );
no02f80 g548306 ( .a(n_20414), .b(x_in_58_7), .o(n_20732) );
in01f80 g548307 ( .a(n_21656), .o(n_21657) );
na02f80 g548308 ( .a(n_21348), .b(n_20992), .o(n_21656) );
na02f80 g548309 ( .a(n_21029), .b(x_in_60_6), .o(n_22100) );
in01f80 g548310 ( .a(n_21346), .o(n_21347) );
no02f80 g548311 ( .a(n_21029), .b(x_in_60_6), .o(n_21346) );
in01f80 g548312 ( .a(n_21344), .o(n_21345) );
no02f80 g548313 ( .a(n_21028), .b(x_in_60_5), .o(n_21344) );
na02f80 g548314 ( .a(n_21028), .b(x_in_60_5), .o(n_22091) );
na02f80 g548315 ( .a(n_20449), .b(n_20073), .o(n_20074) );
no02f80 g548316 ( .a(n_20095), .b(n_19698), .o(n_19699) );
no02f80 g548317 ( .a(n_20815), .b(n_20412), .o(n_20413) );
no02f80 g548318 ( .a(n_20447), .b(n_20071), .o(n_20072) );
no02f80 g548319 ( .a(n_20448), .b(n_20069), .o(n_20070) );
na02f80 g548320 ( .a(n_20094), .b(n_19696), .o(n_19697) );
no02f80 g548321 ( .a(n_21092), .b(n_20730), .o(n_20731) );
no02f80 g548322 ( .a(n_20093), .b(n_19694), .o(n_19695) );
no02f80 g548323 ( .a(n_20446), .b(n_20067), .o(n_20068) );
na02f80 g548324 ( .a(n_19718), .b(n_19390), .o(n_19391) );
no02f80 g548325 ( .a(n_20429), .b(n_20411), .o(n_21496) );
no02f80 g548326 ( .a(n_20775), .b(n_20729), .o(n_21838) );
no02f80 g548327 ( .a(n_20434), .b(n_20410), .o(n_21499) );
na02f80 g548328 ( .a(n_20065), .b(n_20410), .o(n_20066) );
no02f80 g548329 ( .a(n_20058), .b(n_20400), .o(n_21498) );
no02f80 g548330 ( .a(n_20433), .b(n_20409), .o(n_21497) );
no02f80 g548331 ( .a(n_20431), .b(n_20408), .o(n_21495) );
na02f80 g548332 ( .a(n_20063), .b(n_20408), .o(n_20064) );
na02f80 g548333 ( .a(n_20061), .b(n_20411), .o(n_20062) );
na02f80 g548334 ( .a(n_20059), .b(n_20409), .o(n_20060) );
na02f80 g548335 ( .a(n_21026), .b(n_21343), .o(n_21027) );
no02f80 g548336 ( .a(n_21404), .b(n_21343), .o(n_22654) );
na02f80 g548337 ( .a(n_20406), .b(n_20405), .o(n_20407) );
na02f80 g548338 ( .a(n_20406), .b(n_19894), .o(n_21781) );
na02f80 g548339 ( .a(n_20403), .b(n_20729), .o(n_20404) );
na02f80 g548340 ( .a(n_20401), .b(n_20400), .o(n_20402) );
no02f80 g548341 ( .a(n_20395), .b(n_20726), .o(n_21837) );
na02f80 g548342 ( .a(n_20727), .b(n_20726), .o(n_20728) );
no02f80 g548343 ( .a(n_20814), .b(n_20398), .o(n_20399) );
no02f80 g548344 ( .a(n_20092), .b(n_19692), .o(n_19693) );
no02f80 g548345 ( .a(n_20091), .b(n_19690), .o(n_19691) );
no02f80 g548346 ( .a(n_21768), .b(n_21341), .o(n_21342) );
no02f80 g548347 ( .a(n_20978), .b(n_21341), .o(n_22397) );
in01f80 g548348 ( .a(n_20396), .o(n_20397) );
na02f80 g548349 ( .a(n_20058), .b(x_in_14_7), .o(n_20396) );
na02f80 g548350 ( .a(n_20401), .b(n_1848), .o(n_21098) );
in01f80 g548351 ( .a(n_20724), .o(n_20725) );
na02f80 g548352 ( .a(n_20395), .b(x_in_12_7), .o(n_20724) );
na02f80 g548353 ( .a(n_20727), .b(n_1863), .o(n_21417) );
no02f80 g548354 ( .a(n_20445), .b(n_20056), .o(n_20057) );
na02f80 g548355 ( .a(n_20090), .b(n_19688), .o(n_19689) );
no02f80 g548356 ( .a(n_20089), .b(n_19686), .o(n_19687) );
no02f80 g548357 ( .a(n_20088), .b(n_19684), .o(n_19685) );
no02f80 g548358 ( .a(n_21077), .b(n_20722), .o(n_20723) );
no02f80 g548359 ( .a(n_20324), .b(n_20722), .o(n_21833) );
na02f80 g548360 ( .a(n_20087), .b(n_19682), .o(n_19683) );
no02f80 g548361 ( .a(n_20054), .b(n_20053), .o(n_20055) );
na02f80 g548362 ( .a(n_19681), .b(n_20053), .o(n_21137) );
no02f80 g548363 ( .a(n_20086), .b(n_19679), .o(n_19680) );
no02f80 g548364 ( .a(n_20720), .b(n_20719), .o(n_20721) );
na02f80 g548365 ( .a(n_20372), .b(n_19924), .o(n_21485) );
na02f80 g548366 ( .a(n_20717), .b(n_20250), .o(n_21831) );
na02f80 g548367 ( .a(n_20717), .b(n_20716), .o(n_20718) );
in01f80 g548368 ( .a(n_20715), .o(n_21462) );
no02f80 g548369 ( .a(n_20430), .b(n_20394), .o(n_20715) );
na02f80 g548370 ( .a(n_20051), .b(n_20394), .o(n_20052) );
in01f80 g548371 ( .a(n_20714), .o(n_21458) );
no02f80 g548372 ( .a(n_20427), .b(n_20393), .o(n_20714) );
no02f80 g548373 ( .a(n_20392), .b(n_19919), .o(n_21823) );
na02f80 g548374 ( .a(n_20375), .b(n_19922), .o(n_21483) );
na02f80 g548375 ( .a(n_20390), .b(n_20389), .o(n_20391) );
na02f80 g548376 ( .a(n_20387), .b(n_19920), .o(n_21482) );
na02f80 g548377 ( .a(n_20387), .b(n_20386), .o(n_20388) );
na02f80 g548378 ( .a(n_20384), .b(n_20708), .o(n_20385) );
no02f80 g548379 ( .a(n_20392), .b(n_20382), .o(n_20383) );
ao12f80 g548380 ( .a(n_10827), .b(n_20050), .c(n_12061), .o(n_21116) );
na02f80 g548381 ( .a(n_20048), .b(n_20378), .o(n_20049) );
no02f80 g548382 ( .a(n_20426), .b(n_20381), .o(n_21473) );
na02f80 g548383 ( .a(n_20379), .b(n_20381), .o(n_20380) );
in01f80 g548384 ( .a(n_20713), .o(n_21479) );
no02f80 g548385 ( .a(n_20414), .b(n_20378), .o(n_20713) );
no02f80 g548386 ( .a(n_20046), .b(n_20045), .o(n_20047) );
in01f80 g548387 ( .a(n_20044), .o(n_20831) );
na02f80 g548388 ( .a(n_19678), .b(n_20045), .o(n_20044) );
in01f80 g548389 ( .a(n_20712), .o(n_21470) );
no02f80 g548390 ( .a(n_20432), .b(n_20377), .o(n_20712) );
na02f80 g548391 ( .a(n_20042), .b(n_20377), .o(n_20043) );
in01f80 g548392 ( .a(n_21340), .o(n_22117) );
no02f80 g548393 ( .a(n_21035), .b(n_21025), .o(n_21340) );
na02f80 g548394 ( .a(n_20710), .b(n_21025), .o(n_20711) );
no02f80 g548395 ( .a(n_20040), .b(n_20039), .o(n_20041) );
no02f80 g548396 ( .a(n_20040), .b(n_19569), .o(n_21467) );
na02f80 g548397 ( .a(n_20375), .b(n_20374), .o(n_20376) );
na02f80 g548398 ( .a(n_20372), .b(n_20371), .o(n_20373) );
ao12f80 g548399 ( .a(n_9423), .b(n_20370), .c(n_9422), .o(n_21465) );
in01f80 g548400 ( .a(n_21024), .o(n_21817) );
no02f80 g548401 ( .a(n_20774), .b(n_20709), .o(n_21024) );
na02f80 g548402 ( .a(n_20368), .b(n_20709), .o(n_20369) );
ao22s80 g548403 ( .a(n_20237), .b(n_13012), .c(n_19937), .d(n_12891), .o(n_21791) );
oa12f80 g548404 ( .a(n_32734), .b(n_21022), .c(n_8896), .o(n_21023) );
na02f80 g548405 ( .a(n_21021), .b(n_20559), .o(n_22651) );
na02f80 g548406 ( .a(n_21021), .b(n_21019), .o(n_21020) );
no02f80 g548407 ( .a(n_20366), .b(n_20365), .o(n_20367) );
in01f80 g548408 ( .a(n_20364), .o(n_21125) );
na02f80 g548409 ( .a(n_20038), .b(n_20365), .o(n_20364) );
na02f80 g548410 ( .a(n_21338), .b(n_20922), .o(n_22390) );
na02f80 g548411 ( .a(n_21338), .b(n_21337), .o(n_21339) );
na02f80 g548412 ( .a(n_20390), .b(n_19921), .o(n_21484) );
in01f80 g548413 ( .a(n_21655), .o(n_22387) );
no02f80 g548414 ( .a(n_21356), .b(n_21336), .o(n_21655) );
na02f80 g548415 ( .a(n_21017), .b(n_21336), .o(n_21018) );
no02f80 g548416 ( .a(n_20787), .b(n_20708), .o(n_21821) );
in01f80 g548417 ( .a(n_20707), .o(n_21486) );
na02f80 g548418 ( .a(n_20363), .b(n_20719), .o(n_20707) );
no02f80 g548419 ( .a(n_20075), .b(n_20037), .o(n_21121) );
na02f80 g548420 ( .a(n_20035), .b(n_20037), .o(n_20036) );
no02f80 g548421 ( .a(n_20361), .b(n_20360), .o(n_20362) );
in01f80 g548422 ( .a(n_20359), .o(n_21118) );
na02f80 g548423 ( .a(n_20034), .b(n_20360), .o(n_20359) );
na02f80 g548424 ( .a(n_20032), .b(n_20393), .o(n_20033) );
na02f80 g548425 ( .a(n_21015), .b(n_20554), .o(n_22116) );
na02f80 g548426 ( .a(n_21015), .b(n_21014), .o(n_21016) );
in01f80 g548427 ( .a(n_23040), .o(n_22607) );
oa12f80 g548428 ( .a(n_21320), .b(n_20657), .c(n_21592), .o(n_23040) );
in01f80 g548429 ( .a(n_23037), .o(n_22947) );
oa12f80 g548430 ( .a(n_21303), .b(n_20655), .c(n_21591), .o(n_23037) );
in01f80 g548431 ( .a(n_22705), .o(n_23257) );
oa12f80 g548432 ( .a(n_21317), .b(n_20631), .c(n_21212), .o(n_22705) );
in01f80 g548433 ( .a(n_23034), .o(n_22946) );
oa12f80 g548434 ( .a(n_20700), .b(n_19987), .c(n_21590), .o(n_23034) );
in01f80 g548435 ( .a(n_23031), .o(n_22945) );
oa12f80 g548436 ( .a(n_20681), .b(n_19982), .c(n_21589), .o(n_23031) );
in01f80 g548437 ( .a(n_22985), .o(n_23584) );
oa12f80 g548438 ( .a(n_21004), .b(n_20311), .c(n_21587), .o(n_22985) );
in01f80 g548439 ( .a(n_22717), .o(n_22606) );
oa12f80 g548440 ( .a(n_20699), .b(n_21219), .c(n_19979), .o(n_22717) );
in01f80 g548441 ( .a(n_22665), .o(n_22605) );
oa12f80 g548442 ( .a(n_20698), .b(n_21213), .c(n_19977), .o(n_22665) );
in01f80 g548443 ( .a(n_22720), .o(n_22604) );
oa12f80 g548444 ( .a(n_21001), .b(n_20306), .c(n_21217), .o(n_22720) );
oa12f80 g548445 ( .a(n_12453), .b(n_20031), .c(n_13661), .o(n_20829) );
in01f80 g548446 ( .a(n_22298), .o(n_22971) );
oa12f80 g548447 ( .a(n_20165), .b(n_22028), .c(n_19427), .o(n_22298) );
in01f80 g548448 ( .a(n_22714), .o(n_22603) );
oa12f80 g548449 ( .a(n_21315), .b(n_20638), .c(n_21216), .o(n_22714) );
in01f80 g548450 ( .a(n_23013), .o(n_22944) );
oa12f80 g548451 ( .a(n_20692), .b(n_19971), .c(n_21586), .o(n_23013) );
in01f80 g548452 ( .a(n_22711), .o(n_22602) );
oa12f80 g548453 ( .a(n_21312), .b(n_20636), .c(n_21215), .o(n_22711) );
in01f80 g548454 ( .a(n_22693), .o(n_23263) );
oa12f80 g548455 ( .a(n_20347), .b(n_21214), .c(n_19643), .o(n_22693) );
in01f80 g548456 ( .a(n_23022), .o(n_22943) );
ao12f80 g548457 ( .a(n_19969), .b(n_20691), .c(n_21585), .o(n_23022) );
in01f80 g548458 ( .a(n_23025), .o(n_22942) );
oa12f80 g548459 ( .a(n_20993), .b(n_20263), .c(n_21584), .o(n_23025) );
in01f80 g548460 ( .a(n_22702), .o(n_22601) );
oa12f80 g548461 ( .a(n_21313), .b(n_20588), .c(n_21211), .o(n_22702) );
in01f80 g548462 ( .a(n_22699), .o(n_22600) );
oa12f80 g548463 ( .a(n_21314), .b(n_20626), .c(n_21210), .o(n_22699) );
in01f80 g548464 ( .a(n_22991), .o(n_22941) );
ao12f80 g548465 ( .a(n_19640), .b(n_20351), .c(n_21588), .o(n_22991) );
in01f80 g548466 ( .a(n_22687), .o(n_22599) );
oa12f80 g548467 ( .a(n_21304), .b(n_20624), .c(n_21209), .o(n_22687) );
in01f80 g548468 ( .a(n_22297), .o(n_22969) );
oa12f80 g548469 ( .a(n_19621), .b(n_22026), .c(n_19012), .o(n_22297) );
in01f80 g548470 ( .a(n_21654), .o(n_22383) );
oa12f80 g548471 ( .a(n_3230), .b(n_21333), .c(n_2179), .o(n_21654) );
in01f80 g548472 ( .a(n_23286), .o(n_23245) );
oa12f80 g548473 ( .a(n_21634), .b(n_20941), .c(n_21983), .o(n_23286) );
oa12f80 g548474 ( .a(n_20349), .b(n_19637), .c(n_21583), .o(n_23266) );
in01f80 g548475 ( .a(n_23605), .o(n_23579) );
oa12f80 g548476 ( .a(n_21000), .b(n_20293), .c(n_22275), .o(n_23605) );
in01f80 g548477 ( .a(n_23008), .o(n_22940) );
ao12f80 g548478 ( .a(n_19635), .b(n_20348), .c(n_21582), .o(n_23008) );
in01f80 g548479 ( .a(n_22690), .o(n_22598) );
ao12f80 g548480 ( .a(n_19966), .b(n_20690), .c(n_21207), .o(n_22690) );
in01f80 g548481 ( .a(n_22708), .o(n_22597) );
oa12f80 g548482 ( .a(n_20695), .b(n_21218), .c(n_19975), .o(n_22708) );
in01f80 g548483 ( .a(n_23005), .o(n_22939) );
oa12f80 g548484 ( .a(n_20346), .b(n_19632), .c(n_21581), .o(n_23005) );
in01f80 g548485 ( .a(n_22684), .o(n_22596) );
oa12f80 g548486 ( .a(n_20689), .b(n_19964), .c(n_21206), .o(n_22684) );
in01f80 g548487 ( .a(n_22595), .o(n_23260) );
oa12f80 g548488 ( .a(n_19265), .b(n_22290), .c(n_18567), .o(n_22595) );
oa12f80 g548489 ( .a(n_20685), .b(n_19962), .c(n_21580), .o(n_23265) );
in01f80 g548490 ( .a(n_23002), .o(n_22938) );
oa12f80 g548491 ( .a(n_20345), .b(n_19628), .c(n_21579), .o(n_23002) );
in01f80 g548492 ( .a(n_22033), .o(n_22647) );
oa12f80 g548493 ( .a(n_16548), .b(n_21650), .c(n_15903), .o(n_22033) );
in01f80 g548494 ( .a(n_22999), .o(n_22296) );
oa12f80 g548495 ( .a(n_21633), .b(n_20939), .c(n_20919), .o(n_22999) );
in01f80 g548496 ( .a(n_22681), .o(n_22295) );
oa12f80 g548497 ( .a(n_21310), .b(n_20604), .c(n_20918), .o(n_22681) );
in01f80 g548498 ( .a(n_22994), .o(n_22937) );
oa12f80 g548499 ( .a(n_20684), .b(n_19960), .c(n_21578), .o(n_22994) );
in01f80 g548500 ( .a(n_21653), .o(n_22381) );
oa12f80 g548501 ( .a(n_3268), .b(n_21330), .c(n_2177), .o(n_21653) );
in01f80 g548502 ( .a(n_22594), .o(n_23252) );
oa12f80 g548503 ( .a(n_20212), .b(n_22288), .c(n_19487), .o(n_22594) );
in01f80 g548504 ( .a(n_22676), .o(n_22032) );
oa12f80 g548505 ( .a(n_20995), .b(n_20271), .c(n_20551), .o(n_22676) );
in01f80 g548506 ( .a(n_22673), .o(n_23254) );
oa12f80 g548507 ( .a(n_20683), .b(n_19956), .c(n_21203), .o(n_22673) );
in01f80 g548508 ( .a(n_21652), .o(n_22378) );
oa12f80 g548509 ( .a(n_19623), .b(n_21327), .c(n_19008), .o(n_21652) );
oa12f80 g548510 ( .a(n_13126), .b(n_20358), .c(n_14272), .o(n_21117) );
in01f80 g548511 ( .a(n_22988), .o(n_22936) );
ao12f80 g548512 ( .a(n_19950), .b(n_21577), .c(n_20682), .o(n_22988) );
in01f80 g548513 ( .a(n_22294), .o(n_22967) );
oa12f80 g548514 ( .a(n_18922), .b(n_22024), .c(n_18305), .o(n_22294) );
in01f80 g548515 ( .a(n_23283), .o(n_23244) );
oa12f80 g548516 ( .a(n_21637), .b(n_20932), .c(n_21982), .o(n_23283) );
oa12f80 g548517 ( .a(n_16913), .b(n_21645), .c(n_16410), .o(n_22385) );
in01f80 g548518 ( .a(n_22723), .o(n_22593) );
oa12f80 g548519 ( .a(n_21299), .b(n_21205), .c(n_20600), .o(n_22723) );
in01f80 g548520 ( .a(n_22980), .o(n_22935) );
oa12f80 g548521 ( .a(n_20680), .b(n_21576), .c(n_19944), .o(n_22980) );
in01f80 g548522 ( .a(n_23278), .o(n_23243) );
oa12f80 g548523 ( .a(n_22013), .b(n_21232), .c(n_21981), .o(n_23278) );
in01f80 g548524 ( .a(n_23275), .o(n_23242) );
oa12f80 g548525 ( .a(n_21625), .b(n_20929), .c(n_21980), .o(n_23275) );
in01f80 g548526 ( .a(n_22977), .o(n_22934) );
oa12f80 g548527 ( .a(n_20679), .b(n_21575), .c(n_19940), .o(n_22977) );
in01f80 g548528 ( .a(n_22660), .o(n_22031) );
oa12f80 g548529 ( .a(n_21298), .b(n_20549), .c(n_20573), .o(n_22660) );
in01f80 g548530 ( .a(n_22657), .o(n_23249) );
oa12f80 g548531 ( .a(n_21297), .b(n_20571), .c(n_21202), .o(n_22657) );
in01f80 g548532 ( .a(n_22293), .o(n_22964) );
oa12f80 g548533 ( .a(n_20924), .b(n_22030), .c(n_20205), .o(n_22293) );
in01f80 g548534 ( .a(n_22292), .o(n_22962) );
oa12f80 g548535 ( .a(n_20175), .b(n_22022), .c(n_19417), .o(n_22292) );
in01f80 g548536 ( .a(n_22726), .o(n_22592) );
oa12f80 g548537 ( .a(n_20693), .b(n_21201), .c(n_19938), .o(n_22726) );
in01f80 g548538 ( .a(n_23028), .o(n_22933) );
oa12f80 g548539 ( .a(n_21316), .b(n_20566), .c(n_21574), .o(n_23028) );
in01f80 g548540 ( .a(n_23043), .o(n_22932) );
oa12f80 g548541 ( .a(n_21309), .b(n_20564), .c(n_21573), .o(n_23043) );
oa12f80 g548542 ( .a(n_11536), .b(n_20357), .c(n_12500), .o(n_21130) );
oa12f80 g548543 ( .a(n_9873), .b(n_19677), .c(n_11175), .o(n_20465) );
in01f80 g548544 ( .a(n_19064), .o(n_19725) );
ao12f80 g548545 ( .a(n_9530), .b(n_18683), .c(n_10814), .o(n_19064) );
oa12f80 g548546 ( .a(n_4383), .b(n_20030), .c(n_6651), .o(n_20827) );
oa12f80 g548547 ( .a(n_11812), .b(n_20029), .c(n_13120), .o(n_20828) );
ao12f80 g548548 ( .a(n_20676), .b(n_21009), .c(n_20675), .o(n_21335) );
in01f80 g548549 ( .a(n_20456), .o(n_20356) );
oa12f80 g548550 ( .a(n_19387), .b(n_19677), .c(n_19386), .o(n_20456) );
in01f80 g548551 ( .a(n_20826), .o(n_20706) );
oa12f80 g548552 ( .a(n_19674), .b(n_20031), .c(n_19673), .o(n_20826) );
ao12f80 g548553 ( .a(n_20007), .b(n_20006), .c(n_20005), .o(n_20705) );
oa12f80 g548554 ( .a(n_20010), .b(n_20009), .c(n_20338), .o(n_21110) );
ao22s80 g548555 ( .a(n_21208), .b(n_19503), .c(n_22290), .d(n_19504), .o(n_22291) );
ao22s80 g548556 ( .a(n_22028), .b(n_20490), .c(n_20920), .d(n_20489), .o(n_22029) );
oa22f80 g548557 ( .a(n_20354), .b(FE_OFN249_n_4162), .c(n_436), .d(FE_OFN92_n_27449), .o(n_20355) );
in01f80 g548558 ( .a(n_21099), .o(n_21421) );
ao12f80 g548559 ( .a(n_20025), .b(n_20357), .c(n_20024), .o(n_21099) );
ao22s80 g548560 ( .a(n_19948), .b(n_20921), .c(n_19949), .d(n_22026), .o(n_22027) );
ao22s80 g548561 ( .a(n_20241), .b(n_3708), .c(n_21333), .d(n_3709), .o(n_21334) );
in01f80 g548562 ( .a(n_21013), .o(n_21810) );
oa12f80 g548563 ( .a(n_20023), .b(n_20050), .c(n_20022), .o(n_21013) );
ao22s80 g548564 ( .a(n_21650), .b(n_16740), .c(n_20552), .d(n_16739), .o(n_21651) );
ao12f80 g548565 ( .a(n_20688), .b(n_20687), .c(n_20686), .o(n_21332) );
ao22s80 g548566 ( .a(n_21330), .b(n_4049), .c(n_20240), .d(n_4048), .o(n_21331) );
in01f80 g548567 ( .a(n_19396), .o(n_19722) );
ao12f80 g548568 ( .a(n_18397), .b(n_18683), .c(n_18396), .o(n_19396) );
in01f80 g548569 ( .a(n_22373), .o(n_22362) );
ao12f80 g548570 ( .a(n_20990), .b(n_21022), .c(n_20989), .o(n_22373) );
ao12f80 g548571 ( .a(n_20999), .b(n_20998), .c(n_20997), .o(n_21649) );
ao12f80 g548572 ( .a(n_20988), .b(n_20987), .c(n_20986), .o(n_21648) );
in01f80 g548573 ( .a(n_21329), .o(n_22109) );
oa12f80 g548574 ( .a(n_20343), .b(n_20370), .c(n_20342), .o(n_21329) );
ao12f80 g548575 ( .a(n_20013), .b(n_20354), .c(n_20012), .o(n_20704) );
ao12f80 g548577 ( .a(n_19670), .b(n_20030), .c(n_19669), .o(n_20821) );
oa12f80 g548578 ( .a(n_20015), .b(n_20016), .c(n_20014), .o(n_21105) );
in01f80 g548579 ( .a(n_21418), .o(n_21796) );
ao12f80 g548580 ( .a(n_20337), .b(n_20336), .c(n_20335), .o(n_21418) );
in01f80 g548581 ( .a(n_22400), .o(n_21647) );
oa12f80 g548582 ( .a(n_20674), .b(n_20673), .c(n_20672), .o(n_22400) );
ao12f80 g548583 ( .a(n_20334), .b(n_20333), .c(n_20332), .o(n_21012) );
in01f80 g548584 ( .a(n_21095), .o(n_21413) );
ao12f80 g548585 ( .a(n_20019), .b(n_20358), .c(n_20018), .o(n_21095) );
ao22s80 g548586 ( .a(n_22288), .b(n_20523), .c(n_21204), .d(n_20522), .o(n_22289) );
ao22s80 g548587 ( .a(n_19955), .b(n_21327), .c(n_19954), .d(n_20239), .o(n_21328) );
in01f80 g548588 ( .a(n_20817), .o(n_21104) );
ao12f80 g548589 ( .a(n_19668), .b(n_20029), .c(n_19667), .o(n_20817) );
ao22s80 g548590 ( .a(n_21645), .b(n_17178), .c(n_20550), .d(n_17177), .o(n_21646) );
ao22s80 g548591 ( .a(n_22024), .b(n_19205), .c(n_20916), .d(n_19204), .o(n_22025) );
ao12f80 g548592 ( .a(n_19063), .b(n_19388), .c(n_19062), .o(n_19676) );
in01f80 g548593 ( .a(n_22354), .o(n_22287) );
oa12f80 g548594 ( .a(n_21296), .b(n_21624), .c(n_21307), .o(n_22354) );
ao22s80 g548595 ( .a(n_22030), .b(n_21223), .c(n_20915), .d(n_21222), .o(n_22286) );
oa12f80 g548596 ( .a(n_20011), .b(n_20017), .c(n_20339), .o(n_21103) );
ao22s80 g548597 ( .a(n_22022), .b(n_20492), .c(n_20914), .d(n_20491), .o(n_22023) );
oa22f80 g548598 ( .a(n_20236), .b(FE_OFN411_n_28303), .c(n_437), .d(FE_OFN129_n_27449), .o(n_21326) );
oa22f80 g548599 ( .a(FE_OFN1031_n_19666), .b(n_22019), .c(n_1762), .d(n_29104), .o(n_20028) );
oa22f80 g548600 ( .a(FE_OFN498_n_20677), .b(n_22019), .c(n_1302), .d(n_29266), .o(n_21011) );
oa22f80 g548601 ( .a(n_19319), .b(FE_OFN249_n_4162), .c(n_1767), .d(n_29261), .o(n_20353) );
oa22f80 g548602 ( .a(FE_OFN789_n_20913), .b(n_22019), .c(n_1538), .d(n_29264), .o(n_22021) );
oa22f80 g548603 ( .a(n_20911), .b(n_22019), .c(n_851), .d(n_27449), .o(n_22020) );
oa22f80 g548604 ( .a(n_21009), .b(FE_OFN303_n_3069), .c(n_1068), .d(n_27709), .o(n_21010) );
oa22f80 g548605 ( .a(n_19893), .b(FE_OFN264_n_4280), .c(n_490), .d(n_29261), .o(n_21008) );
oa22f80 g548606 ( .a(n_20546), .b(FE_OFN314_n_3069), .c(n_1369), .d(FE_OFN330_n_4860), .o(n_21644) );
oa22f80 g548607 ( .a(n_20344), .b(FE_OFN240_n_4162), .c(n_1703), .d(FE_OFN138_n_27449), .o(n_20703) );
oa22f80 g548608 ( .a(n_20235), .b(FE_OFN259_n_4280), .c(n_1484), .d(FE_OFN76_n_27012), .o(n_21325) );
oa22f80 g548609 ( .a(n_20233), .b(FE_OFN253_n_4280), .c(n_917), .d(FE_OFN1121_rst), .o(n_21324) );
oa22f80 g548610 ( .a(n_19388), .b(FE_OFN266_n_4280), .c(n_526), .d(n_29264), .o(n_19389) );
oa22f80 g548611 ( .a(n_20544), .b(FE_OFN225_n_21642), .c(n_624), .d(FE_OFN104_n_27449), .o(n_21643) );
oa22f80 g548612 ( .a(n_19896), .b(FE_OFN223_n_21642), .c(n_1404), .d(FE_OFN360_n_4860), .o(n_21007) );
oa22f80 g548613 ( .a(n_20543), .b(FE_OFN223_n_21642), .c(n_465), .d(FE_OFN76_n_27012), .o(n_21641) );
oa22f80 g548614 ( .a(n_19318), .b(FE_OFN223_n_21642), .c(n_110), .d(FE_OFN92_n_27449), .o(n_20352) );
oa22f80 g548615 ( .a(n_20232), .b(FE_OFN260_n_4280), .c(n_1411), .d(rst), .o(n_21323) );
oa22f80 g548616 ( .a(n_21623), .b(FE_OFN268_n_4280), .c(n_1423), .d(FE_OFN124_n_27449), .o(n_22018) );
oa22f80 g548617 ( .a(n_21200), .b(FE_OFN268_n_4280), .c(n_873), .d(FE_OFN124_n_27449), .o(n_22285) );
oa22f80 g548618 ( .a(n_20231), .b(FE_OFN223_n_21642), .c(n_845), .d(FE_OFN72_n_27012), .o(n_21322) );
oa22f80 g548619 ( .a(n_20542), .b(FE_OFN225_n_21642), .c(n_1424), .d(FE_OFN104_n_27449), .o(n_21640) );
oa22f80 g548620 ( .a(n_20230), .b(FE_OFN224_n_21642), .c(n_1004), .d(n_27449), .o(n_21321) );
oa22f80 g548621 ( .a(n_20541), .b(FE_OFN402_n_28303), .c(n_1434), .d(FE_OFN134_n_27449), .o(n_21639) );
oa22f80 g548622 ( .a(n_19898), .b(FE_OFN224_n_21642), .c(n_365), .d(n_29264), .o(n_21006) );
oa22f80 g548623 ( .a(n_18675), .b(FE_OFN224_n_21642), .c(n_1096), .d(FE_OFN335_n_4860), .o(n_19675) );
oa22f80 g548624 ( .a(n_21199), .b(FE_OFN223_n_21642), .c(n_1442), .d(FE_OFN65_n_27012), .o(n_22284) );
oa22f80 g548625 ( .a(n_20910), .b(FE_OFN402_n_28303), .c(n_133), .d(FE_OFN134_n_27449), .o(n_22017) );
in01f80 g548656 ( .a(n_20701), .o(n_20702) );
no02f80 g548657 ( .a(n_20405), .b(x_in_24_10), .o(n_20701) );
na02f80 g548658 ( .a(n_21320), .b(n_20658), .o(n_21760) );
na02f80 g548659 ( .a(n_21637), .b(n_20933), .o(n_22047) );
in01f80 g548660 ( .a(n_21318), .o(n_21319) );
na02f80 g548661 ( .a(n_21005), .b(n_20274), .o(n_21318) );
na02f80 g548662 ( .a(n_20700), .b(n_19988), .o(n_21752) );
na02f80 g548663 ( .a(n_21004), .b(n_20312), .o(n_21743) );
na02f80 g548664 ( .a(n_20699), .b(n_19980), .o(n_21396) );
na02f80 g548665 ( .a(n_21317), .b(n_20632), .o(n_21714) );
na02f80 g548666 ( .a(n_20698), .b(n_19978), .o(n_21354) );
na02f80 g548667 ( .a(n_20351), .b(n_19641), .o(n_21732) );
na02f80 g548668 ( .a(n_21316), .b(n_20567), .o(n_21681) );
na02f80 g548669 ( .a(n_20031), .b(n_19673), .o(n_19674) );
na02f80 g548670 ( .a(n_20350), .b(x_in_38_9), .o(n_21061) );
in01f80 g548671 ( .a(n_20696), .o(n_20697) );
no02f80 g548672 ( .a(n_20350), .b(x_in_38_9), .o(n_20696) );
na02f80 g548673 ( .a(n_20695), .b(n_19976), .o(n_21376) );
na02f80 g548674 ( .a(n_20694), .b(x_in_38_8), .o(n_21398) );
in01f80 g548675 ( .a(n_21002), .o(n_21003) );
no02f80 g548676 ( .a(n_20694), .b(x_in_38_8), .o(n_21002) );
in01f80 g548677 ( .a(n_20026), .o(n_20027) );
no02f80 g548678 ( .a(n_19672), .b(x_in_24_9), .o(n_20026) );
na02f80 g548679 ( .a(n_21315), .b(n_20639), .o(n_21749) );
na02f80 g548680 ( .a(n_21314), .b(n_20627), .o(n_21717) );
na02f80 g548681 ( .a(n_20693), .b(n_19939), .o(n_21390) );
na02f80 g548682 ( .a(n_21313), .b(n_20589), .o(n_21720) );
na02f80 g548683 ( .a(n_21312), .b(n_20637), .o(n_21729) );
na02f80 g548684 ( .a(n_21001), .b(n_20307), .o(n_21402) );
na02f80 g548685 ( .a(n_20405), .b(x_in_24_10), .o(n_21049) );
na02f80 g548686 ( .a(n_19672), .b(x_in_24_9), .o(n_20428) );
no02f80 g548687 ( .a(n_20357), .b(n_20024), .o(n_20025) );
na02f80 g548688 ( .a(n_20692), .b(n_19972), .o(n_21709) );
in01f80 g548689 ( .a(n_21635), .o(n_21636) );
na02f80 g548690 ( .a(n_21311), .b(n_20623), .o(n_21635) );
na02f80 g548691 ( .a(n_21634), .b(n_20942), .o(n_22035) );
na02f80 g548692 ( .a(n_20349), .b(n_19638), .o(n_21704) );
na02f80 g548693 ( .a(n_20691), .b(n_19970), .o(n_21723) );
na02f80 g548694 ( .a(n_20348), .b(n_19636), .o(n_21701) );
na02f80 g548695 ( .a(n_20347), .b(n_19644), .o(n_21386) );
na02f80 g548696 ( .a(n_21000), .b(n_20294), .o(n_22305) );
na02f80 g548697 ( .a(n_20050), .b(n_20022), .o(n_20023) );
na02f80 g548698 ( .a(n_20690), .b(n_19967), .o(n_21383) );
na02f80 g548699 ( .a(n_20346), .b(n_19633), .o(n_21698) );
no02f80 g548700 ( .a(n_18395), .b(n_19062), .o(n_19721) );
na02f80 g548701 ( .a(n_20345), .b(n_19629), .o(n_21695) );
na02f80 g548702 ( .a(n_20689), .b(n_19965), .o(n_21380) );
na02f80 g548703 ( .a(n_21633), .b(n_20940), .o(n_22044) );
no02f80 g548704 ( .a(n_20687), .b(n_20686), .o(n_20688) );
na02f80 g548705 ( .a(n_20344), .b(n_20686), .o(n_21437) );
na02f80 g548706 ( .a(n_21310), .b(n_20605), .o(n_21690) );
na02f80 g548707 ( .a(n_20685), .b(n_19963), .o(n_21687) );
na02f80 g548708 ( .a(n_21309), .b(n_20565), .o(n_21763) );
no02f80 g548709 ( .a(n_20998), .b(n_20997), .o(n_20999) );
in01f80 g548710 ( .a(n_21631), .o(n_21632) );
na02f80 g548711 ( .a(n_21308), .b(n_20603), .o(n_21631) );
na02f80 g548712 ( .a(n_21307), .b(x_in_44_8), .o(n_22042) );
in01f80 g548713 ( .a(n_21629), .o(n_21630) );
no02f80 g548714 ( .a(n_21307), .b(x_in_44_8), .o(n_21629) );
na02f80 g548715 ( .a(n_20684), .b(n_19961), .o(n_21684) );
na02f80 g548716 ( .a(n_20370), .b(n_20342), .o(n_20343) );
in01f80 g548717 ( .a(n_21305), .o(n_21306) );
na02f80 g548718 ( .a(n_20996), .b(n_20276), .o(n_21305) );
na02f80 g548719 ( .a(n_21304), .b(n_20625), .o(n_21737) );
na02f80 g548720 ( .a(n_20995), .b(n_20272), .o(n_21365) );
na02f80 g548721 ( .a(n_19671), .b(x_in_24_7), .o(n_20424) );
in01f80 g548722 ( .a(n_20020), .o(n_20021) );
no02f80 g548723 ( .a(n_19671), .b(x_in_24_7), .o(n_20020) );
in01f80 g548724 ( .a(n_22282), .o(n_22283) );
na02f80 g548725 ( .a(n_22016), .b(n_21228), .o(n_22282) );
na02f80 g548726 ( .a(n_21303), .b(n_20656), .o(n_21757) );
no02f80 g548727 ( .a(n_20358), .b(n_20018), .o(n_20019) );
na02f80 g548728 ( .a(n_20683), .b(n_19957), .o(n_21362) );
in01f80 g548729 ( .a(n_22014), .o(n_22015) );
na02f80 g548730 ( .a(n_21628), .b(n_20935), .o(n_22014) );
na02f80 g548731 ( .a(n_20017), .b(x_in_28_9), .o(n_20737) );
in01f80 g548732 ( .a(n_20340), .o(n_20341) );
no02f80 g548733 ( .a(n_20017), .b(x_in_28_9), .o(n_20340) );
in01f80 g548734 ( .a(n_21301), .o(n_21302) );
na02f80 g548735 ( .a(n_20994), .b(n_20266), .o(n_21301) );
na02f80 g548736 ( .a(n_20993), .b(n_20264), .o(n_21726) );
na02f80 g548737 ( .a(n_20682), .b(n_19951), .o(n_21678) );
in01f80 g548738 ( .a(n_21626), .o(n_21627) );
na02f80 g548739 ( .a(n_21300), .b(n_20586), .o(n_21626) );
na02f80 g548740 ( .a(n_20681), .b(n_19983), .o(n_21746) );
na02f80 g548741 ( .a(n_21299), .b(n_20601), .o(n_21740) );
na02f80 g548742 ( .a(n_20680), .b(n_19945), .o(n_21672) );
na02f80 g548743 ( .a(n_22013), .b(n_21233), .o(n_22300) );
na02f80 g548744 ( .a(n_21625), .b(n_20930), .o(n_22038) );
na02f80 g548745 ( .a(n_21298), .b(n_20574), .o(n_21667) );
na02f80 g548746 ( .a(n_20679), .b(n_19941), .o(n_21664) );
no02f80 g548747 ( .a(n_19388), .b(n_19062), .o(n_19063) );
na02f80 g548748 ( .a(n_21297), .b(n_20572), .o(n_21661) );
na02f80 g548749 ( .a(n_20678), .b(x_in_28_8), .o(n_21348) );
in01f80 g548750 ( .a(n_20991), .o(n_20992) );
no02f80 g548751 ( .a(n_20678), .b(x_in_28_8), .o(n_20991) );
no02f80 g548752 ( .a(n_21022), .b(n_20989), .o(n_20990) );
na02f80 g548753 ( .a(n_19677), .b(n_19386), .o(n_19387) );
no02f80 g548754 ( .a(n_18683), .b(n_18396), .o(n_18397) );
no02f80 g548755 ( .a(n_20987), .b(n_20986), .o(n_20988) );
na02f80 g548756 ( .a(FE_OFN498_n_20677), .b(n_20986), .o(n_21782) );
no02f80 g548757 ( .a(n_19320), .b(n_20012), .o(n_21100) );
no02f80 g548758 ( .a(n_21009), .b(n_20675), .o(n_20676) );
no02f80 g548759 ( .a(n_19899), .b(n_20675), .o(n_21420) );
no02f80 g548760 ( .a(n_20016), .b(n_19672), .o(n_20406) );
na02f80 g548761 ( .a(n_20016), .b(n_20014), .o(n_20015) );
no02f80 g548762 ( .a(n_20354), .b(n_20012), .o(n_20013) );
na02f80 g548763 ( .a(n_21624), .b(n_21307), .o(n_21296) );
na02f80 g548764 ( .a(n_21624), .b(n_21623), .o(n_22352) );
no02f80 g548765 ( .a(n_20246), .b(n_7109), .o(n_20985) );
na02f80 g548766 ( .a(n_19562), .b(n_20339), .o(n_21097) );
na02f80 g548767 ( .a(n_20017), .b(n_20339), .o(n_20011) );
no02f80 g548768 ( .a(n_20030), .b(n_19669), .o(n_19670) );
no02f80 g548769 ( .a(n_20029), .b(n_19667), .o(n_19668) );
na02f80 g548770 ( .a(n_20009), .b(n_20338), .o(n_20010) );
no02f80 g548771 ( .a(n_20350), .b(n_20338), .o(n_21096) );
in01f80 g548772 ( .a(n_20008), .o(n_20454) );
na02f80 g548773 ( .a(FE_OFN1031_n_19666), .b(n_20005), .o(n_20008) );
no02f80 g548774 ( .a(n_20006), .b(n_20005), .o(n_20007) );
no02f80 g548775 ( .a(n_20336), .b(n_20335), .o(n_20337) );
na02f80 g548776 ( .a(n_20673), .b(n_20672), .o(n_20674) );
oa12f80 g548777 ( .a(n_11512), .b(n_19061), .c(n_12492), .o(n_19719) );
no02f80 g548778 ( .a(n_20333), .b(n_20332), .o(n_20334) );
no02f80 g548779 ( .a(n_20333), .b(n_19524), .o(n_21412) );
in01f80 g548780 ( .a(n_22281), .o(n_22953) );
oa12f80 g548781 ( .a(n_19886), .b(n_22010), .c(n_19192), .o(n_22281) );
ao12f80 g548782 ( .a(n_15569), .b(n_19665), .c(n_16262), .o(n_20452) );
ao12f80 g548783 ( .a(n_13608), .b(n_19664), .c(n_14785), .o(n_20453) );
oa12f80 g548784 ( .a(n_15557), .b(n_19060), .c(n_16261), .o(n_19720) );
oa12f80 g548785 ( .a(n_14778), .b(n_19663), .c(n_15414), .o(n_20451) );
oa12f80 g548786 ( .a(n_14764), .b(n_19385), .c(n_15418), .o(n_20104) );
in01f80 g548787 ( .a(n_21622), .o(n_22318) );
ao12f80 g548788 ( .a(n_19272), .b(n_19869), .c(n_21280), .o(n_21622) );
oa12f80 g548789 ( .a(n_14752), .b(n_19384), .c(n_15407), .o(n_20099) );
oa12f80 g548790 ( .a(n_14741), .b(n_19383), .c(n_15397), .o(n_20103) );
ao12f80 g548791 ( .a(n_14380), .b(n_19382), .c(n_15142), .o(n_20102) );
oa12f80 g548792 ( .a(n_14713), .b(n_19381), .c(n_15385), .o(n_20101) );
oa12f80 g548793 ( .a(n_14687), .b(n_19380), .c(n_15367), .o(n_20100) );
in01f80 g548794 ( .a(n_20984), .o(n_21779) );
oa12f80 g548795 ( .a(n_20277), .b(n_19528), .c(n_19540), .o(n_20984) );
ao12f80 g548796 ( .a(n_13152), .b(n_19662), .c(n_14317), .o(n_20450) );
in01f80 g548797 ( .a(n_22012), .o(n_22623) );
oa12f80 g548798 ( .a(n_19881), .b(n_21613), .c(n_19225), .o(n_22012) );
ao12f80 g548799 ( .a(n_12304), .b(n_20669), .c(n_12954), .o(n_21039) );
oa12f80 g548800 ( .a(n_16100), .b(n_20331), .c(n_16680), .o(n_21094) );
in01f80 g548801 ( .a(n_20983), .o(n_21776) );
ao12f80 g548802 ( .a(n_11018), .b(n_20668), .c(n_12121), .o(n_20983) );
in01f80 g548803 ( .a(n_21621), .o(n_22324) );
oa12f80 g548804 ( .a(n_19535), .b(n_21276), .c(n_18932), .o(n_21621) );
in01f80 g548805 ( .a(n_21620), .o(n_22321) );
oa12f80 g548806 ( .a(n_19874), .b(n_21273), .c(n_19213), .o(n_21620) );
oa12f80 g548807 ( .a(n_15533), .b(n_20330), .c(n_16250), .o(n_21093) );
ao12f80 g548808 ( .a(n_12254), .b(n_19379), .c(n_12436), .o(n_20098) );
ao12f80 g548809 ( .a(n_11423), .b(n_19378), .c(n_12429), .o(n_20097) );
ao12f80 g548810 ( .a(n_14216), .b(n_19377), .c(n_15086), .o(n_20096) );
ao12f80 g548811 ( .a(n_14707), .b(n_19661), .c(n_15372), .o(n_20449) );
ao12f80 g548812 ( .a(n_14347), .b(n_19376), .c(n_15131), .o(n_20095) );
ao12f80 g548813 ( .a(n_16081), .b(n_20004), .c(n_16673), .o(n_20815) );
ao12f80 g548814 ( .a(n_14305), .b(n_19660), .c(n_15113), .o(n_20448) );
oa12f80 g548815 ( .a(n_8828), .b(n_19659), .c(n_9526), .o(n_20447) );
oa12f80 g548816 ( .a(n_13199), .b(n_19375), .c(n_14405), .o(n_20094) );
ao12f80 g548817 ( .a(n_13183), .b(n_20329), .c(n_14367), .o(n_21092) );
oa12f80 g548818 ( .a(n_14444), .b(n_19374), .c(n_15161), .o(n_20093) );
oa12f80 g548819 ( .a(n_14417), .b(n_19658), .c(n_15155), .o(n_20446) );
oa12f80 g548820 ( .a(n_11492), .b(n_19059), .c(n_11790), .o(n_19718) );
ao12f80 g548821 ( .a(n_13163), .b(n_20003), .c(n_14327), .o(n_20814) );
ao12f80 g548822 ( .a(n_14257), .b(n_19373), .c(n_15179), .o(n_20092) );
ao12f80 g548823 ( .a(n_13899), .b(n_19372), .c(n_14910), .o(n_20091) );
ao12f80 g548824 ( .a(n_11477), .b(n_19657), .c(n_12459), .o(n_20445) );
ao12f80 g548825 ( .a(n_15522), .b(n_19371), .c(n_16258), .o(n_20090) );
ao12f80 g548826 ( .a(n_13881), .b(n_19370), .c(n_14941), .o(n_20089) );
oa12f80 g548827 ( .a(n_13957), .b(n_19369), .c(n_14932), .o(n_20088) );
ao12f80 g548828 ( .a(n_10669), .b(n_19368), .c(n_11801), .o(n_20087) );
oa12f80 g548829 ( .a(n_8278), .b(n_19367), .c(n_9465), .o(n_20086) );
ao12f80 g548830 ( .a(n_19588), .b(FE_OFN1061_n_19587), .c(n_19586), .o(n_20328) );
ao12f80 g548831 ( .a(n_21598), .b(n_21597), .c(n_21596), .o(n_22280) );
oa12f80 g548832 ( .a(n_19338), .b(n_19337), .c(n_19585), .o(n_20421) );
ao12f80 g548833 ( .a(n_20955), .b(n_20954), .c(n_20953), .o(n_21619) );
oa12f80 g548834 ( .a(n_19574), .b(n_19573), .c(n_19923), .o(n_20792) );
ao12f80 g548835 ( .a(n_20952), .b(n_20951), .c(n_20950), .o(n_21618) );
ao12f80 g548836 ( .a(n_20563), .b(n_20562), .c(n_20561), .o(n_21295) );
ao12f80 g548837 ( .a(n_20949), .b(n_20948), .c(n_20947), .o(n_21617) );
ao22s80 g548838 ( .a(n_20216), .b(n_20905), .c(n_20217), .d(n_22010), .o(n_22011) );
oa12f80 g548839 ( .a(n_19565), .b(n_19564), .c(n_19563), .o(n_20791) );
ao12f80 g548840 ( .a(n_19986), .b(n_19985), .c(n_19984), .o(n_20671) );
ao12f80 g548841 ( .a(n_20651), .b(n_20650), .c(n_20649), .o(n_21294) );
oa12f80 g548842 ( .a(n_19584), .b(n_19583), .c(n_19582), .o(n_20788) );
ao12f80 g548843 ( .a(n_20635), .b(n_20634), .c(n_20633), .o(n_21293) );
in01f80 g548844 ( .a(n_20384), .o(n_20787) );
ao12f80 g548845 ( .a(n_19365), .b(n_19665), .c(n_19364), .o(n_20384) );
ao12f80 g548846 ( .a(n_19918), .b(FE_OFN918_n_19575), .c(n_19916), .o(n_20670) );
ao12f80 g548847 ( .a(n_20648), .b(n_20647), .c(n_20646), .o(n_21292) );
oa12f80 g548848 ( .a(n_19324), .b(n_19323), .c(n_19581), .o(n_20439) );
ao12f80 g548849 ( .a(n_20310), .b(n_20309), .c(n_20308), .o(n_20982) );
oa12f80 g548850 ( .a(n_19334), .b(n_19333), .c(n_19580), .o(n_20438) );
ao12f80 g548851 ( .a(n_20297), .b(n_20296), .c(n_20295), .o(n_20981) );
oa12f80 g548852 ( .a(n_19328), .b(n_19327), .c(n_19579), .o(n_20437) );
ao12f80 g548853 ( .a(n_20645), .b(n_20644), .c(n_20643), .o(n_21291) );
oa12f80 g548854 ( .a(n_19596), .b(n_19595), .c(n_19603), .o(n_20776) );
ao12f80 g548855 ( .a(n_20642), .b(n_20641), .c(n_20640), .o(n_21290) );
ao12f80 g548856 ( .a(n_20946), .b(n_20945), .c(n_20944), .o(n_21616) );
oa12f80 g548857 ( .a(n_19578), .b(n_19577), .c(n_19576), .o(n_20761) );
ao12f80 g548858 ( .a(n_20280), .b(n_20279), .c(n_20278), .o(n_20980) );
oa12f80 g548859 ( .a(n_19567), .b(n_19901), .c(n_19566), .o(n_20780) );
in01f80 g548860 ( .a(n_20065), .o(n_20434) );
ao12f80 g548861 ( .a(n_19058), .b(n_19385), .c(n_19057), .o(n_20065) );
ao12f80 g548862 ( .a(n_21248), .b(n_21247), .c(n_21246), .o(n_22009) );
in01f80 g548863 ( .a(n_20363), .o(n_20720) );
ao12f80 g548864 ( .a(n_19363), .b(n_19664), .c(n_19362), .o(n_20363) );
oa12f80 g548865 ( .a(n_19604), .b(n_19642), .c(n_19931), .o(n_20779) );
ao12f80 g548866 ( .a(n_21262), .b(n_21261), .c(n_21260), .o(n_22008) );
in01f80 g548867 ( .a(n_20372), .o(n_20436) );
ao12f80 g548868 ( .a(n_19036), .b(n_19374), .c(n_19035), .o(n_20372) );
in01f80 g548869 ( .a(n_20035), .o(n_20075) );
ao12f80 g548870 ( .a(n_18682), .b(n_19060), .c(n_18681), .o(n_20035) );
in01f80 g548871 ( .a(n_20403), .o(n_20775) );
ao12f80 g548872 ( .a(n_19360), .b(n_19663), .c(n_19359), .o(n_20403) );
ao12f80 g548873 ( .a(n_21257), .b(n_21256), .c(n_21255), .o(n_22007) );
in01f80 g548874 ( .a(n_20002), .o(n_20801) );
oa12f80 g548875 ( .a(n_19046), .b(n_19379), .c(n_19045), .o(n_20002) );
oa12f80 g548876 ( .a(n_19598), .b(n_19597), .c(n_19602), .o(n_20752) );
ao12f80 g548877 ( .a(n_20630), .b(n_20629), .c(n_20628), .o(n_21289) );
oa12f80 g548878 ( .a(n_19600), .b(n_19599), .c(n_19601), .o(n_20758) );
oa12f80 g548879 ( .a(n_19593), .b(n_19592), .c(n_19605), .o(n_20757) );
ao12f80 g548880 ( .a(n_21254), .b(n_21253), .c(n_21252), .o(n_22006) );
ao12f80 g548881 ( .a(n_21251), .b(n_21250), .c(n_21249), .o(n_22005) );
oa12f80 g548882 ( .a(n_19608), .b(n_19607), .c(n_19606), .o(n_20771) );
ao12f80 g548883 ( .a(n_20621), .b(n_20620), .c(n_20619), .o(n_21288) );
ao12f80 g548884 ( .a(n_20654), .b(n_20653), .c(n_20652), .o(n_21287) );
ao12f80 g548885 ( .a(n_21236), .b(n_21235), .c(n_21234), .o(n_22004) );
in01f80 g548886 ( .a(n_20058), .o(n_20401) );
oa12f80 g548887 ( .a(n_19056), .b(n_19384), .c(n_19055), .o(n_20058) );
in01f80 g548888 ( .a(n_20034), .o(n_20361) );
ao12f80 g548889 ( .a(n_19038), .b(n_19375), .c(n_19037), .o(n_20034) );
ao12f80 g548890 ( .a(n_20618), .b(n_20617), .c(n_20616), .o(n_21286) );
in01f80 g548891 ( .a(n_20717), .o(n_20770) );
ao12f80 g548892 ( .a(n_19347), .b(n_19658), .c(n_19346), .o(n_20717) );
in01f80 g548893 ( .a(n_20059), .o(n_20433) );
ao12f80 g548894 ( .a(n_19054), .b(n_19383), .c(n_19053), .o(n_20059) );
ao12f80 g548895 ( .a(n_20615), .b(n_20614), .c(n_20613), .o(n_21285) );
in01f80 g548896 ( .a(n_20042), .o(n_20432) );
ao12f80 g548897 ( .a(n_19052), .b(n_19382), .c(n_19051), .o(n_20042) );
ao12f80 g548898 ( .a(n_20292), .b(n_20291), .c(n_20290), .o(n_20979) );
in01f80 g548899 ( .a(n_20978), .o(n_21768) );
oa12f80 g548900 ( .a(n_19934), .b(n_20329), .c(n_19933), .o(n_20978) );
ao12f80 g548901 ( .a(n_21245), .b(n_21244), .c(n_21243), .o(n_22003) );
ao12f80 g548902 ( .a(n_20289), .b(n_20288), .c(n_20287), .o(n_20977) );
in01f80 g548903 ( .a(n_20063), .o(n_20431) );
ao12f80 g548904 ( .a(n_19050), .b(n_19381), .c(n_19049), .o(n_20063) );
in01f80 g548905 ( .a(n_20051), .o(n_20430) );
ao12f80 g548906 ( .a(n_19040), .b(n_19376), .c(n_19039), .o(n_20051) );
ao12f80 g548907 ( .a(n_20612), .b(n_20611), .c(n_20610), .o(n_21284) );
in01f80 g548908 ( .a(n_20395), .o(n_20727) );
oa12f80 g548909 ( .a(n_19353), .b(n_19661), .c(n_19352), .o(n_20395) );
in01f80 g548910 ( .a(n_20061), .o(n_20429) );
ao12f80 g548911 ( .a(n_19048), .b(n_19380), .c(n_19047), .o(n_20061) );
ao12f80 g548912 ( .a(n_21242), .b(n_21241), .c(n_21240), .o(n_22002) );
ao12f80 g548913 ( .a(n_20609), .b(n_20608), .c(n_20607), .o(n_21283) );
in01f80 g548914 ( .a(n_20327), .o(n_21081) );
oa12f80 g548915 ( .a(n_19342), .b(n_19657), .c(n_19341), .o(n_20327) );
ao12f80 g548916 ( .a(n_20286), .b(n_20285), .c(n_20284), .o(n_20976) );
oa12f80 g548917 ( .a(n_20249), .b(n_20248), .c(n_20247), .o(n_21378) );
ao12f80 g548918 ( .a(n_19020), .b(FE_OFN724_n_19019), .c(n_19018), .o(n_19656) );
ao12f80 g548919 ( .a(n_21239), .b(n_21238), .c(n_21237), .o(n_22001) );
oa12f80 g548920 ( .a(n_19915), .b(n_19914), .c(n_19913), .o(n_21042) );
ao12f80 g548921 ( .a(n_20938), .b(n_20937), .c(n_20936), .o(n_21615) );
in01f80 g548922 ( .a(n_20032), .o(n_20427) );
ao12f80 g548923 ( .a(n_19026), .b(n_19369), .c(n_19025), .o(n_20032) );
in01f80 g548924 ( .a(n_20710), .o(n_21035) );
ao12f80 g548925 ( .a(n_19591), .b(n_20003), .c(n_19590), .o(n_20710) );
oa12f80 g548926 ( .a(n_19911), .b(n_19912), .c(n_19910), .o(n_21041) );
ao12f80 g548927 ( .a(n_20260), .b(n_20259), .c(n_20258), .o(n_20975) );
ao12f80 g548928 ( .a(n_20599), .b(n_20598), .c(n_20597), .o(n_21282) );
ao12f80 g548929 ( .a(n_19572), .b(n_19571), .c(n_19570), .o(n_20326) );
in01f80 g548930 ( .a(n_20040), .o(n_20001) );
oa12f80 g548931 ( .a(n_19022), .b(n_19367), .c(n_19021), .o(n_20040) );
in01f80 g548932 ( .a(n_21026), .o(n_21404) );
ao22s80 g548933 ( .a(n_19523), .b(n_13507), .c(n_20669), .d(n_13506), .o(n_21026) );
ao22s80 g548934 ( .a(n_20202), .b(n_21280), .c(n_20201), .d(n_20200), .o(n_21281) );
oa12f80 g548935 ( .a(n_19932), .b(n_19989), .c(n_20253), .o(n_21040) );
in01f80 g548936 ( .a(n_20392), .o(n_20325) );
oa12f80 g548937 ( .a(n_19357), .b(n_19662), .c(n_19356), .o(n_20392) );
ao12f80 g548938 ( .a(n_20596), .b(n_20595), .c(n_20594), .o(n_21279) );
ao22s80 g548939 ( .a(n_20214), .b(n_21613), .c(n_20213), .d(n_20519), .o(n_21614) );
in01f80 g548940 ( .a(n_20368), .o(n_20774) );
ao12f80 g548941 ( .a(n_19349), .b(n_19660), .c(n_19348), .o(n_20368) );
oa12f80 g548942 ( .a(n_19909), .b(n_19908), .c(n_19907), .o(n_21038) );
in01f80 g548943 ( .a(n_20379), .o(n_20426) );
ao12f80 g548944 ( .a(n_19030), .b(n_19371), .c(n_19029), .o(n_20379) );
ao12f80 g548945 ( .a(n_20592), .b(n_20591), .c(n_20590), .o(n_21278) );
oa12f80 g548946 ( .a(n_19344), .b(n_19345), .c(n_19343), .o(n_20425) );
in01f80 g548947 ( .a(n_19678), .o(n_20046) );
ao12f80 g548948 ( .a(n_18680), .b(n_19061), .c(n_18679), .o(n_19678) );
ao12f80 g548949 ( .a(n_20269), .b(n_20268), .c(n_20267), .o(n_20974) );
in01f80 g548950 ( .a(n_21021), .o(n_21392) );
ao22s80 g548951 ( .a(n_19522), .b(n_12544), .c(n_20668), .d(n_12543), .o(n_21021) );
oa12f80 g548952 ( .a(n_19906), .b(n_19905), .c(n_20245), .o(n_21036) );
in01f80 g548953 ( .a(n_20375), .o(n_20423) );
ao12f80 g548954 ( .a(n_19034), .b(n_19373), .c(n_19033), .o(n_20375) );
ao12f80 g548955 ( .a(n_19331), .b(n_19330), .c(n_19329), .o(n_20000) );
in01f80 g548956 ( .a(n_20038), .o(n_20366) );
ao12f80 g548957 ( .a(n_19024), .b(n_19368), .c(n_19023), .o(n_20038) );
ao22s80 g548958 ( .a(n_19879), .b(n_21276), .c(n_19878), .d(n_20198), .o(n_21277) );
in01f80 g548959 ( .a(n_21017), .o(n_21356) );
ao12f80 g548960 ( .a(n_19947), .b(n_20331), .c(n_19946), .o(n_21017) );
ao12f80 g548961 ( .a(n_20584), .b(n_20583), .c(n_20582), .o(n_21275) );
ao22s80 g548962 ( .a(n_20211), .b(n_21273), .c(n_20210), .d(n_20197), .o(n_21274) );
ao12f80 g548963 ( .a(n_19340), .b(n_19654), .c(n_19339), .o(n_19999) );
in01f80 g548964 ( .a(n_19681), .o(n_20054) );
ao12f80 g548965 ( .a(n_18678), .b(n_19059), .c(n_18677), .o(n_19681) );
in01f80 g548966 ( .a(n_20390), .o(n_20420) );
ao12f80 g548967 ( .a(n_19032), .b(n_19372), .c(n_19031), .o(n_20390) );
in01f80 g548968 ( .a(n_21338), .o(n_21388) );
ao12f80 g548969 ( .a(n_19943), .b(n_20330), .c(n_19942), .o(n_21338) );
in01f80 g548970 ( .a(n_20324), .o(n_21077) );
oa12f80 g548971 ( .a(n_19351), .b(n_19659), .c(n_19350), .o(n_20324) );
oa12f80 g548972 ( .a(n_20557), .b(n_20556), .c(n_20558), .o(n_21674) );
ao12f80 g548973 ( .a(n_20580), .b(n_20579), .c(n_20578), .o(n_21272) );
ao12f80 g548974 ( .a(n_19619), .b(n_19618), .c(n_19617), .o(n_20323) );
ao12f80 g548975 ( .a(n_21595), .b(n_21594), .c(n_21593), .o(n_22279) );
oa12f80 g548976 ( .a(n_20244), .b(n_20555), .c(n_20243), .o(n_21352) );
in01f80 g548977 ( .a(n_20387), .o(n_20417) );
ao12f80 g548978 ( .a(n_19028), .b(n_19370), .c(n_19027), .o(n_20387) );
ao12f80 g548979 ( .a(n_19615), .b(n_19614), .c(n_19613), .o(n_20322) );
ao12f80 g548980 ( .a(n_21986), .b(n_21985), .c(n_21984), .o(n_22590) );
oa12f80 g548981 ( .a(n_19904), .b(n_19903), .c(n_19902), .o(n_21032) );
ao12f80 g548982 ( .a(n_19326), .b(n_19335), .c(n_19325), .o(n_19998) );
ao12f80 g548983 ( .a(n_20928), .b(n_20927), .c(n_20926), .o(n_21612) );
oa12f80 g548984 ( .a(n_19594), .b(n_19630), .c(n_19930), .o(n_20734) );
ao12f80 g548985 ( .a(n_20570), .b(n_20569), .c(n_20568), .o(n_21271) );
ao12f80 g548986 ( .a(n_21231), .b(n_21230), .c(n_21229), .o(n_22000) );
in01f80 g548987 ( .a(n_21349), .o(n_21270) );
oa12f80 g548988 ( .a(n_20251), .b(n_20560), .c(n_20660), .o(n_21349) );
ao12f80 g548989 ( .a(n_21226), .b(n_21225), .c(n_21224), .o(n_21999) );
in01f80 g548990 ( .a(n_20048), .o(n_20414) );
ao12f80 g548991 ( .a(n_19044), .b(n_19377), .c(n_19043), .o(n_20048) );
ao12f80 g548992 ( .a(n_19929), .b(n_19928), .c(n_19927), .o(n_20667) );
in01f80 g548993 ( .a(n_21015), .o(n_21029) );
ao12f80 g548994 ( .a(n_19610), .b(n_20004), .c(n_19609), .o(n_21015) );
oa12f80 g548995 ( .a(n_19926), .b(n_19925), .c(n_20242), .o(n_21028) );
in01f80 g548996 ( .a(n_19997), .o(n_20795) );
oa12f80 g548997 ( .a(n_19042), .b(n_19378), .c(n_19041), .o(n_19997) );
oa22f80 g548998 ( .a(n_19521), .b(FE_OFN223_n_21642), .c(n_772), .d(FE_OFN193_n_28928), .o(n_20666) );
oa22f80 g548999 ( .a(FE_OFN1035_n_21194), .b(n_29664), .c(n_1896), .d(FE_OFN347_n_4860), .o(n_22278) );
oa22f80 g549000 ( .a(FE_OFN432_n_20518), .b(n_29664), .c(n_1897), .d(FE_OFN336_n_4860), .o(n_21611) );
oa22f80 g549001 ( .a(n_20196), .b(FE_OFN311_n_3069), .c(n_1245), .d(FE_OFN1174_n_4860), .o(n_21269) );
oa22f80 g549002 ( .a(FE_OFN740_n_20195), .b(n_23291), .c(n_350), .d(FE_OFN95_n_27449), .o(n_21268) );
oa22f80 g549003 ( .a(n_19520), .b(n_23291), .c(n_23), .d(FE_OFN193_n_28928), .o(n_20665) );
oa22f80 g549004 ( .a(n_20517), .b(FE_OFN313_n_3069), .c(n_1457), .d(FE_OFN139_n_27449), .o(n_21610) );
oa22f80 g549005 ( .a(FE_OFN490_n_20516), .b(n_22960), .c(n_210), .d(n_29266), .o(n_21609) );
oa22f80 g549006 ( .a(n_19519), .b(FE_OFN311_n_3069), .c(n_407), .d(FE_OFN1174_n_4860), .o(n_20664) );
oa22f80 g549007 ( .a(FE_OFN590_n_20904), .b(n_29664), .c(n_1765), .d(FE_OFN96_n_27449), .o(n_21998) );
oa22f80 g549008 ( .a(FE_OFN917_n_19297), .b(n_29664), .c(n_1117), .d(FE_OFN347_n_4860), .o(n_20321) );
oa22f80 g549009 ( .a(FE_OFN903_n_20903), .b(n_23291), .c(n_1528), .d(n_29266), .o(n_21997) );
oa22f80 g549010 ( .a(n_20514), .b(FE_OFN299_n_3069), .c(n_1177), .d(FE_OFN136_n_27449), .o(n_21607) );
oa22f80 g549011 ( .a(n_19296), .b(n_29664), .c(n_1478), .d(n_27449), .o(n_20320) );
oa22f80 g549012 ( .a(n_20513), .b(n_29664), .c(n_1366), .d(n_27449), .o(n_21606) );
oa22f80 g549013 ( .a(n_20194), .b(FE_OFN223_n_21642), .c(n_708), .d(FE_OFN330_n_4860), .o(n_21267) );
oa22f80 g549014 ( .a(n_20512), .b(FE_OFN293_n_3069), .c(n_1327), .d(n_29204), .o(n_21605) );
oa22f80 g549015 ( .a(n_20511), .b(FE_OFN300_n_3069), .c(n_118), .d(FE_OFN1110_rst), .o(n_21604) );
oa22f80 g549016 ( .a(n_20902), .b(FE_OFN206_n_28771), .c(n_1362), .d(FE_OFN336_n_4860), .o(n_21996) );
oa22f80 g549017 ( .a(n_20901), .b(FE_OFN253_n_4280), .c(n_1447), .d(FE_OFN136_n_27449), .o(n_21995) );
oa22f80 g549018 ( .a(n_20900), .b(FE_OFN257_n_4280), .c(n_794), .d(n_28607), .o(n_21994) );
oa22f80 g549019 ( .a(n_19861), .b(FE_OFN264_n_4280), .c(n_1919), .d(FE_OFN65_n_27012), .o(n_20973) );
oa22f80 g549020 ( .a(n_19860), .b(FE_OFN253_n_4280), .c(n_334), .d(FE_OFN1119_rst), .o(n_20972) );
oa22f80 g549021 ( .a(n_20896), .b(FE_OFN260_n_4280), .c(n_719), .d(FE_OFN125_n_27449), .o(n_21993) );
oa22f80 g549022 ( .a(n_20899), .b(FE_OFN204_n_28771), .c(n_1476), .d(FE_OFN98_n_27449), .o(n_21992) );
oa22f80 g549023 ( .a(n_20898), .b(FE_OFN206_n_28771), .c(n_1878), .d(FE_OFN1144_n_27012), .o(n_21991) );
oa22f80 g549024 ( .a(n_20895), .b(FE_OFN257_n_4280), .c(n_185), .d(FE_OFN1106_rst), .o(n_21990) );
oa22f80 g549025 ( .a(n_19844), .b(FE_OFN230_n_4162), .c(n_1105), .d(FE_OFN95_n_27449), .o(n_20971) );
oa22f80 g549026 ( .a(n_19859), .b(FE_OFN265_n_4280), .c(n_144), .d(FE_OFN128_n_27449), .o(n_20970) );
oa22f80 g549027 ( .a(n_18992), .b(FE_OFN269_n_4280), .c(n_1465), .d(FE_OFN115_n_27449), .o(n_19996) );
oa22f80 g549028 ( .a(FE_OFN1003_n_19855), .b(FE_OFN266_n_4280), .c(n_728), .d(n_29104), .o(n_20969) );
oa22f80 g549029 ( .a(n_19654), .b(FE_OFN405_n_28303), .c(n_629), .d(FE_OFN92_n_27449), .o(n_19655) );
oa22f80 g549030 ( .a(n_19354), .b(n_4280), .c(n_1495), .d(FE_OFN99_n_27449), .o(n_19653) );
oa22f80 g549031 ( .a(n_20897), .b(n_21988), .c(n_212), .d(n_29104), .o(n_21989) );
oa22f80 g549032 ( .a(n_18997), .b(n_21988), .c(n_1241), .d(n_25680), .o(n_19995) );
oa22f80 g549033 ( .a(n_19858), .b(FE_OFN260_n_4280), .c(n_1782), .d(FE_OFN125_n_27449), .o(n_20968) );
oa22f80 g549034 ( .a(n_19857), .b(FE_OFN171_n_22948), .c(n_1512), .d(FE_OFN98_n_27449), .o(n_20967) );
oa22f80 g549035 ( .a(n_20193), .b(FE_OFN169_n_22948), .c(n_269), .d(FE_OFN130_n_27449), .o(n_21266) );
oa22f80 g549036 ( .a(FE_OFN750_n_20252), .b(FE_OFN173_n_22948), .c(n_886), .d(FE_OFN139_n_27449), .o(n_20663) );
oa22f80 g549037 ( .a(n_20510), .b(FE_OFN254_n_4280), .c(n_156), .d(FE_OFN77_n_27012), .o(n_21603) );
oa22f80 g549038 ( .a(n_19856), .b(FE_OFN169_n_22948), .c(n_232), .d(FE_OFN136_n_27449), .o(n_20966) );
oa22f80 g549039 ( .a(FE_OFN696_n_19853), .b(n_27933), .c(n_1258), .d(FE_OFN63_n_27012), .o(n_20965) );
oa22f80 g549040 ( .a(n_19852), .b(n_27933), .c(n_1297), .d(n_27449), .o(n_20964) );
oa22f80 g549041 ( .a(n_19639), .b(FE_OFN416_n_28303), .c(n_1209), .d(FE_OFN1123_rst), .o(n_19994) );
oa22f80 g549042 ( .a(n_19518), .b(n_28771), .c(n_1276), .d(FE_OFN131_n_27449), .o(n_20662) );
oa22f80 g549043 ( .a(FE_OFN718_n_18993), .b(n_27933), .c(n_875), .d(FE_OFN102_n_27449), .o(n_19993) );
oa22f80 g549044 ( .a(FE_OFN710_n_20192), .b(n_27933), .c(n_644), .d(FE_OFN336_n_4860), .o(n_21265) );
oa22f80 g549045 ( .a(n_20509), .b(FE_OFN299_n_3069), .c(n_927), .d(FE_OFN136_n_27449), .o(n_21602) );
oa22f80 g549046 ( .a(n_19851), .b(FE_OFN206_n_28771), .c(n_652), .d(FE_OFN364_n_4860), .o(n_20963) );
oa22f80 g549047 ( .a(n_19293), .b(n_28771), .c(n_76), .d(FE_OFN138_n_27449), .o(n_20319) );
oa22f80 g549048 ( .a(FE_OFN919_n_19575), .b(FE_OFN309_n_3069), .c(n_1278), .d(FE_OFN190_n_28362), .o(n_19992) );
oa22f80 g549049 ( .a(FE_OFN911_n_19850), .b(n_21988), .c(n_906), .d(FE_OFN347_n_4860), .o(n_20962) );
oa22f80 g549050 ( .a(n_20508), .b(FE_OFN295_n_3069), .c(n_1545), .d(FE_OFN1120_rst), .o(n_21601) );
oa22f80 g549051 ( .a(n_18370), .b(FE_OFN312_n_3069), .c(n_1296), .d(FE_OFN1111_rst), .o(n_19366) );
oa22f80 g549052 ( .a(n_20191), .b(FE_OFN314_n_3069), .c(n_605), .d(FE_OFN1111_rst), .o(n_21264) );
oa22f80 g549053 ( .a(n_18648), .b(n_21988), .c(n_1012), .d(FE_OFN349_n_4860), .o(n_19652) );
oa22f80 g549054 ( .a(n_20660), .b(FE_OFN312_n_3069), .c(n_231), .d(FE_OFN329_n_4860), .o(n_20661) );
oa22f80 g549055 ( .a(n_20507), .b(FE_OFN297_n_3069), .c(n_233), .d(FE_OFN142_n_27449), .o(n_21600) );
oa22f80 g549056 ( .a(n_19288), .b(FE_OFN310_n_3069), .c(n_1524), .d(FE_OFN1143_n_27012), .o(n_20318) );
oa22f80 g549057 ( .a(n_19516), .b(FE_OFN230_n_4162), .c(n_153), .d(FE_OFN102_n_27449), .o(n_20659) );
oa22f80 g549058 ( .a(n_19849), .b(FE_OFN310_n_3069), .c(n_1309), .d(FE_OFN1113_rst), .o(n_20961) );
oa22f80 g549059 ( .a(FE_OFN512_n_19847), .b(n_21988), .c(n_864), .d(FE_OFN68_n_27012), .o(n_20960) );
oa22f80 g549060 ( .a(FE_OFN899_n_19332), .b(n_21988), .c(n_1779), .d(FE_OFN1115_rst), .o(n_19651) );
oa22f80 g549061 ( .a(n_18991), .b(FE_OFN405_n_28303), .c(n_142), .d(FE_OFN60_n_27012), .o(n_19991) );
oa22f80 g549062 ( .a(n_19589), .b(FE_OFN230_n_4162), .c(n_852), .d(FE_OFN102_n_27449), .o(n_19990) );
oa22f80 g549063 ( .a(n_19845), .b(FE_OFN170_n_22948), .c(n_363), .d(n_28607), .o(n_20959) );
oa22f80 g549064 ( .a(n_19287), .b(FE_OFN169_n_22948), .c(n_61), .d(FE_OFN99_n_27449), .o(n_20317) );
oa22f80 g549065 ( .a(n_21193), .b(n_27933), .c(n_564), .d(FE_OFN1109_rst), .o(n_22276) );
oa22f80 g549066 ( .a(n_19286), .b(FE_OFN247_n_4162), .c(n_408), .d(FE_OFN134_n_27449), .o(n_20316) );
oa22f80 g549067 ( .a(n_21571), .b(FE_OFN244_n_4162), .c(n_1924), .d(FE_OFN134_n_27449), .o(n_22589) );
oa22f80 g549068 ( .a(n_19285), .b(FE_OFN239_n_4162), .c(n_802), .d(FE_OFN135_n_27449), .o(n_20315) );
oa22f80 g549069 ( .a(n_20190), .b(FE_OFN239_n_4162), .c(n_1010), .d(FE_OFN130_n_27449), .o(n_21263) );
oa22f80 g549070 ( .a(n_19846), .b(FE_OFN303_n_3069), .c(n_1172), .d(FE_OFN1108_rst), .o(n_20958) );
oa22f80 g549071 ( .a(n_19843), .b(n_27933), .c(n_754), .d(FE_OFN105_n_27449), .o(n_20957) );
oa22f80 g549072 ( .a(FE_OFN518_n_20894), .b(n_27933), .c(n_1706), .d(FE_OFN56_n_27012), .o(n_21987) );
oa22f80 g549073 ( .a(n_20506), .b(n_27933), .c(n_1872), .d(FE_OFN64_n_27012), .o(n_21599) );
oa22f80 g549074 ( .a(n_19842), .b(FE_OFN412_n_28303), .c(n_1870), .d(FE_OFN330_n_4860), .o(n_20956) );
oa22f80 g549075 ( .a(FE_OFN630_n_19358), .b(FE_OFN311_n_3069), .c(n_1858), .d(n_28362), .o(n_19650) );
no02f80 g549153 ( .a(n_21597), .b(n_21596), .o(n_21598) );
na02f80 g549154 ( .a(n_20314), .b(x_in_2_5), .o(n_21320) );
in01f80 g549155 ( .a(n_20657), .o(n_20658) );
no02f80 g549156 ( .a(n_20314), .b(x_in_2_5), .o(n_20657) );
no02f80 g549157 ( .a(n_20954), .b(n_20953), .o(n_20955) );
na02f80 g549158 ( .a(n_20254), .b(x_in_60_4), .o(n_21309) );
na02f80 g549159 ( .a(n_20313), .b(x_in_34_5), .o(n_21303) );
in01f80 g549160 ( .a(n_20655), .o(n_20656) );
no02f80 g549161 ( .a(n_20313), .b(x_in_34_5), .o(n_20655) );
no02f80 g549162 ( .a(n_20951), .b(n_20950), .o(n_20952) );
no02f80 g549163 ( .a(n_20653), .b(n_20652), .o(n_20654) );
no02f80 g549164 ( .a(n_20948), .b(n_20947), .o(n_20949) );
na02f80 g549165 ( .a(n_19989), .b(x_in_8_8), .o(n_21005) );
na02f80 g549166 ( .a(n_19649), .b(x_in_18_5), .o(n_20700) );
in01f80 g549167 ( .a(n_19987), .o(n_19988) );
no02f80 g549168 ( .a(n_19649), .b(x_in_18_5), .o(n_19987) );
no02f80 g549169 ( .a(n_19985), .b(n_19984), .o(n_19986) );
no02f80 g549170 ( .a(n_20650), .b(n_20649), .o(n_20651) );
in01f80 g549171 ( .a(n_19982), .o(n_19983) );
no02f80 g549172 ( .a(n_19612), .b(x_in_50_5), .o(n_19982) );
no02f80 g549173 ( .a(n_19665), .b(n_19364), .o(n_19365) );
na02f80 g549174 ( .a(n_19981), .b(x_in_6_5), .o(n_21004) );
in01f80 g549175 ( .a(n_20311), .o(n_20312) );
no02f80 g549176 ( .a(n_19981), .b(x_in_6_5), .o(n_20311) );
no02f80 g549177 ( .a(n_20647), .b(n_20646), .o(n_20648) );
na02f80 g549178 ( .a(n_19648), .b(x_in_10_5), .o(n_20699) );
in01f80 g549179 ( .a(n_19979), .o(n_19980) );
no02f80 g549180 ( .a(n_19648), .b(x_in_10_5), .o(n_19979) );
na02f80 g549181 ( .a(n_20298), .b(x_in_56_7), .o(n_21311) );
no02f80 g549182 ( .a(n_20309), .b(n_20308), .o(n_20310) );
na02f80 g549183 ( .a(n_19647), .b(x_in_42_5), .o(n_20698) );
in01f80 g549184 ( .a(n_19977), .o(n_19978) );
no02f80 g549185 ( .a(n_19647), .b(x_in_42_5), .o(n_19977) );
na02f80 g549186 ( .a(n_19645), .b(x_in_2_6), .o(n_20692) );
na02f80 g549187 ( .a(n_20281), .b(x_in_26_5), .o(n_21299) );
no02f80 g549188 ( .a(n_20644), .b(n_20643), .o(n_20645) );
no02f80 g549189 ( .a(n_20945), .b(n_20944), .o(n_20946) );
no02f80 g549190 ( .a(n_20641), .b(n_20640), .o(n_20642) );
na02f80 g549191 ( .a(n_19646), .b(x_in_58_5), .o(n_20695) );
in01f80 g549192 ( .a(n_19975), .o(n_19976) );
no02f80 g549193 ( .a(n_19646), .b(x_in_58_5), .o(n_19975) );
na02f80 g549194 ( .a(n_19974), .b(x_in_6_4), .o(n_21001) );
in01f80 g549195 ( .a(n_20306), .o(n_20307) );
no02f80 g549196 ( .a(n_19974), .b(x_in_6_4), .o(n_20306) );
no02f80 g549197 ( .a(n_21261), .b(n_21260), .o(n_21262) );
no02f80 g549198 ( .a(n_19385), .b(n_19057), .o(n_19058) );
in01f80 g549199 ( .a(n_21258), .o(n_21259) );
na02f80 g549200 ( .a(n_20943), .b(n_20219), .o(n_21258) );
no02f80 g549201 ( .a(n_19664), .b(n_19362), .o(n_19363) );
in01f80 g549202 ( .a(n_20304), .o(n_20305) );
na02f80 g549203 ( .a(n_19973), .b(n_19314), .o(n_20304) );
na02f80 g549204 ( .a(n_20303), .b(x_in_22_5), .o(n_21315) );
in01f80 g549205 ( .a(n_20638), .o(n_20639) );
no02f80 g549206 ( .a(n_20303), .b(x_in_22_5), .o(n_20638) );
na02f80 g549207 ( .a(n_20302), .b(x_in_54_5), .o(n_21312) );
in01f80 g549208 ( .a(n_20636), .o(n_20637) );
no02f80 g549209 ( .a(n_20302), .b(x_in_54_5), .o(n_20636) );
in01f80 g549210 ( .a(n_19971), .o(n_19972) );
no02f80 g549211 ( .a(n_19645), .b(x_in_2_6), .o(n_19971) );
na02f80 g549212 ( .a(n_19361), .b(x_in_52_5), .o(n_20347) );
in01f80 g549213 ( .a(n_19643), .o(n_19644) );
no02f80 g549214 ( .a(n_19361), .b(x_in_52_5), .o(n_19643) );
no02f80 g549215 ( .a(n_19663), .b(n_19359), .o(n_19360) );
in01f80 g549216 ( .a(n_19969), .o(n_19970) );
no02f80 g549217 ( .a(n_19642), .b(x_in_22_6), .o(n_19969) );
na02f80 g549218 ( .a(n_19642), .b(x_in_22_6), .o(n_20691) );
no02f80 g549219 ( .a(n_21256), .b(n_21255), .o(n_21257) );
na02f80 g549220 ( .a(n_19952), .b(x_in_40_5), .o(n_20993) );
no02f80 g549221 ( .a(n_20634), .b(n_20633), .o(n_20635) );
na02f80 g549222 ( .a(n_20301), .b(x_in_14_5), .o(n_21317) );
in01f80 g549223 ( .a(n_20631), .o(n_20632) );
no02f80 g549224 ( .a(n_20301), .b(x_in_14_5), .o(n_20631) );
no02f80 g549225 ( .a(n_20629), .b(n_20628), .o(n_20630) );
na02f80 g549226 ( .a(n_20270), .b(x_in_46_5), .o(n_21313) );
no02f80 g549227 ( .a(n_21253), .b(n_21252), .o(n_21254) );
na02f80 g549228 ( .a(n_20300), .b(x_in_30_5), .o(n_21314) );
in01f80 g549229 ( .a(n_20626), .o(n_20627) );
no02f80 g549230 ( .a(n_20300), .b(x_in_30_5), .o(n_20626) );
no02f80 g549231 ( .a(n_21250), .b(n_21249), .o(n_21251) );
in01f80 g549232 ( .a(n_19640), .o(n_19641) );
no02f80 g549233 ( .a(n_19595), .b(x_in_54_6), .o(n_19640) );
no02f80 g549234 ( .a(n_19060), .b(n_18681), .o(n_18682) );
na02f80 g549235 ( .a(n_19595), .b(x_in_54_6), .o(n_20351) );
na02f80 g549236 ( .a(n_20299), .b(x_in_62_5), .o(n_21304) );
in01f80 g549237 ( .a(n_20624), .o(n_20625) );
no02f80 g549238 ( .a(n_20299), .b(x_in_62_5), .o(n_20624) );
na02f80 g549239 ( .a(n_19639), .b(n_19984), .o(n_20789) );
na02f80 g549240 ( .a(n_20255), .b(x_in_60_5), .o(n_21316) );
in01f80 g549241 ( .a(n_20622), .o(n_20623) );
no02f80 g549242 ( .a(n_20298), .b(x_in_56_7), .o(n_20622) );
no02f80 g549243 ( .a(n_20296), .b(n_20295), .o(n_20297) );
in01f80 g549244 ( .a(n_20941), .o(n_20942) );
no02f80 g549245 ( .a(n_20587), .b(x_in_36_5), .o(n_20941) );
no02f80 g549246 ( .a(n_20620), .b(n_20619), .o(n_20621) );
na02f80 g549247 ( .a(n_19384), .b(n_19055), .o(n_19056) );
na02f80 g549248 ( .a(n_19597), .b(x_in_14_6), .o(n_20349) );
in01f80 g549249 ( .a(n_19637), .o(n_19638) );
no02f80 g549250 ( .a(n_19597), .b(x_in_14_6), .o(n_19637) );
no02f80 g549251 ( .a(n_21247), .b(n_21246), .o(n_21248) );
no02f80 g549252 ( .a(n_20617), .b(n_20616), .o(n_20618) );
na02f80 g549253 ( .a(n_19968), .b(x_in_34_6), .o(n_21000) );
in01f80 g549254 ( .a(n_20293), .o(n_20294) );
no02f80 g549255 ( .a(n_19968), .b(x_in_34_6), .o(n_20293) );
no02f80 g549256 ( .a(n_19383), .b(n_19053), .o(n_19054) );
na02f80 g549257 ( .a(FE_OFN630_n_19358), .b(n_19613), .o(n_20415) );
in01f80 g549258 ( .a(n_19635), .o(n_19636) );
no02f80 g549259 ( .a(n_19599), .b(x_in_46_6), .o(n_19635) );
na02f80 g549260 ( .a(n_19599), .b(x_in_46_6), .o(n_20348) );
no02f80 g549261 ( .a(n_20614), .b(n_20613), .o(n_20615) );
no02f80 g549262 ( .a(n_19382), .b(n_19051), .o(n_19052) );
in01f80 g549263 ( .a(n_19966), .o(n_19967) );
no02f80 g549264 ( .a(n_19634), .b(x_in_16_6), .o(n_19966) );
na02f80 g549265 ( .a(n_19634), .b(x_in_16_6), .o(n_20690) );
no02f80 g549266 ( .a(n_20291), .b(n_20290), .o(n_20292) );
no02f80 g549267 ( .a(n_21244), .b(n_21243), .o(n_21245) );
no02f80 g549268 ( .a(n_20288), .b(n_20287), .o(n_20289) );
no02f80 g549269 ( .a(n_19381), .b(n_19049), .o(n_19050) );
na02f80 g549270 ( .a(n_19592), .b(x_in_30_6), .o(n_20346) );
in01f80 g549271 ( .a(n_19632), .o(n_19633) );
no02f80 g549272 ( .a(n_19592), .b(x_in_30_6), .o(n_19632) );
na02f80 g549273 ( .a(n_19631), .b(x_in_18_6), .o(n_20689) );
in01f80 g549274 ( .a(n_19964), .o(n_19965) );
no02f80 g549275 ( .a(n_19631), .b(x_in_18_6), .o(n_19964) );
no02f80 g549276 ( .a(n_20611), .b(n_20610), .o(n_20612) );
na02f80 g549277 ( .a(n_19630), .b(x_in_12_6), .o(n_20685) );
in01f80 g549278 ( .a(n_19962), .o(n_19963) );
no02f80 g549279 ( .a(n_19630), .b(x_in_12_6), .o(n_19962) );
no02f80 g549280 ( .a(n_19380), .b(n_19047), .o(n_19048) );
na02f80 g549281 ( .a(n_19607), .b(x_in_62_6), .o(n_20345) );
in01f80 g549282 ( .a(n_19628), .o(n_19629) );
no02f80 g549283 ( .a(n_19607), .b(x_in_62_6), .o(n_19628) );
no02f80 g549284 ( .a(n_21241), .b(n_21240), .o(n_21242) );
no02f80 g549285 ( .a(n_20608), .b(n_20607), .o(n_20609) );
no02f80 g549286 ( .a(n_20285), .b(n_20284), .o(n_20286) );
na02f80 g549287 ( .a(n_20606), .b(x_in_32_4), .o(n_21633) );
in01f80 g549288 ( .a(n_20939), .o(n_20940) );
no02f80 g549289 ( .a(n_20606), .b(x_in_32_4), .o(n_20939) );
no02f80 g549290 ( .a(n_21238), .b(n_21237), .o(n_21239) );
na02f80 g549291 ( .a(n_20283), .b(x_in_16_5), .o(n_21310) );
in01f80 g549292 ( .a(n_20604), .o(n_20605) );
no02f80 g549293 ( .a(n_20283), .b(x_in_16_5), .o(n_20604) );
no02f80 g549294 ( .a(n_20937), .b(n_20936), .o(n_20938) );
na02f80 g549295 ( .a(n_19627), .b(x_in_50_6), .o(n_20684) );
in01f80 g549296 ( .a(n_19960), .o(n_19961) );
no02f80 g549297 ( .a(n_19627), .b(x_in_50_6), .o(n_19960) );
in01f80 g549298 ( .a(n_20602), .o(n_20603) );
no02f80 g549299 ( .a(n_20282), .b(x_in_48_4), .o(n_20602) );
na02f80 g549300 ( .a(n_20282), .b(x_in_48_4), .o(n_21308) );
in01f80 g549301 ( .a(n_20600), .o(n_20601) );
no02f80 g549302 ( .a(n_20281), .b(x_in_26_5), .o(n_20600) );
no02f80 g549303 ( .a(n_20598), .b(n_20597), .o(n_20599) );
no02f80 g549304 ( .a(n_20279), .b(n_20278), .o(n_20280) );
na02f80 g549305 ( .a(n_20277), .b(n_19541), .o(n_20998) );
na02f80 g549306 ( .a(n_19959), .b(x_in_8_7), .o(n_20996) );
in01f80 g549307 ( .a(n_20275), .o(n_20276) );
no02f80 g549308 ( .a(n_19959), .b(x_in_8_7), .o(n_20275) );
na02f80 g549309 ( .a(n_19662), .b(n_19356), .o(n_19357) );
na02f80 g549310 ( .a(n_20593), .b(x_in_44_7), .o(n_21628) );
in01f80 g549311 ( .a(n_20273), .o(n_20274) );
no02f80 g549312 ( .a(n_19989), .b(x_in_8_8), .o(n_20273) );
in01f80 g549313 ( .a(n_19625), .o(n_19626) );
na02f80 g549314 ( .a(n_19355), .b(n_18669), .o(n_19625) );
no02f80 g549315 ( .a(n_20595), .b(n_20594), .o(n_20596) );
in01f80 g549316 ( .a(n_20934), .o(n_20935) );
no02f80 g549317 ( .a(n_20593), .b(x_in_44_7), .o(n_20934) );
na02f80 g549318 ( .a(n_19958), .b(x_in_40_4), .o(n_20995) );
in01f80 g549319 ( .a(n_20271), .o(n_20272) );
no02f80 g549320 ( .a(n_19958), .b(x_in_40_4), .o(n_20271) );
na02f80 g549321 ( .a(n_19624), .b(x_in_32_5), .o(n_20683) );
in01f80 g549322 ( .a(n_19956), .o(n_19957) );
no02f80 g549323 ( .a(n_19624), .b(x_in_32_5), .o(n_19956) );
no02f80 g549324 ( .a(n_21235), .b(n_21234), .o(n_21236) );
no02f80 g549325 ( .a(n_20591), .b(n_20590), .o(n_20592) );
in01f80 g549326 ( .a(n_20588), .o(n_20589) );
no02f80 g549327 ( .a(n_20270), .b(x_in_46_5), .o(n_20588) );
na02f80 g549328 ( .a(n_20587), .b(x_in_36_5), .o(n_21634) );
no02f80 g549329 ( .a(n_20268), .b(n_20267), .o(n_20269) );
in01f80 g549330 ( .a(n_19954), .o(n_19955) );
na02f80 g549331 ( .a(n_19623), .b(n_19009), .o(n_19954) );
na02f80 g549332 ( .a(n_19953), .b(x_in_56_6), .o(n_20994) );
in01f80 g549333 ( .a(n_20265), .o(n_20266) );
no02f80 g549334 ( .a(n_19953), .b(x_in_56_6), .o(n_20265) );
in01f80 g549335 ( .a(n_20263), .o(n_20264) );
no02f80 g549336 ( .a(n_19952), .b(x_in_40_5), .o(n_20263) );
in01f80 g549337 ( .a(n_19950), .o(n_19951) );
no02f80 g549338 ( .a(n_19622), .b(x_in_10_6), .o(n_19950) );
na02f80 g549339 ( .a(n_19622), .b(x_in_10_6), .o(n_20682) );
in01f80 g549340 ( .a(n_19948), .o(n_19949) );
na02f80 g549341 ( .a(n_19621), .b(n_19013), .o(n_19948) );
na02f80 g549342 ( .a(n_20262), .b(x_in_48_5), .o(n_21300) );
in01f80 g549343 ( .a(n_20585), .o(n_20586) );
no02f80 g549344 ( .a(n_20262), .b(x_in_48_5), .o(n_20585) );
no02f80 g549345 ( .a(n_20331), .b(n_19946), .o(n_19947) );
no02f80 g549346 ( .a(n_20583), .b(n_20582), .o(n_20584) );
na02f80 g549347 ( .a(n_20581), .b(x_in_20_5), .o(n_21637) );
in01f80 g549348 ( .a(n_20932), .o(n_20933) );
no02f80 g549349 ( .a(n_20581), .b(x_in_20_5), .o(n_20932) );
no02f80 g549350 ( .a(n_21985), .b(n_21984), .o(n_21986) );
na02f80 g549351 ( .a(n_19620), .b(x_in_42_6), .o(n_20680) );
in01f80 g549352 ( .a(n_19944), .o(n_19945) );
no02f80 g549353 ( .a(n_19620), .b(x_in_42_6), .o(n_19944) );
no02f80 g549354 ( .a(n_20330), .b(n_19942), .o(n_19943) );
na02f80 g549355 ( .a(n_20931), .b(x_in_36_4), .o(n_22013) );
in01f80 g549356 ( .a(n_21232), .o(n_21233) );
no02f80 g549357 ( .a(n_20931), .b(x_in_36_4), .o(n_21232) );
no02f80 g549358 ( .a(n_20579), .b(n_20578), .o(n_20580) );
no02f80 g549359 ( .a(n_19618), .b(n_19617), .o(n_19619) );
na02f80 g549360 ( .a(n_19379), .b(n_19045), .o(n_19046) );
na02f80 g549361 ( .a(n_19354), .b(n_19617), .o(n_20418) );
no02f80 g549362 ( .a(n_21594), .b(n_21593), .o(n_21595) );
in01f80 g549363 ( .a(n_20576), .o(n_20577) );
na02f80 g549364 ( .a(n_20261), .b(n_19537), .o(n_20576) );
na02f80 g549365 ( .a(n_20575), .b(x_in_20_4), .o(n_21625) );
in01f80 g549366 ( .a(n_20929), .o(n_20930) );
no02f80 g549367 ( .a(n_20575), .b(x_in_20_4), .o(n_20929) );
na02f80 g549368 ( .a(n_19616), .b(x_in_26_6), .o(n_20679) );
in01f80 g549369 ( .a(n_19940), .o(n_19941) );
no02f80 g549370 ( .a(n_19616), .b(x_in_26_6), .o(n_19940) );
no02f80 g549371 ( .a(n_19614), .b(n_19613), .o(n_19615) );
no02f80 g549372 ( .a(n_20259), .b(n_20258), .o(n_20260) );
na02f80 g549373 ( .a(n_19612), .b(x_in_50_5), .o(n_20681) );
na02f80 g549374 ( .a(n_20257), .b(x_in_52_4), .o(n_21298) );
in01f80 g549375 ( .a(n_20573), .o(n_20574) );
no02f80 g549376 ( .a(n_20257), .b(x_in_52_4), .o(n_20573) );
no02f80 g549377 ( .a(n_20927), .b(n_20926), .o(n_20928) );
na02f80 g549378 ( .a(n_20256), .b(x_in_12_5), .o(n_21297) );
in01f80 g549379 ( .a(n_20571), .o(n_20572) );
no02f80 g549380 ( .a(n_20256), .b(x_in_12_5), .o(n_20571) );
no02f80 g549381 ( .a(n_20569), .b(n_20568), .o(n_20570) );
no02f80 g549382 ( .a(n_21230), .b(n_21229), .o(n_21231) );
na02f80 g549383 ( .a(n_20925), .b(x_in_44_6), .o(n_22016) );
in01f80 g549384 ( .a(n_21227), .o(n_21228) );
no02f80 g549385 ( .a(n_20925), .b(x_in_44_6), .o(n_21227) );
no02f80 g549386 ( .a(n_21225), .b(n_21224), .o(n_21226) );
in01f80 g549387 ( .a(n_21222), .o(n_21223) );
na02f80 g549388 ( .a(n_20924), .b(n_20206), .o(n_21222) );
no02f80 g549389 ( .a(n_19377), .b(n_19043), .o(n_19044) );
na02f80 g549390 ( .a(n_19611), .b(x_in_58_6), .o(n_20693) );
in01f80 g549391 ( .a(n_19938), .o(n_19939) );
no02f80 g549392 ( .a(n_19611), .b(x_in_58_6), .o(n_19938) );
in01f80 g549393 ( .a(n_21220), .o(n_21221) );
na02f80 g549394 ( .a(n_20923), .b(n_20204), .o(n_21220) );
in01f80 g549395 ( .a(n_20566), .o(n_20567) );
no02f80 g549396 ( .a(n_20255), .b(x_in_60_5), .o(n_20566) );
in01f80 g549397 ( .a(n_20564), .o(n_20565) );
no02f80 g549398 ( .a(n_20254), .b(x_in_60_4), .o(n_20564) );
na02f80 g549399 ( .a(n_19378), .b(n_19041), .o(n_19042) );
na02f80 g549400 ( .a(n_19661), .b(n_19352), .o(n_19353) );
no02f80 g549401 ( .a(n_19061), .b(n_18679), .o(n_18680) );
no02f80 g549402 ( .a(n_19376), .b(n_19039), .o(n_19040) );
no02f80 g549403 ( .a(n_20004), .b(n_19609), .o(n_19610) );
na02f80 g549404 ( .a(n_19936), .b(n_19935), .o(n_19937) );
na02f80 g549405 ( .a(n_19659), .b(n_19350), .o(n_19351) );
no02f80 g549406 ( .a(n_19660), .b(n_19348), .o(n_19349) );
no02f80 g549407 ( .a(n_19375), .b(n_19037), .o(n_19038) );
na02f80 g549408 ( .a(n_20329), .b(n_19933), .o(n_19934) );
no02f80 g549409 ( .a(n_19374), .b(n_19035), .o(n_19036) );
no02f80 g549410 ( .a(n_19658), .b(n_19346), .o(n_19347) );
no02f80 g549411 ( .a(n_19059), .b(n_18677), .o(n_18678) );
na02f80 g549412 ( .a(n_19607), .b(n_19606), .o(n_19608) );
na02f80 g549413 ( .a(n_18995), .b(n_19605), .o(n_20408) );
na02f80 g549414 ( .a(n_19642), .b(n_19931), .o(n_19604) );
na02f80 g549415 ( .a(n_18999), .b(n_19603), .o(n_20410) );
na02f80 g549416 ( .a(n_18998), .b(n_19602), .o(n_20400) );
na02f80 g549417 ( .a(n_18996), .b(n_19601), .o(n_20409) );
na02f80 g549418 ( .a(n_19599), .b(n_19601), .o(n_19600) );
na02f80 g549419 ( .a(n_18994), .b(n_19606), .o(n_20411) );
na02f80 g549420 ( .a(n_19517), .b(n_20253), .o(n_21343) );
na02f80 g549421 ( .a(n_19989), .b(n_20253), .o(n_19932) );
na02f80 g549422 ( .a(n_19345), .b(n_18043), .o(n_20016) );
na02f80 g549423 ( .a(n_19345), .b(n_19343), .o(n_19344) );
na02f80 g549424 ( .a(n_19597), .b(n_19602), .o(n_19598) );
na02f80 g549425 ( .a(n_19595), .b(n_19603), .o(n_19596) );
na02f80 g549426 ( .a(n_19295), .b(n_19931), .o(n_20729) );
na02f80 g549427 ( .a(n_19294), .b(n_19930), .o(n_20726) );
na02f80 g549428 ( .a(n_19630), .b(n_19930), .o(n_19594) );
na02f80 g549429 ( .a(n_19592), .b(n_19605), .o(n_19593) );
no02f80 g549430 ( .a(n_20003), .b(n_19590), .o(n_19591) );
no02f80 g549431 ( .a(n_19373), .b(n_19033), .o(n_19034) );
no02f80 g549432 ( .a(n_19372), .b(n_19031), .o(n_19032) );
no02f80 g549433 ( .a(n_20562), .b(n_20561), .o(n_20563) );
na02f80 g549434 ( .a(FE_OFN751_n_20252), .b(n_20561), .o(n_21341) );
no02f80 g549435 ( .a(n_20560), .b(n_20593), .o(n_21624) );
na02f80 g549436 ( .a(n_20560), .b(n_20660), .o(n_20251) );
na02f80 g549437 ( .a(n_19657), .b(n_19341), .o(n_19342) );
no02f80 g549438 ( .a(n_19371), .b(n_19029), .o(n_19030) );
no02f80 g549439 ( .a(n_19370), .b(n_19027), .o(n_19028) );
no02f80 g549440 ( .a(n_19369), .b(n_19025), .o(n_19026) );
no02f80 g549441 ( .a(n_19928), .b(n_19927), .o(n_19929) );
na02f80 g549442 ( .a(n_19589), .b(n_19927), .o(n_20722) );
no02f80 g549443 ( .a(n_19368), .b(n_19023), .o(n_19024) );
no02f80 g549444 ( .a(n_19654), .b(n_19339), .o(n_19340) );
no02f80 g549445 ( .a(n_18647), .b(n_19339), .o(n_20053) );
na02f80 g549446 ( .a(n_19367), .b(n_19021), .o(n_19022) );
no02f80 g549447 ( .a(FE_OFN1061_n_19587), .b(n_19586), .o(n_19588) );
na02f80 g549448 ( .a(n_19925), .b(n_20242), .o(n_19926) );
in01f80 g549449 ( .a(n_19924), .o(n_20371) );
no02f80 g549450 ( .a(n_19645), .b(n_19585), .o(n_19924) );
na02f80 g549451 ( .a(n_19337), .b(n_19585), .o(n_19338) );
in01f80 g549452 ( .a(n_20250), .o(n_20716) );
no02f80 g549453 ( .a(n_19968), .b(n_19923), .o(n_20250) );
ao12f80 g549454 ( .a(n_11575), .b(n_19336), .c(n_12511), .o(n_20357) );
na02f80 g549455 ( .a(n_19564), .b(n_18866), .o(n_20394) );
na02f80 g549456 ( .a(n_19583), .b(n_18880), .o(n_20393) );
na02f80 g549457 ( .a(n_19583), .b(n_19582), .o(n_19584) );
in01f80 g549458 ( .a(n_19922), .o(n_20374) );
no02f80 g549459 ( .a(n_19622), .b(n_19581), .o(n_19922) );
in01f80 g549460 ( .a(n_19921), .o(n_20389) );
no02f80 g549461 ( .a(n_19620), .b(n_19580), .o(n_19921) );
in01f80 g549462 ( .a(n_19920), .o(n_20386) );
no02f80 g549463 ( .a(n_19616), .b(n_19579), .o(n_19920) );
na02f80 g549464 ( .a(n_19577), .b(n_18872), .o(n_20378) );
na02f80 g549465 ( .a(n_19577), .b(n_19576), .o(n_19578) );
in01f80 g549466 ( .a(n_19919), .o(n_20382) );
na02f80 g549467 ( .a(n_19575), .b(n_19916), .o(n_19919) );
no02f80 g549468 ( .a(FE_OFN918_n_19575), .b(n_19916), .o(n_19918) );
no02f80 g549469 ( .a(n_19335), .b(n_18588), .o(n_20360) );
na02f80 g549470 ( .a(n_19573), .b(n_19923), .o(n_19574) );
na02f80 g549471 ( .a(n_20248), .b(n_19459), .o(n_20381) );
na02f80 g549472 ( .a(n_20248), .b(n_20247), .o(n_20249) );
na02f80 g549473 ( .a(n_19333), .b(n_19580), .o(n_19334) );
no02f80 g549474 ( .a(FE_OFN724_n_19019), .b(n_19018), .o(n_19020) );
no02f80 g549475 ( .a(FE_OFN724_n_19019), .b(n_18330), .o(n_20045) );
na02f80 g549476 ( .a(n_19914), .b(n_19184), .o(n_20377) );
na02f80 g549477 ( .a(n_19914), .b(n_19913), .o(n_19915) );
na02f80 g549478 ( .a(n_19912), .b(n_19183), .o(n_21025) );
na02f80 g549479 ( .a(n_19912), .b(n_19910), .o(n_19911) );
no02f80 g549480 ( .a(n_19571), .b(n_19570), .o(n_19572) );
in01f80 g549481 ( .a(n_19569), .o(n_20039) );
na02f80 g549482 ( .a(FE_OFN899_n_19332), .b(n_19570), .o(n_19569) );
no02f80 g549483 ( .a(FE_OFN1061_n_19587), .b(n_18879), .o(n_20719) );
ao12f80 g549484 ( .a(n_8404), .b(n_19568), .c(n_9562), .o(n_20370) );
na02f80 g549485 ( .a(n_19908), .b(n_19182), .o(n_20709) );
na02f80 g549486 ( .a(n_19908), .b(n_19907), .o(n_19909) );
in01f80 g549487 ( .a(n_20673), .o(n_20246) );
na02f80 g549488 ( .a(n_19291), .b(n_12624), .o(n_20673) );
in01f80 g549489 ( .a(n_20559), .o(n_21019) );
no02f80 g549490 ( .a(n_20298), .b(n_20245), .o(n_20559) );
na02f80 g549491 ( .a(n_19905), .b(n_20245), .o(n_19906) );
no02f80 g549492 ( .a(n_19330), .b(n_19329), .o(n_19331) );
no02f80 g549493 ( .a(n_19330), .b(n_18589), .o(n_20365) );
na02f80 g549494 ( .a(n_19901), .b(n_19566), .o(n_19567) );
na02f80 g549495 ( .a(n_19327), .b(n_19579), .o(n_19328) );
in01f80 g549496 ( .a(n_20922), .o(n_21337) );
no02f80 g549497 ( .a(n_20587), .b(n_20558), .o(n_20922) );
na02f80 g549498 ( .a(n_20556), .b(n_20558), .o(n_20557) );
na02f80 g549499 ( .a(n_20555), .b(n_19772), .o(n_21336) );
na02f80 g549500 ( .a(n_20555), .b(n_20243), .o(n_20244) );
na02f80 g549501 ( .a(n_19903), .b(n_19179), .o(n_20037) );
na02f80 g549502 ( .a(n_19903), .b(n_19902), .o(n_19904) );
no02f80 g549503 ( .a(n_19335), .b(n_19325), .o(n_19326) );
na02f80 g549504 ( .a(n_19901), .b(n_19177), .o(n_20708) );
na02f80 g549505 ( .a(n_19564), .b(n_19563), .o(n_19565) );
na02f80 g549506 ( .a(n_19323), .b(n_19581), .o(n_19324) );
in01f80 g549507 ( .a(n_20554), .o(n_21014) );
no02f80 g549508 ( .a(n_20255), .b(n_20242), .o(n_20554) );
in01f80 g549509 ( .a(n_21759), .o(n_21592) );
oa12f80 g549510 ( .a(n_20221), .b(n_19510), .c(n_20130), .o(n_21759) );
in01f80 g549511 ( .a(n_21756), .o(n_21591) );
oa12f80 g549512 ( .a(n_20208), .b(n_19508), .c(n_20127), .o(n_21756) );
in01f80 g549513 ( .a(n_21751), .o(n_21590) );
oa12f80 g549514 ( .a(n_19883), .b(n_19269), .c(n_20128), .o(n_21751) );
in01f80 g549515 ( .a(n_21745), .o(n_21589) );
oa12f80 g549516 ( .a(n_19872), .b(n_19267), .c(n_20126), .o(n_21745) );
in01f80 g549517 ( .a(n_21731), .o(n_21588) );
oa12f80 g549518 ( .a(n_19550), .b(n_18962), .c(n_20129), .o(n_21731) );
in01f80 g549519 ( .a(n_21742), .o(n_21587) );
oa12f80 g549520 ( .a(n_19554), .b(n_18973), .c(n_20124), .o(n_21742) );
in01f80 g549521 ( .a(n_21395), .o(n_21219) );
oa12f80 g549522 ( .a(n_19556), .b(n_19771), .c(n_18971), .o(n_21395) );
ao12f80 g549523 ( .a(n_12469), .b(n_19017), .c(n_13614), .o(n_20031) );
in01f80 g549524 ( .a(n_21375), .o(n_21218) );
oa12f80 g549525 ( .a(n_19553), .b(n_19769), .c(n_18967), .o(n_21375) );
in01f80 g549526 ( .a(n_20921), .o(n_22026) );
ao12f80 g549527 ( .a(n_17795), .b(n_20545), .c(n_18358), .o(n_20921) );
in01f80 g549528 ( .a(n_21401), .o(n_21217) );
oa12f80 g549529 ( .a(n_20526), .b(n_19812), .c(n_19774), .o(n_21401) );
in01f80 g549530 ( .a(n_20920), .o(n_22028) );
oa12f80 g549531 ( .a(n_19429), .b(n_20553), .c(n_18782), .o(n_20920) );
in01f80 g549532 ( .a(n_21748), .o(n_21216) );
oa12f80 g549533 ( .a(n_20530), .b(n_19810), .c(n_19767), .o(n_21748) );
in01f80 g549534 ( .a(n_21728), .o(n_21215) );
oa12f80 g549535 ( .a(n_20528), .b(n_19808), .c(n_19766), .o(n_21728) );
in01f80 g549536 ( .a(n_21708), .o(n_21586) );
oa12f80 g549537 ( .a(n_19551), .b(n_18965), .c(n_20117), .o(n_21708) );
in01f80 g549538 ( .a(n_21385), .o(n_21214) );
oa12f80 g549539 ( .a(n_19316), .b(n_19764), .c(n_18639), .o(n_21385) );
in01f80 g549540 ( .a(n_21722), .o(n_21585) );
oa12f80 g549541 ( .a(n_19885), .b(n_19263), .c(n_20125), .o(n_21722) );
in01f80 g549542 ( .a(n_21725), .o(n_21584) );
oa12f80 g549543 ( .a(n_19888), .b(n_19236), .c(n_20123), .o(n_21725) );
in01f80 g549544 ( .a(n_21353), .o(n_21213) );
oa12f80 g549545 ( .a(n_19555), .b(n_19770), .c(n_18969), .o(n_21353) );
in01f80 g549546 ( .a(n_21713), .o(n_21212) );
oa12f80 g549547 ( .a(n_20524), .b(n_19806), .c(n_19759), .o(n_21713) );
in01f80 g549548 ( .a(n_21719), .o(n_21211) );
oa12f80 g549549 ( .a(n_20529), .b(n_19804), .c(n_19765), .o(n_21719) );
in01f80 g549550 ( .a(n_21716), .o(n_21210) );
oa12f80 g549551 ( .a(n_20531), .b(n_19802), .c(n_19763), .o(n_21716) );
in01f80 g549552 ( .a(n_21736), .o(n_21209) );
oa12f80 g549553 ( .a(n_20520), .b(n_19800), .c(n_19762), .o(n_21736) );
in01f80 g549554 ( .a(n_20241), .o(n_21333) );
ao12f80 g549555 ( .a(n_2162), .b(n_19897), .c(n_2748), .o(n_20241) );
in01f80 g549556 ( .a(n_22034), .o(n_21983) );
oa12f80 g549557 ( .a(n_20527), .b(n_19798), .c(n_20478), .o(n_22034) );
in01f80 g549558 ( .a(n_21208), .o(n_22290) );
ao12f80 g549559 ( .a(n_17418), .b(n_20912), .c(n_18002), .o(n_21208) );
in01f80 g549560 ( .a(n_21703), .o(n_21583) );
oa12f80 g549561 ( .a(n_19549), .b(n_18959), .c(n_20122), .o(n_21703) );
in01f80 g549562 ( .a(n_22304), .o(n_22275) );
oa12f80 g549563 ( .a(n_19884), .b(n_19252), .c(n_20878), .o(n_22304) );
in01f80 g549564 ( .a(n_21700), .o(n_21582) );
oa12f80 g549565 ( .a(n_19548), .b(n_18956), .c(n_20121), .o(n_21700) );
in01f80 g549566 ( .a(n_21382), .o(n_21207) );
oa12f80 g549567 ( .a(n_19547), .b(n_18954), .c(n_19761), .o(n_21382) );
oa12f80 g549568 ( .a(n_10750), .b(n_19322), .c(n_11937), .o(n_20050) );
in01f80 g549569 ( .a(n_21697), .o(n_21581) );
oa12f80 g549570 ( .a(n_19546), .b(n_18952), .c(n_20120), .o(n_21697) );
in01f80 g549571 ( .a(n_21379), .o(n_21206) );
oa12f80 g549572 ( .a(n_19544), .b(n_18950), .c(n_19760), .o(n_21379) );
in01f80 g549573 ( .a(n_21686), .o(n_21580) );
oa12f80 g549574 ( .a(n_19882), .b(n_19241), .c(n_20119), .o(n_21686) );
in01f80 g549575 ( .a(n_21694), .o(n_21579) );
oa12f80 g549576 ( .a(n_19545), .b(n_18947), .c(n_20118), .o(n_21694) );
in01f80 g549577 ( .a(n_20552), .o(n_21650) );
oa12f80 g549578 ( .a(n_16188), .b(n_20234), .c(n_15658), .o(n_20552) );
in01f80 g549579 ( .a(n_22043), .o(n_20919) );
oa12f80 g549580 ( .a(n_20525), .b(n_19793), .c(n_19185), .o(n_22043) );
in01f80 g549581 ( .a(n_21689), .o(n_20918) );
oa12f80 g549582 ( .a(n_20215), .b(n_19489), .c(n_19455), .o(n_21689) );
in01f80 g549583 ( .a(n_21683), .o(n_21578) );
oa12f80 g549584 ( .a(n_19539), .b(n_18941), .c(n_20116), .o(n_21683) );
in01f80 g549585 ( .a(n_20240), .o(n_21330) );
oa12f80 g549586 ( .a(n_3155), .b(n_19895), .c(n_2166), .o(n_20240) );
in01f80 g549587 ( .a(n_21739), .o(n_21205) );
oa12f80 g549588 ( .a(n_20209), .b(n_19758), .c(n_19506), .o(n_21739) );
in01f80 g549589 ( .a(n_21204), .o(n_22288) );
oa12f80 g549590 ( .a(n_19783), .b(n_20917), .c(n_19137), .o(n_21204) );
in01f80 g549591 ( .a(n_21364), .o(n_20551) );
oa12f80 g549592 ( .a(n_19880), .b(n_19220), .c(n_19181), .o(n_21364) );
in01f80 g549593 ( .a(n_21361), .o(n_21203) );
oa12f80 g549594 ( .a(n_19538), .b(n_18935), .c(n_19756), .o(n_21361) );
in01f80 g549595 ( .a(n_20239), .o(n_21327) );
oa12f80 g549596 ( .a(n_18934), .b(n_19900), .c(n_18307), .o(n_20239) );
ao12f80 g549597 ( .a(n_13128), .b(n_19321), .c(n_14276), .o(n_20358) );
in01f80 g549598 ( .a(n_21677), .o(n_21577) );
oa12f80 g549599 ( .a(n_19534), .b(n_20115), .c(n_18930), .o(n_21677) );
in01f80 g549600 ( .a(n_20916), .o(n_22024) );
oa12f80 g549601 ( .a(n_18236), .b(n_20540), .c(n_17685), .o(n_20916) );
in01f80 g549602 ( .a(n_22046), .o(n_21982) );
oa12f80 g549603 ( .a(n_20220), .b(n_19483), .c(n_20477), .o(n_22046) );
in01f80 g549604 ( .a(n_20550), .o(n_21645) );
oa12f80 g549605 ( .a(n_15899), .b(n_20229), .c(n_15278), .o(n_20550) );
in01f80 g549606 ( .a(n_21671), .o(n_21576) );
oa12f80 g549607 ( .a(n_19533), .b(n_20114), .c(n_18925), .o(n_21671) );
in01f80 g549608 ( .a(n_22299), .o(n_21981) );
oa12f80 g549609 ( .a(n_20906), .b(n_20146), .c(n_20480), .o(n_22299) );
in01f80 g549610 ( .a(n_22037), .o(n_21980) );
oa12f80 g549611 ( .a(n_21195), .b(n_20487), .c(n_20479), .o(n_22037) );
in01f80 g549612 ( .a(n_21663), .o(n_21575) );
oa12f80 g549613 ( .a(n_19532), .b(n_20113), .c(n_18920), .o(n_21663) );
in01f80 g549614 ( .a(n_21666), .o(n_20549) );
oa12f80 g549615 ( .a(n_20207), .b(n_19178), .c(n_19478), .o(n_21666) );
in01f80 g549616 ( .a(n_21660), .o(n_21202) );
oa12f80 g549617 ( .a(n_20521), .b(n_19776), .c(n_19755), .o(n_21660) );
in01f80 g549618 ( .a(n_20915), .o(n_22030) );
oa12f80 g549619 ( .a(n_19778), .b(n_20548), .c(n_19133), .o(n_20915) );
in01f80 g549620 ( .a(n_20914), .o(n_22022) );
oa12f80 g549621 ( .a(n_19434), .b(n_20547), .c(n_18758), .o(n_20914) );
in01f80 g549622 ( .a(n_21389), .o(n_21201) );
oa12f80 g549623 ( .a(n_19552), .b(n_19754), .c(n_18939), .o(n_21389) );
in01f80 g549624 ( .a(n_21680), .o(n_21574) );
oa12f80 g549625 ( .a(n_19873), .b(n_19190), .c(n_20112), .o(n_21680) );
in01f80 g549626 ( .a(n_21762), .o(n_21573) );
oa12f80 g549627 ( .a(n_20907), .b(n_20135), .c(n_20131), .o(n_21762) );
oa12f80 g549628 ( .a(n_8834), .b(n_20238), .c(n_10345), .o(n_21022) );
oa12f80 g549629 ( .a(n_5129), .b(n_17810), .c(n_6648), .o(n_18683) );
ao12f80 g549630 ( .a(n_9866), .b(n_18676), .c(n_11173), .o(n_19677) );
na03f80 g549631 ( .a(n_19935), .b(n_19936), .c(n_12890), .o(n_20237) );
ao12f80 g549632 ( .a(n_3675), .b(n_19016), .c(n_19015), .o(n_20030) );
in01f80 g549633 ( .a(n_19320), .o(n_20354) );
oa22f80 g549634 ( .a(n_19016), .b(n_6292), .c(n_18045), .d(n_19015), .o(n_19320) );
ao12f80 g549635 ( .a(n_11988), .b(n_19014), .c(n_13113), .o(n_20029) );
ao12f80 g549636 ( .a(n_19531), .b(n_19530), .c(n_19529), .o(n_20236) );
in01f80 g549637 ( .a(FE_OFN1031_n_19666), .o(n_20006) );
ao12f80 g549638 ( .a(n_18394), .b(n_18676), .c(n_18393), .o(n_19666) );
in01f80 g549639 ( .a(n_20009), .o(n_20350) );
ao12f80 g549640 ( .a(n_18671), .b(n_19017), .c(n_18670), .o(n_20009) );
ao12f80 g549641 ( .a(n_18659), .b(n_18660), .c(n_18658), .o(n_19319) );
oa12f80 g549642 ( .a(n_19305), .b(n_19304), .c(n_19303), .o(n_20694) );
ao22s80 g549643 ( .a(n_20912), .b(n_18262), .c(n_19768), .d(n_18261), .o(n_20913) );
ao22s80 g549644 ( .a(n_19742), .b(n_20553), .c(n_19741), .d(n_19457), .o(n_20911) );
in01f80 g549645 ( .a(n_19899), .o(n_21009) );
oa12f80 g549646 ( .a(n_19005), .b(n_19336), .c(n_19004), .o(n_19899) );
ao22s80 g549647 ( .a(n_18619), .b(n_20545), .c(n_18618), .d(n_19456), .o(n_20546) );
ao22s80 g549648 ( .a(n_19897), .b(n_3831), .c(n_18861), .d(n_3830), .o(n_19898) );
in01f80 g549649 ( .a(n_20344), .o(n_20687) );
ao12f80 g549650 ( .a(n_19011), .b(n_19322), .c(n_19010), .o(n_20344) );
ao22s80 g549651 ( .a(n_20234), .b(n_16419), .c(n_19175), .d(n_16418), .o(n_20235) );
ao12f80 g549652 ( .a(n_19543), .b(n_19891), .c(n_19542), .o(n_20233) );
in01f80 g549653 ( .a(n_18395), .o(n_19388) );
oa12f80 g549654 ( .a(n_17496), .b(n_17810), .c(n_17495), .o(n_18395) );
ao12f80 g549655 ( .a(n_19864), .b(n_19863), .c(n_19862), .o(n_20544) );
in01f80 g549656 ( .a(n_21307), .o(n_21623) );
oa12f80 g549657 ( .a(n_19866), .b(n_20238), .c(n_19865), .o(n_21307) );
ao22s80 g549658 ( .a(n_19895), .b(n_4008), .c(n_18860), .d(n_4007), .o(n_19896) );
ao12f80 g549659 ( .a(n_19868), .b(n_20226), .c(n_19867), .o(n_20543) );
in01f80 g549660 ( .a(FE_OFN498_n_20677), .o(n_20987) );
ao12f80 g549661 ( .a(n_19312), .b(n_19568), .c(n_19311), .o(n_20677) );
ao12f80 g549662 ( .a(n_18665), .b(n_18664), .c(n_18663), .o(n_19318) );
in01f80 g549663 ( .a(n_20405), .o(n_19894) );
oa12f80 g549664 ( .a(n_19003), .b(n_19290), .c(n_19002), .o(n_20405) );
in01f80 g549665 ( .a(n_20014), .o(n_19672) );
ao12f80 g549666 ( .a(n_18094), .b(n_18093), .c(n_18092), .o(n_20014) );
oa12f80 g549667 ( .a(n_18392), .b(n_18391), .c(n_18666), .o(n_19671) );
ao12f80 g549668 ( .a(n_10700), .b(n_18598), .c(n_11831), .o(n_20336) );
ao12f80 g549669 ( .a(n_19527), .b(n_19526), .c(n_19525), .o(n_20232) );
in01f80 g549670 ( .a(n_20333), .o(n_19893) );
oa12f80 g549671 ( .a(n_19007), .b(n_19321), .c(n_19006), .o(n_20333) );
ao22s80 g549672 ( .a(n_20149), .b(n_20917), .c(n_20148), .d(n_19757), .o(n_21200) );
ao22s80 g549673 ( .a(n_19219), .b(n_19900), .c(n_19218), .d(n_18859), .o(n_20231) );
in01f80 g549674 ( .a(n_20017), .o(n_19562) );
oa12f80 g549675 ( .a(n_18662), .b(n_19014), .c(n_18661), .o(n_20017) );
ao12f80 g549676 ( .a(n_19877), .b(n_19876), .c(n_19875), .o(n_20542) );
ao22s80 g549677 ( .a(n_20229), .b(n_16176), .c(n_19174), .d(n_16175), .o(n_20230) );
ao22s80 g549678 ( .a(n_20540), .b(n_18470), .c(n_19453), .d(n_18469), .o(n_20541) );
ao12f80 g549679 ( .a(n_18097), .b(n_18096), .c(n_18095), .o(n_18675) );
ao22s80 g549680 ( .a(n_20145), .b(n_20548), .c(n_20144), .d(n_19452), .o(n_21199) );
oa12f80 g549681 ( .a(n_19308), .b(n_19307), .c(n_19306), .o(n_20678) );
ao22s80 g549682 ( .a(n_19744), .b(n_20547), .c(n_19743), .d(n_19451), .o(n_20910) );
oa22f80 g549683 ( .a(n_19753), .b(FE_OFN314_n_3069), .c(n_532), .d(FE_OFN330_n_4860), .o(n_20909) );
oa22f80 g549684 ( .a(n_19172), .b(n_27933), .c(n_1881), .d(FE_OFN96_n_27449), .o(n_20228) );
oa22f80 g549685 ( .a(n_18325), .b(FE_OFN300_n_3069), .c(n_48), .d(FE_OFN1110_rst), .o(n_19317) );
oa22f80 g549686 ( .a(n_20226), .b(FE_OFN406_n_28303), .c(n_1467), .d(FE_OFN76_n_27012), .o(n_20227) );
oa22f80 g549687 ( .a(n_18577), .b(FE_OFN300_n_3069), .c(n_573), .d(FE_OFN1110_rst), .o(n_19561) );
oa22f80 g549688 ( .a(n_19309), .b(FE_OFN1152_n_3069), .c(n_192), .d(FE_OFN1182_rst), .o(n_19560) );
oa22f80 g549689 ( .a(n_19450), .b(FE_OFN311_n_3069), .c(n_833), .d(FE_OFN122_n_27449), .o(n_20539) );
oa22f80 g549690 ( .a(n_19449), .b(FE_OFN400_n_28303), .c(n_1373), .d(FE_OFN1108_rst), .o(n_20538) );
oa22f80 g549691 ( .a(n_20111), .b(FE_OFN257_n_4280), .c(n_1738), .d(FE_OFN1108_rst), .o(n_21198) );
oa22f80 g549692 ( .a(n_18390), .b(FE_OFN249_n_4162), .c(n_1186), .d(FE_OFN92_n_27449), .o(n_18674) );
oa22f80 g549693 ( .a(n_19302), .b(FE_OFN236_n_4162), .c(n_1323), .d(rst), .o(n_19559) );
oa22f80 g549694 ( .a(n_19171), .b(FE_OFN268_n_4280), .c(n_613), .d(FE_OFN72_n_27012), .o(n_20225) );
oa22f80 g549695 ( .a(n_18581), .b(FE_OFN400_n_28303), .c(n_165), .d(FE_OFN20_n_27452), .o(n_19558) );
oa22f80 g549696 ( .a(n_19891), .b(FE_OFN413_n_28303), .c(n_788), .d(FE_OFN1121_rst), .o(n_19892) );
oa22f80 g549697 ( .a(n_18857), .b(FE_OFN259_n_4280), .c(n_893), .d(FE_OFN1120_rst), .o(n_19890) );
oa22f80 g549698 ( .a(FE_OFN586_n_19447), .b(n_21988), .c(n_1640), .d(FE_OFN1115_rst), .o(n_20536) );
oa22f80 g549699 ( .a(FE_OFN540_n_17809), .b(n_21988), .c(n_1126), .d(FE_OFN347_n_4860), .o(n_18098) );
oa22f80 g549700 ( .a(n_18579), .b(FE_OFN259_n_4280), .c(n_881), .d(FE_OFN130_n_27449), .o(n_19557) );
oa22f80 g549701 ( .a(n_19446), .b(FE_OFN406_n_28303), .c(n_1802), .d(FE_OFN355_n_4860), .o(n_20534) );
oa22f80 g549702 ( .a(n_19168), .b(FE_OFN260_n_4280), .c(n_545), .d(FE_OFN94_n_27449), .o(n_20224) );
oa22f80 g549703 ( .a(n_19752), .b(FE_OFN314_n_3069), .c(n_898), .d(FE_OFN124_n_27449), .o(n_20908) );
oa22f80 g549704 ( .a(FE_OFN660_n_19445), .b(n_21988), .c(n_314), .d(n_27449), .o(n_20533) );
oa22f80 g549705 ( .a(n_19167), .b(FE_OFN258_n_4280), .c(n_275), .d(FE_OFN77_n_27012), .o(n_20223) );
oa22f80 g549706 ( .a(n_18855), .b(FE_OFN266_n_4280), .c(n_1959), .d(FE_OFN190_n_28362), .o(n_19889) );
oa22f80 g549707 ( .a(FE_OFN767_n_20476), .b(n_21988), .c(n_416), .d(n_25680), .o(n_21572) );
oa22f80 g549708 ( .a(n_19166), .b(FE_OFN311_n_3069), .c(n_1082), .d(FE_OFN134_n_27449), .o(n_20222) );
oa22f80 g549709 ( .a(FE_OFN614_n_20110), .b(n_22960), .c(n_1123), .d(FE_OFN336_n_4860), .o(n_21197) );
oa22f80 g549710 ( .a(FE_OFN536_n_17798), .b(n_22960), .c(n_1436), .d(FE_OFN335_n_4860), .o(n_18673) );
oa22f80 g549711 ( .a(n_19444), .b(FE_OFN223_n_21642), .c(n_635), .d(FE_OFN1111_rst), .o(n_20532) );
oa22f80 g549712 ( .a(FE_OFN688_n_20109), .b(FE_OFN235_n_4162), .c(n_168), .d(n_29264), .o(n_21196) );
na02f80 g549758 ( .a(n_20531), .b(n_19803), .o(n_21250) );
na02f80 g549759 ( .a(n_19888), .b(n_19237), .o(n_20634) );
na02f80 g549760 ( .a(n_20221), .b(n_19511), .o(n_20954) );
na02f80 g549761 ( .a(n_20220), .b(n_19484), .o(n_20951) );
na02f80 g549762 ( .a(n_19556), .b(n_18972), .o(n_20309) );
na02f80 g549763 ( .a(n_19555), .b(n_18970), .o(n_20296) );
na02f80 g549764 ( .a(n_19554), .b(n_18974), .o(n_20644) );
na02f80 g549765 ( .a(n_18672), .b(x_in_24_7), .o(n_19621) );
in01f80 g549766 ( .a(n_19012), .o(n_19013) );
no02f80 g549767 ( .a(n_18672), .b(x_in_24_7), .o(n_19012) );
no02f80 g549768 ( .a(n_19017), .b(n_18670), .o(n_18671) );
na02f80 g549769 ( .a(n_19553), .b(n_18968), .o(n_20279) );
in01f80 g549770 ( .a(n_18668), .o(n_18669) );
no02f80 g549771 ( .a(n_19343), .b(x_in_24_8), .o(n_18668) );
na02f80 g549772 ( .a(n_19887), .b(x_in_38_7), .o(n_20943) );
in01f80 g549773 ( .a(n_20218), .o(n_20219) );
no02f80 g549774 ( .a(n_19887), .b(x_in_38_7), .o(n_20218) );
in01f80 g549775 ( .a(n_20216), .o(n_20217) );
na02f80 g549776 ( .a(n_19886), .b(n_19193), .o(n_20216) );
na02f80 g549777 ( .a(n_19343), .b(x_in_24_8), .o(n_19355) );
na02f80 g549778 ( .a(n_20530), .b(n_19811), .o(n_21261) );
na02f80 g549779 ( .a(n_19552), .b(n_18940), .o(n_20259) );
na02f80 g549780 ( .a(n_19885), .b(n_19264), .o(n_20629) );
na02f80 g549781 ( .a(n_20529), .b(n_19805), .o(n_21253) );
na02f80 g549782 ( .a(n_19551), .b(n_18966), .o(n_20653) );
na02f80 g549783 ( .a(n_20528), .b(n_19809), .o(n_21256) );
na02f80 g549784 ( .a(n_20527), .b(n_19799), .o(n_21235) );
na02f80 g549785 ( .a(n_20526), .b(n_19813), .o(n_21247) );
na02f80 g549786 ( .a(n_19550), .b(n_18963), .o(n_20620) );
na02f80 g549787 ( .a(n_19549), .b(n_18960), .o(n_20617) );
na02f80 g549788 ( .a(n_19548), .b(n_18957), .o(n_20614) );
na02f80 g549789 ( .a(n_19316), .b(n_18640), .o(n_20291) );
na02f80 g549790 ( .a(n_19884), .b(n_19253), .o(n_21244) );
no02f80 g549791 ( .a(n_19322), .b(n_19010), .o(n_19011) );
na02f80 g549792 ( .a(n_19547), .b(n_18955), .o(n_20288) );
na02f80 g549793 ( .a(n_19546), .b(n_18953), .o(n_20611) );
na02f80 g549794 ( .a(n_19545), .b(n_18948), .o(n_20608) );
na02f80 g549795 ( .a(n_19544), .b(n_18951), .o(n_20285) );
na02f80 g549796 ( .a(n_20525), .b(n_19794), .o(n_21238) );
na02f80 g549797 ( .a(n_20524), .b(n_19807), .o(n_21241) );
no02f80 g549798 ( .a(n_19891), .b(n_19542), .o(n_19543) );
no02f80 g549799 ( .a(n_18858), .b(n_19542), .o(n_20686) );
na02f80 g549800 ( .a(n_20215), .b(n_19490), .o(n_20937) );
na02f80 g549801 ( .a(n_17809), .b(n_18095), .o(n_19062) );
na02f80 g549802 ( .a(n_17810), .b(n_17495), .o(n_17496) );
na02f80 g549803 ( .a(n_19315), .b(x_in_48_3), .o(n_20277) );
in01f80 g549804 ( .a(n_19540), .o(n_19541) );
no02f80 g549805 ( .a(n_19315), .b(x_in_48_3), .o(n_19540) );
na02f80 g549806 ( .a(n_19883), .b(n_19270), .o(n_20650) );
na02f80 g549807 ( .a(n_19882), .b(n_19242), .o(n_20598) );
in01f80 g549808 ( .a(n_19313), .o(n_19314) );
no02f80 g549809 ( .a(n_19304), .b(x_in_38_8), .o(n_19313) );
na02f80 g549810 ( .a(n_20907), .b(n_20136), .o(n_21597) );
na02f80 g549811 ( .a(n_19539), .b(n_18942), .o(n_20595) );
no02f80 g549812 ( .a(n_19568), .b(n_19311), .o(n_19312) );
in01f80 g549813 ( .a(n_20213), .o(n_20214) );
na02f80 g549814 ( .a(n_19881), .b(n_19226), .o(n_20213) );
na02f80 g549815 ( .a(n_19880), .b(n_19221), .o(n_20591) );
in01f80 g549816 ( .a(n_19008), .o(n_19009) );
no02f80 g549817 ( .a(n_18667), .b(x_in_24_6), .o(n_19008) );
na02f80 g549818 ( .a(n_18667), .b(x_in_24_6), .o(n_19623) );
na02f80 g549819 ( .a(n_19321), .b(n_19006), .o(n_19007) );
na02f80 g549820 ( .a(n_19538), .b(n_18936), .o(n_20268) );
in01f80 g549821 ( .a(n_20522), .o(n_20523) );
na02f80 g549822 ( .a(n_20212), .b(n_19488), .o(n_20522) );
na02f80 g549823 ( .a(n_19304), .b(x_in_38_8), .o(n_19973) );
na02f80 g549824 ( .a(n_19310), .b(x_in_28_8), .o(n_20261) );
in01f80 g549825 ( .a(n_19536), .o(n_19537) );
no02f80 g549826 ( .a(n_19310), .b(x_in_28_8), .o(n_19536) );
in01f80 g549827 ( .a(n_19878), .o(n_19879) );
na02f80 g549828 ( .a(n_19535), .b(n_18933), .o(n_19878) );
na02f80 g549829 ( .a(n_19534), .b(n_18931), .o(n_20583) );
no02f80 g549830 ( .a(n_19876), .b(n_19875), .o(n_19877) );
in01f80 g549831 ( .a(n_20210), .o(n_20211) );
na02f80 g549832 ( .a(n_19874), .b(n_19214), .o(n_20210) );
na02f80 g549833 ( .a(n_20209), .b(n_19507), .o(n_20945) );
na02f80 g549834 ( .a(n_19873), .b(n_19191), .o(n_20641) );
na02f80 g549835 ( .a(n_19533), .b(n_18926), .o(n_20579) );
na02f80 g549836 ( .a(n_20906), .b(n_20147), .o(n_21594) );
na02f80 g549837 ( .a(n_20208), .b(n_19509), .o(n_20948) );
na02f80 g549838 ( .a(n_21195), .b(n_20488), .o(n_21985) );
na02f80 g549839 ( .a(n_20207), .b(n_19479), .o(n_20927) );
na02f80 g549840 ( .a(n_19532), .b(n_18921), .o(n_20569) );
no02f80 g549841 ( .a(n_18096), .b(n_18095), .o(n_18097) );
na02f80 g549842 ( .a(n_20521), .b(n_19777), .o(n_21230) );
na02f80 g549843 ( .a(n_19872), .b(n_19268), .o(n_20647) );
na02f80 g549844 ( .a(n_19871), .b(x_in_44_5), .o(n_20924) );
in01f80 g549845 ( .a(n_20205), .o(n_20206) );
no02f80 g549846 ( .a(n_19871), .b(x_in_44_5), .o(n_20205) );
na02f80 g549847 ( .a(n_20520), .b(n_19801), .o(n_21225) );
in01f80 g549848 ( .a(n_20203), .o(n_20204) );
no02f80 g549849 ( .a(n_19870), .b(x_in_28_7), .o(n_20203) );
na02f80 g549850 ( .a(n_19870), .b(x_in_28_7), .o(n_20923) );
in01f80 g549851 ( .a(n_20201), .o(n_20202) );
na02f80 g549852 ( .a(n_19869), .b(n_19273), .o(n_20201) );
no02f80 g549853 ( .a(n_18676), .b(n_18393), .o(n_18394) );
no02f80 g549854 ( .a(n_20226), .b(n_19867), .o(n_19868) );
no02f80 g549855 ( .a(n_19169), .b(n_19867), .o(n_20986) );
na02f80 g549856 ( .a(n_19336), .b(n_19004), .o(n_19005) );
na02f80 g549857 ( .a(n_19309), .b(n_19529), .o(n_20675) );
no02f80 g549858 ( .a(n_19530), .b(n_19529), .o(n_19531) );
no02f80 g549859 ( .a(n_18672), .b(n_18666), .o(n_19345) );
na02f80 g549860 ( .a(n_18391), .b(n_18666), .o(n_18392) );
na02f80 g549861 ( .a(n_19307), .b(n_19306), .o(n_19308) );
no02f80 g549862 ( .a(n_19310), .b(n_19306), .o(n_20339) );
na02f80 g549863 ( .a(n_20238), .b(n_19865), .o(n_19866) );
no02f80 g549864 ( .a(n_18664), .b(n_18663), .o(n_18665) );
na02f80 g549865 ( .a(n_18390), .b(n_18663), .o(n_20012) );
na02f80 g549866 ( .a(n_19014), .b(n_18661), .o(n_18662) );
na02f80 g549867 ( .a(n_19304), .b(n_19303), .o(n_19305) );
na02f80 g549868 ( .a(n_18582), .b(n_19303), .o(n_20338) );
no02f80 g549869 ( .a(n_19863), .b(n_19862), .o(n_19864) );
no02f80 g549870 ( .a(n_18660), .b(n_18031), .o(n_20005) );
in01f80 g549871 ( .a(n_20997), .o(n_19528) );
oa12f80 g549872 ( .a(n_19228), .b(n_18562), .c(n_17619), .o(n_20997) );
na02f80 g549873 ( .a(n_19290), .b(n_19002), .o(n_19003) );
no02f80 g549874 ( .a(n_18093), .b(n_18092), .o(n_18094) );
no02f80 g549875 ( .a(n_19526), .b(n_19525), .o(n_19527) );
in01f80 g549876 ( .a(n_19524), .o(n_20332) );
na02f80 g549877 ( .a(n_19302), .b(n_19525), .o(n_19524) );
no02f80 g549878 ( .a(n_18660), .b(n_18658), .o(n_18659) );
in01f80 g549879 ( .a(n_20905), .o(n_22010) );
ao12f80 g549880 ( .a(n_17771), .b(n_20515), .c(n_18320), .o(n_20905) );
oa12f80 g549881 ( .a(n_15841), .b(n_18657), .c(n_16494), .o(n_19665) );
oa12f80 g549882 ( .a(n_13669), .b(n_18656), .c(n_14786), .o(n_19664) );
ao12f80 g549883 ( .a(n_15553), .b(n_18091), .c(n_16244), .o(n_19060) );
ao12f80 g549884 ( .a(n_14776), .b(n_18655), .c(n_15342), .o(n_19663) );
ao12f80 g549885 ( .a(n_14754), .b(n_18389), .c(n_15423), .o(n_19385) );
in01f80 g549886 ( .a(n_20200), .o(n_21280) );
oa12f80 g549887 ( .a(n_18565), .b(n_19854), .c(n_17986), .o(n_20200) );
oa12f80 g549888 ( .a(n_12262), .b(n_18388), .c(n_12437), .o(n_19379) );
ao12f80 g549889 ( .a(n_14651), .b(n_18387), .c(n_15406), .o(n_19384) );
ao12f80 g549890 ( .a(n_14739), .b(n_18386), .c(n_15396), .o(n_19383) );
oa12f80 g549891 ( .a(n_14378), .b(n_18385), .c(n_15141), .o(n_19382) );
ao12f80 g549892 ( .a(n_14711), .b(n_18384), .c(n_15384), .o(n_19381) );
ao12f80 g549893 ( .a(n_14685), .b(n_18383), .c(n_15366), .o(n_19380) );
oa12f80 g549894 ( .a(n_13150), .b(n_18654), .c(n_14318), .o(n_19662) );
in01f80 g549895 ( .a(n_19523), .o(n_20669) );
ao12f80 g549896 ( .a(n_12302), .b(n_19292), .c(n_12953), .o(n_19523) );
in01f80 g549897 ( .a(n_20519), .o(n_21613) );
oa12f80 g549898 ( .a(n_19139), .b(n_20199), .c(n_18478), .o(n_20519) );
ao12f80 g549899 ( .a(n_16098), .b(n_19301), .c(n_16679), .o(n_20331) );
in01f80 g549900 ( .a(n_19522), .o(n_20668) );
ao12f80 g549901 ( .a(n_11016), .b(n_19289), .c(n_12120), .o(n_19522) );
in01f80 g549902 ( .a(n_20198), .o(n_21276) );
oa12f80 g549903 ( .a(n_18570), .b(n_19848), .c(n_17977), .o(n_20198) );
in01f80 g549904 ( .a(n_20197), .o(n_21273) );
oa12f80 g549905 ( .a(n_19209), .b(n_18821), .c(n_18557), .o(n_20197) );
ao12f80 g549906 ( .a(n_15501), .b(n_19300), .c(n_16247), .o(n_20330) );
oa12f80 g549907 ( .a(n_11421), .b(n_18382), .c(n_12430), .o(n_19378) );
oa12f80 g549908 ( .a(n_14674), .b(n_18381), .c(n_15348), .o(n_19377) );
oa12f80 g549909 ( .a(n_14699), .b(n_18653), .c(n_15371), .o(n_19661) );
ao12f80 g549910 ( .a(n_11497), .b(n_18090), .c(n_12485), .o(n_19061) );
oa12f80 g549911 ( .a(n_14345), .b(n_18380), .c(n_15130), .o(n_19376) );
oa12f80 g549912 ( .a(n_15761), .b(n_19001), .c(n_16491), .o(n_20004) );
ao12f80 g549913 ( .a(n_8308), .b(n_18652), .c(n_8943), .o(n_19659) );
oa12f80 g549914 ( .a(n_15060), .b(n_19299), .c(n_14661), .o(n_19936) );
oa12f80 g549915 ( .a(n_14303), .b(n_18651), .c(n_15112), .o(n_19660) );
ao12f80 g549916 ( .a(n_13201), .b(n_18379), .c(n_14412), .o(n_19375) );
oa12f80 g549917 ( .a(n_13181), .b(n_19298), .c(n_14368), .o(n_20329) );
ao12f80 g549918 ( .a(n_14442), .b(n_18378), .c(n_15115), .o(n_19374) );
ao12f80 g549919 ( .a(n_14415), .b(n_18650), .c(n_15154), .o(n_19658) );
ao12f80 g549920 ( .a(n_10655), .b(n_18089), .c(n_11791), .o(n_19059) );
oa12f80 g549921 ( .a(n_13161), .b(n_19000), .c(n_14326), .o(n_20003) );
oa12f80 g549922 ( .a(n_14255), .b(n_18377), .c(n_15099), .o(n_19373) );
oa12f80 g549923 ( .a(n_14248), .b(n_18376), .c(n_15094), .o(n_19372) );
oa12f80 g549924 ( .a(n_11502), .b(n_18649), .c(n_12487), .o(n_19657) );
oa12f80 g549925 ( .a(n_15520), .b(n_18375), .c(n_16257), .o(n_19371) );
oa12f80 g549926 ( .a(n_13879), .b(n_18374), .c(n_14925), .o(n_19370) );
ao12f80 g549927 ( .a(n_14672), .b(n_18373), .c(n_15354), .o(n_19369) );
oa12f80 g549928 ( .a(n_10769), .b(n_18372), .c(n_11803), .o(n_19368) );
ao12f80 g549929 ( .a(n_8823), .b(n_18371), .c(n_10342), .o(n_19367) );
ao12f80 g549930 ( .a(n_18889), .b(n_18888), .c(n_18887), .o(n_19521) );
ao12f80 g549931 ( .a(n_20486), .b(n_20485), .c(n_20484), .o(n_21194) );
ao12f80 g549932 ( .a(n_19825), .b(n_19824), .c(n_19823), .o(n_20518) );
ao12f80 g549933 ( .a(n_19495), .b(n_19494), .c(n_19493), .o(n_20196) );
oa12f80 g549934 ( .a(n_18883), .b(n_18882), .c(n_18881), .o(n_20313) );
ao12f80 g549935 ( .a(n_19476), .b(n_19835), .c(n_19475), .o(n_20195) );
oa12f80 g549936 ( .a(n_18893), .b(n_18892), .c(n_18894), .o(n_20256) );
ao12f80 g549937 ( .a(n_18981), .b(n_18980), .c(n_18979), .o(n_19520) );
ao12f80 g549938 ( .a(n_19822), .b(n_19821), .c(n_19820), .o(n_20517) );
ao22s80 g549939 ( .a(n_18572), .b(n_20515), .c(n_18571), .d(n_19413), .o(n_20516) );
oa12f80 g549940 ( .a(n_18344), .b(n_18343), .c(n_18596), .o(n_19649) );
ao12f80 g549941 ( .a(n_18977), .b(n_19282), .c(n_18976), .o(n_19519) );
ao12f80 g549942 ( .a(n_20174), .b(n_20173), .c(n_20172), .o(n_20904) );
oa12f80 g549943 ( .a(n_18868), .b(n_18918), .c(n_19189), .o(n_20254) );
oa12f80 g549944 ( .a(n_18342), .b(n_18341), .c(n_18611), .o(n_19612) );
ao12f80 g549945 ( .a(n_18607), .b(n_18608), .c(n_18606), .o(n_19297) );
ao12f80 g549946 ( .a(n_20171), .b(n_20170), .c(n_20169), .o(n_20903) );
oa12f80 g549947 ( .a(n_18340), .b(n_18609), .c(n_18339), .o(n_19648) );
ao12f80 g549948 ( .a(n_19819), .b(n_19818), .c(n_19817), .o(n_20514) );
oa12f80 g549949 ( .a(n_18338), .b(n_18597), .c(n_18337), .o(n_19647) );
in01f80 g549950 ( .a(FE_OFN1061_n_19587), .o(n_19296) );
oa12f80 g549951 ( .a(n_18365), .b(n_18656), .c(n_18364), .o(n_19587) );
ao12f80 g549952 ( .a(n_19789), .b(n_19788), .c(n_19787), .o(n_20513) );
oa12f80 g549953 ( .a(n_18878), .b(n_18877), .c(n_18876), .o(n_20281) );
in01f80 g549954 ( .a(n_19595), .o(n_18999) );
oa12f80 g549955 ( .a(n_18086), .b(n_18389), .c(n_18085), .o(n_19595) );
ao12f80 g549956 ( .a(n_19262), .b(n_19261), .c(n_19260), .o(n_19861) );
ao12f80 g549957 ( .a(n_19482), .b(n_19481), .c(n_19480), .o(n_20194) );
ao12f80 g549958 ( .a(n_19816), .b(n_19815), .c(n_19814), .o(n_20512) );
ao12f80 g549959 ( .a(n_19782), .b(n_19781), .c(n_19780), .o(n_20511) );
oa12f80 g549960 ( .a(n_18601), .b(n_18644), .c(n_18862), .o(n_19974) );
ao12f80 g549961 ( .a(n_20134), .b(n_20133), .c(n_20132), .o(n_20902) );
oa12f80 g549962 ( .a(n_18909), .b(n_18908), .c(n_18910), .o(n_20303) );
ao12f80 g549963 ( .a(n_20155), .b(n_20154), .c(n_20153), .o(n_20901) );
oa12f80 g549964 ( .a(n_18886), .b(n_18885), .c(n_18884), .o(n_20314) );
in01f80 g549965 ( .a(n_19337), .o(n_19645) );
ao12f80 g549966 ( .a(n_18064), .b(n_18378), .c(n_18063), .o(n_19337) );
oa12f80 g549967 ( .a(n_18913), .b(n_18912), .c(n_18911), .o(n_20302) );
in01f80 g549968 ( .a(n_19903), .o(n_19361) );
ao12f80 g549969 ( .a(n_17808), .b(n_18091), .c(n_17807), .o(n_19903) );
in01f80 g549970 ( .a(n_19642), .o(n_19295) );
oa12f80 g549971 ( .a(n_18362), .b(n_18655), .c(n_18361), .o(n_19642) );
ao12f80 g549972 ( .a(n_20164), .b(n_20163), .c(n_20162), .o(n_20900) );
oa12f80 g549973 ( .a(n_18903), .b(n_18902), .c(n_18904), .o(n_20270) );
oa12f80 g549974 ( .a(n_18906), .b(n_18905), .c(n_18907), .o(n_20301) );
oa22f80 g549975 ( .a(n_18087), .b(FE_OFN249_n_4162), .c(n_617), .d(FE_OFN1111_rst), .o(n_18088) );
ao12f80 g549976 ( .a(n_19259), .b(n_19258), .c(n_19257), .o(n_19860) );
in01f80 g549977 ( .a(n_19901), .o(n_19981) );
ao12f80 g549978 ( .a(n_18367), .b(n_18657), .c(n_18366), .o(n_19901) );
ao12f80 g549979 ( .a(n_20158), .b(n_20157), .c(n_20156), .o(n_20899) );
oa12f80 g549980 ( .a(n_18900), .b(n_18899), .c(n_18901), .o(n_20300) );
ao12f80 g549981 ( .a(n_20161), .b(n_20160), .c(n_20159), .o(n_20898) );
oa12f80 g549982 ( .a(n_18897), .b(n_18896), .c(n_18898), .o(n_20299) );
ao12f80 g549983 ( .a(n_19202), .b(n_19201), .c(n_19200), .o(n_19859) );
ao12f80 g549984 ( .a(n_20168), .b(n_20167), .c(n_20166), .o(n_20897) );
in01f80 g549985 ( .a(n_19597), .o(n_18998) );
oa12f80 g549986 ( .a(n_18082), .b(n_18387), .c(n_18081), .o(n_19597) );
in01f80 g549987 ( .a(n_19335), .o(n_18997) );
oa12f80 g549988 ( .a(n_18066), .b(n_18379), .c(n_18065), .o(n_19335) );
ao12f80 g549989 ( .a(n_19256), .b(n_19255), .c(n_19254), .o(n_19858) );
in01f80 g549990 ( .a(n_19573), .o(n_19968) );
ao12f80 g549991 ( .a(n_18351), .b(n_18650), .c(n_18350), .o(n_19573) );
in01f80 g549992 ( .a(n_19599), .o(n_18996) );
oa12f80 g549993 ( .a(n_18080), .b(n_18386), .c(n_18079), .o(n_19599) );
ao12f80 g549994 ( .a(n_19251), .b(n_19250), .c(n_19249), .o(n_19857) );
in01f80 g549995 ( .a(n_19914), .o(n_19634) );
ao12f80 g549996 ( .a(n_18078), .b(n_18385), .c(n_18077), .o(n_19914) );
ao12f80 g549997 ( .a(n_19498), .b(n_19497), .c(n_19496), .o(n_20193) );
oa12f80 g549998 ( .a(n_18336), .b(n_18335), .c(n_18605), .o(n_19646) );
in01f80 g549999 ( .a(FE_OFN751_n_20252), .o(n_20562) );
ao12f80 g550000 ( .a(n_18915), .b(n_19298), .c(n_18914), .o(n_20252) );
ao12f80 g550001 ( .a(n_19797), .b(n_19796), .c(n_19795), .o(n_20510) );
ao12f80 g550002 ( .a(n_19248), .b(n_19247), .c(n_19246), .o(n_19856) );
in01f80 g550003 ( .a(n_19592), .o(n_18995) );
oa12f80 g550004 ( .a(n_18076), .b(n_18384), .c(n_18075), .o(n_19592) );
in01f80 g550005 ( .a(n_19564), .o(n_19631) );
ao12f80 g550006 ( .a(n_18068), .b(n_18380), .c(n_18067), .o(n_19564) );
ao22s80 g550007 ( .a(n_18842), .b(n_19854), .c(n_18841), .d(n_18820), .o(n_19855) );
ao12f80 g550008 ( .a(n_19245), .b(n_19244), .c(n_19243), .o(n_19853) );
in01f80 g550009 ( .a(n_19630), .o(n_19294) );
oa12f80 g550010 ( .a(n_18357), .b(n_18653), .c(n_18356), .o(n_19630) );
in01f80 g550011 ( .a(n_19607), .o(n_18994) );
oa12f80 g550012 ( .a(n_18074), .b(n_18383), .c(n_18073), .o(n_19607) );
ao12f80 g550013 ( .a(n_19240), .b(n_19239), .c(n_19238), .o(n_19852) );
in01f80 g550014 ( .a(n_19639), .o(n_19985) );
ao12f80 g550015 ( .a(n_18349), .b(n_18649), .c(n_18348), .o(n_19639) );
ao12f80 g550016 ( .a(n_18946), .b(n_18945), .c(n_18944), .o(n_19518) );
oa12f80 g550017 ( .a(n_19187), .b(n_19186), .c(n_19188), .o(n_20606) );
ao12f80 g550018 ( .a(n_18333), .b(n_18332), .c(n_18331), .o(n_18993) );
ao12f80 g550019 ( .a(n_19470), .b(n_19469), .c(n_19468), .o(n_20192) );
oa12f80 g550020 ( .a(n_18874), .b(n_18873), .c(n_18875), .o(n_20283) );
ao12f80 g550021 ( .a(n_19792), .b(n_19791), .c(n_19790), .o(n_20509) );
in01f80 g550022 ( .a(n_19583), .o(n_19627) );
ao12f80 g550023 ( .a(n_18054), .b(n_18373), .c(n_18053), .o(n_19583) );
in01f80 g550024 ( .a(n_19912), .o(n_20262) );
ao12f80 g550025 ( .a(n_18613), .b(n_19000), .c(n_18612), .o(n_19912) );
oa12f80 g550026 ( .a(n_18870), .b(n_18871), .c(n_18869), .o(n_20282) );
ao12f80 g550027 ( .a(n_20152), .b(n_20151), .c(n_20150), .o(n_20896) );
ao12f80 g550028 ( .a(n_19234), .b(n_19233), .c(n_19232), .o(n_19851) );
ao12f80 g550029 ( .a(n_18604), .b(n_18603), .c(n_18602), .o(n_19293) );
in01f80 g550030 ( .a(FE_OFN899_n_19332), .o(n_19571) );
ao12f80 g550031 ( .a(n_18049), .b(n_18371), .c(n_18048), .o(n_19332) );
in01f80 g550032 ( .a(n_19989), .o(n_19517) );
oa22f80 g550033 ( .a(n_19292), .b(n_13504), .c(n_18300), .d(n_13505), .o(n_19989) );
oa12f80 g550034 ( .a(n_18615), .b(n_18614), .c(n_18895), .o(n_19959) );
ao12f80 g550036 ( .a(n_18360), .b(n_18654), .c(n_18359), .o(n_19575) );
in01f80 g550037 ( .a(n_20660), .o(n_20593) );
ao12f80 g550038 ( .a(n_18917), .b(n_19299), .c(n_18916), .o(n_20660) );
ao12f80 g550039 ( .a(n_19224), .b(n_19223), .c(n_19222), .o(n_19850) );
ao22s80 g550040 ( .a(n_19422), .b(n_20199), .c(n_19421), .d(n_19128), .o(n_20508) );
in01f80 g550041 ( .a(n_19908), .o(n_19952) );
ao12f80 g550042 ( .a(n_18353), .b(n_18651), .c(n_18352), .o(n_19908) );
oa12f80 g550043 ( .a(n_18600), .b(n_18599), .c(n_18867), .o(n_19958) );
in01f80 g550044 ( .a(n_20248), .o(n_19624) );
ao12f80 g550045 ( .a(n_18058), .b(n_18375), .c(n_18057), .o(n_20248) );
ao12f80 g550046 ( .a(n_17802), .b(n_18087), .c(n_17801), .o(n_18370) );
ao12f80 g550047 ( .a(n_19467), .b(n_19466), .c(n_19465), .o(n_20191) );
in01f80 g550048 ( .a(FE_OFN724_n_19019), .o(n_18648) );
oa12f80 g550049 ( .a(n_17806), .b(n_18090), .c(n_17805), .o(n_19019) );
na03f80 g550050 ( .a(n_11830), .b(n_19290), .c(n_12340), .o(n_19291) );
in01f80 g550051 ( .a(n_19577), .o(n_19611) );
ao12f80 g550052 ( .a(n_18072), .b(n_18381), .c(n_18071), .o(n_19577) );
ao12f80 g550053 ( .a(n_19786), .b(n_19785), .c(n_19784), .o(n_20507) );
ao12f80 g550054 ( .a(n_20139), .b(n_20138), .c(n_20137), .o(n_20895) );
in01f80 g550055 ( .a(n_19905), .o(n_20298) );
ao22s80 g550056 ( .a(n_18298), .b(n_12542), .c(n_19289), .d(n_12541), .o(n_19905) );
oa12f80 g550057 ( .a(n_18594), .b(n_18595), .c(n_18593), .o(n_19953) );
in01f80 g550058 ( .a(n_19323), .o(n_19622) );
ao12f80 g550059 ( .a(n_18062), .b(n_18377), .c(n_18061), .o(n_19323) );
ao12f80 g550060 ( .a(n_18592), .b(n_18591), .c(n_18590), .o(n_19288) );
in01f80 g550061 ( .a(n_19330), .o(n_18992) );
oa12f80 g550062 ( .a(n_18052), .b(n_18372), .c(n_18051), .o(n_19330) );
ao22s80 g550063 ( .a(n_18845), .b(n_19848), .c(n_18844), .d(n_18818), .o(n_19849) );
ao12f80 g550064 ( .a(n_19212), .b(n_19211), .c(n_19210), .o(n_19847) );
in01f80 g550065 ( .a(n_20555), .o(n_20581) );
ao12f80 g550066 ( .a(n_18928), .b(n_19301), .c(n_18927), .o(n_20555) );
ao12f80 g550067 ( .a(n_18347), .b(n_18346), .c(n_18345), .o(n_18991) );
in01f80 g550068 ( .a(n_18647), .o(n_19654) );
oa12f80 g550069 ( .a(n_17804), .b(n_18089), .c(n_17803), .o(n_18647) );
in01f80 g550070 ( .a(n_19333), .o(n_19620) );
ao12f80 g550071 ( .a(n_18060), .b(n_18376), .c(n_18059), .o(n_19333) );
in01f80 g550072 ( .a(n_19589), .o(n_19928) );
ao12f80 g550073 ( .a(n_18355), .b(n_18652), .c(n_18354), .o(n_19589) );
in01f80 g550074 ( .a(n_20556), .o(n_20587) );
ao12f80 g550075 ( .a(n_18924), .b(n_19300), .c(n_18923), .o(n_20556) );
oa12f80 g550076 ( .a(n_19461), .b(n_19773), .c(n_19460), .o(n_20931) );
ao12f80 g550077 ( .a(n_19231), .b(n_19230), .c(n_19229), .o(n_19846) );
ao12f80 g550078 ( .a(n_19208), .b(n_19207), .c(n_19206), .o(n_19845) );
ao12f80 g550079 ( .a(n_19217), .b(n_19216), .c(n_19215), .o(n_19844) );
ao12f80 g550080 ( .a(n_18624), .b(n_18988), .c(n_18623), .o(n_19287) );
in01f80 g550081 ( .a(n_19354), .o(n_19618) );
ao12f80 g550082 ( .a(n_18070), .b(n_18388), .c(n_18069), .o(n_19354) );
ao12f80 g550083 ( .a(n_20483), .b(n_20482), .c(n_20481), .o(n_21193) );
oa12f80 g550084 ( .a(n_19180), .b(n_19271), .c(n_19458), .o(n_20575) );
in01f80 g550085 ( .a(n_19327), .o(n_19616) );
ao12f80 g550086 ( .a(n_18056), .b(n_18374), .c(n_18055), .o(n_19327) );
ao12f80 g550087 ( .a(n_18621), .b(n_18982), .c(n_18620), .o(n_19286) );
ao12f80 g550088 ( .a(n_20881), .b(n_20880), .c(n_20879), .o(n_21571) );
oa12f80 g550089 ( .a(n_18864), .b(n_18865), .c(n_18863), .o(n_20257) );
ao12f80 g550090 ( .a(n_18587), .b(n_18586), .c(n_18585), .o(n_19285) );
ao12f80 g550091 ( .a(n_19464), .b(n_19463), .c(n_19462), .o(n_20190) );
ao12f80 g550092 ( .a(n_19199), .b(n_19198), .c(n_19197), .o(n_19843) );
ao12f80 g550093 ( .a(n_20142), .b(n_20141), .c(n_20140), .o(n_20894) );
in01f80 g550094 ( .a(n_20925), .o(n_20506) );
oa12f80 g550095 ( .a(n_19472), .b(n_19474), .c(n_19471), .o(n_20925) );
ao12f80 g550096 ( .a(n_19196), .b(n_19195), .c(n_19194), .o(n_19842) );
ao12f80 g550097 ( .a(n_18891), .b(n_19278), .c(n_18890), .o(n_19516) );
in01f80 g550098 ( .a(FE_OFN630_n_19358), .o(n_19614) );
ao12f80 g550099 ( .a(n_18084), .b(n_18382), .c(n_18083), .o(n_19358) );
in01f80 g550100 ( .a(n_19925), .o(n_20255) );
ao12f80 g550101 ( .a(n_18617), .b(n_19001), .c(n_18616), .o(n_19925) );
oa22f80 g550102 ( .a(FE_OFN1057_n_18817), .b(n_23291), .c(n_1075), .d(FE_OFN324_n_4860), .o(n_19841) );
oa22f80 g550103 ( .a(n_19408), .b(n_22960), .c(n_352), .d(FE_OFN89_n_27449), .o(n_20505) );
oa22f80 g550104 ( .a(n_19736), .b(FE_OFN225_n_21642), .c(n_1555), .d(FE_OFN134_n_27449), .o(n_20893) );
oa22f80 g550105 ( .a(n_19412), .b(n_22960), .c(n_953), .d(FE_OFN122_n_27449), .o(n_20504) );
oa22f80 g550106 ( .a(n_19127), .b(FE_OFN313_n_3069), .c(n_27), .d(FE_OFN139_n_27449), .o(n_20189) );
oa22f80 g550107 ( .a(n_18816), .b(FE_OFN264_n_4280), .c(n_1699), .d(FE_OFN1110_rst), .o(n_19840) );
oa22f80 g550108 ( .a(n_19411), .b(FE_OFN417_n_28303), .c(n_869), .d(FE_OFN285_n_29266), .o(n_20503) );
oa22f80 g550109 ( .a(n_19126), .b(FE_OFN406_n_28303), .c(n_974), .d(FE_OFN21_n_27452), .o(n_20188) );
oa22f80 g550110 ( .a(n_18537), .b(FE_OFN256_n_4280), .c(n_887), .d(FE_OFN80_n_27012), .o(n_19515) );
oa22f80 g550111 ( .a(n_19735), .b(FE_OFN254_n_4280), .c(n_1073), .d(FE_OFN131_n_27449), .o(n_20892) );
oa22f80 g550112 ( .a(n_19734), .b(FE_OFN411_n_28303), .c(n_817), .d(FE_OFN129_n_27449), .o(n_20891) );
oa22f80 g550113 ( .a(n_19410), .b(FE_OFN259_n_4280), .c(n_1113), .d(FE_OFN1119_rst), .o(n_20502) );
oa22f80 g550114 ( .a(FE_OFN1059_n_18610), .b(FE_OFN405_n_28303), .c(n_262), .d(n_29264), .o(n_18990) );
oa22f80 g550115 ( .a(n_19409), .b(FE_OFN400_n_28303), .c(n_1474), .d(n_27449), .o(n_20501) );
oa22f80 g550116 ( .a(n_18815), .b(FE_OFN234_n_4162), .c(n_1584), .d(FE_OFN122_n_27449), .o(n_19839) );
oa22f80 g550117 ( .a(n_19124), .b(FE_OFN268_n_4280), .c(n_1205), .d(FE_OFN93_n_27449), .o(n_20187) );
oa22f80 g550118 ( .a(n_19120), .b(n_21076), .c(n_1218), .d(n_27449), .o(n_20186) );
oa22f80 g550119 ( .a(n_18050), .b(FE_OFN267_n_4280), .c(n_462), .d(FE_OFN92_n_27449), .o(n_18369) );
oa22f80 g550120 ( .a(n_19123), .b(n_22019), .c(n_718), .d(n_27449), .o(n_20185) );
oa22f80 g550121 ( .a(n_19407), .b(FE_OFN253_n_4280), .c(n_764), .d(FE_OFN136_n_27449), .o(n_20500) );
oa22f80 g550122 ( .a(n_19406), .b(FE_OFN257_n_4280), .c(n_1407), .d(FE_OFN349_n_4860), .o(n_20499) );
oa22f80 g550123 ( .a(n_19733), .b(FE_OFN239_n_4162), .c(n_856), .d(FE_OFN136_n_27449), .o(n_20890) );
oa22f80 g550124 ( .a(n_19405), .b(FE_OFN260_n_4280), .c(n_394), .d(FE_OFN125_n_27449), .o(n_20498) );
oa22f80 g550125 ( .a(n_19404), .b(FE_OFN251_n_4162), .c(n_367), .d(FE_OFN98_n_27449), .o(n_20497) );
oa22f80 g550126 ( .a(n_19403), .b(n_22615), .c(n_1354), .d(FE_OFN287_n_29266), .o(n_20496) );
oa22f80 g550127 ( .a(n_19402), .b(n_22615), .c(n_1855), .d(FE_OFN324_n_4860), .o(n_20495) );
oa22f80 g550128 ( .a(n_18293), .b(FE_OFN235_n_4162), .c(n_1643), .d(FE_OFN287_n_29266), .o(n_19284) );
oa22f80 g550129 ( .a(n_19732), .b(FE_OFN257_n_4280), .c(n_383), .d(FE_OFN95_n_27449), .o(n_20889) );
oa22f80 g550130 ( .a(FE_OFN444_n_19118), .b(n_21076), .c(n_1264), .d(FE_OFN96_n_27449), .o(n_20184) );
oa22f80 g550131 ( .a(n_18329), .b(n_4162), .c(n_469), .d(FE_OFN115_n_27449), .o(n_18646) );
oa22f80 g550132 ( .a(n_18807), .b(n_4162), .c(n_696), .d(FE_OFN353_n_4860), .o(n_19838) );
oa22f80 g550133 ( .a(n_18328), .b(FE_OFN239_n_4162), .c(n_28), .d(FE_OFN74_n_27012), .o(n_18645) );
oa22f80 g550134 ( .a(n_18988), .b(n_26454), .c(n_1298), .d(FE_OFN99_n_27449), .o(n_18989) );
oa22f80 g550135 ( .a(n_19401), .b(FE_OFN236_n_4162), .c(n_1290), .d(FE_OFN99_n_27449), .o(n_20494) );
oa22f80 g550136 ( .a(n_19731), .b(n_26454), .c(n_1109), .d(FE_OFN72_n_27012), .o(n_20888) );
oa22f80 g550137 ( .a(n_19730), .b(FE_OFN264_n_4280), .c(n_1358), .d(FE_OFN98_n_27449), .o(n_20887) );
oa22f80 g550138 ( .a(n_18813), .b(FE_OFN239_n_4162), .c(n_1252), .d(FE_OFN130_n_27449), .o(n_19837) );
oa22f80 g550139 ( .a(n_19835), .b(FE_OFN254_n_4280), .c(n_1941), .d(FE_OFN139_n_27449), .o(n_19836) );
oa22f80 g550140 ( .a(n_19122), .b(FE_OFN417_n_28303), .c(n_148), .d(FE_OFN139_n_27449), .o(n_20183) );
oa22f80 g550141 ( .a(n_19121), .b(FE_OFN413_n_28303), .c(n_1473), .d(FE_OFN136_n_27449), .o(n_20182) );
oa22f80 g550142 ( .a(n_19729), .b(FE_OFN235_n_4162), .c(n_43), .d(FE_OFN1181_rst), .o(n_20886) );
oa22f80 g550143 ( .a(n_19728), .b(FE_OFN405_n_28303), .c(n_801), .d(FE_OFN324_n_4860), .o(n_20885) );
oa22f80 g550144 ( .a(n_19282), .b(FE_OFN416_n_28303), .c(n_1904), .d(FE_OFN1174_n_4860), .o(n_19283) );
oa22f80 g550145 ( .a(n_18811), .b(FE_OFN417_n_28303), .c(n_420), .d(FE_OFN80_n_27012), .o(n_19834) );
oa22f80 g550146 ( .a(n_18810), .b(FE_OFN149_n_25677), .c(n_294), .d(FE_OFN1124_rst), .o(n_19833) );
oa22f80 g550147 ( .a(n_18026), .b(FE_OFN149_n_25677), .c(n_234), .d(FE_OFN77_n_27012), .o(n_18987) );
oa22f80 g550148 ( .a(FE_OFN580_n_19119), .b(n_23291), .c(n_198), .d(FE_OFN68_n_27012), .o(n_20181) );
oa22f80 g550149 ( .a(n_19727), .b(FE_OFN265_n_4280), .c(n_92), .d(FE_OFN134_n_27449), .o(n_20883) );
oa22f80 g550150 ( .a(n_18809), .b(n_28771), .c(n_1472), .d(FE_OFN11_n_29204), .o(n_19832) );
oa22f80 g550151 ( .a(FE_OFN889_n_18291), .b(n_23813), .c(n_1626), .d(FE_OFN1115_rst), .o(n_19281) );
oa22f80 g550152 ( .a(n_18290), .b(FE_OFN221_n_23315), .c(n_1613), .d(FE_OFN116_n_27449), .o(n_19280) );
oa22f80 g550153 ( .a(n_18536), .b(FE_OFN411_n_28303), .c(n_962), .d(FE_OFN335_n_4860), .o(n_19514) );
oa22f80 g550154 ( .a(n_19726), .b(FE_OFN406_n_28303), .c(n_523), .d(FE_OFN76_n_27012), .o(n_20882) );
oa22f80 g550155 ( .a(n_19117), .b(FE_OFN312_n_3069), .c(n_954), .d(FE_OFN65_n_27012), .o(n_20180) );
oa22f80 g550156 ( .a(n_18047), .b(n_23315), .c(n_590), .d(FE_OFN77_n_27012), .o(n_18368) );
oa22f80 g550157 ( .a(n_18808), .b(FE_OFN297_n_3069), .c(n_1611), .d(FE_OFN358_n_4860), .o(n_19831) );
oa22f80 g550158 ( .a(n_19473), .b(FE_OFN198_n_29637), .c(n_359), .d(FE_OFN124_n_27449), .o(n_19830) );
oa22f80 g550159 ( .a(n_18535), .b(FE_OFN198_n_29637), .c(n_827), .d(FE_OFN124_n_27449), .o(n_19513) );
oa22f80 g550160 ( .a(n_18021), .b(FE_OFN308_n_3069), .c(n_1314), .d(n_29264), .o(n_18986) );
oa22f80 g550161 ( .a(n_19116), .b(FE_OFN269_n_4280), .c(n_424), .d(FE_OFN353_n_4860), .o(n_20179) );
oa22f80 g550162 ( .a(n_18806), .b(FE_OFN259_n_4280), .c(n_618), .d(FE_OFN1119_rst), .o(n_19829) );
oa22f80 g550163 ( .a(n_18024), .b(FE_OFN297_n_3069), .c(n_1659), .d(FE_OFN352_n_4860), .o(n_18985) );
oa22f80 g550164 ( .a(n_18814), .b(FE_OFN312_n_3069), .c(n_1185), .d(FE_OFN124_n_27449), .o(n_19828) );
oa22f80 g550165 ( .a(n_18020), .b(FE_OFN156_n_28014), .c(n_454), .d(FE_OFN330_n_4860), .o(n_18984) );
oa22f80 g550166 ( .a(n_19278), .b(n_28608), .c(n_1742), .d(FE_OFN122_n_27449), .o(n_19279) );
oa22f80 g550167 ( .a(n_18804), .b(FE_OFN199_n_29637), .c(n_1713), .d(n_28607), .o(n_19827) );
oa22f80 g550168 ( .a(n_18288), .b(FE_OFN198_n_29637), .c(n_940), .d(FE_OFN99_n_27449), .o(n_19277) );
oa22f80 g550169 ( .a(n_18287), .b(FE_OFN256_n_4280), .c(n_973), .d(n_27452), .o(n_19276) );
oa22f80 g550170 ( .a(n_18803), .b(FE_OFN295_n_3069), .c(n_986), .d(FE_OFN130_n_27449), .o(n_19826) );
oa22f80 g550171 ( .a(n_18286), .b(FE_OFN259_n_4280), .c(n_1712), .d(FE_OFN135_n_27449), .o(n_19275) );
oa22f80 g550172 ( .a(n_19115), .b(FE_OFN293_n_3069), .c(n_184), .d(FE_OFN105_n_27449), .o(n_20178) );
oa22f80 g550173 ( .a(n_19400), .b(FE_OFN309_n_3069), .c(n_1089), .d(FE_OFN134_n_27449), .o(n_20493) );
oa22f80 g550174 ( .a(n_19114), .b(FE_OFN268_n_4280), .c(n_594), .d(FE_OFN98_n_27449), .o(n_20177) );
oa22f80 g550175 ( .a(n_18534), .b(FE_OFN311_n_3069), .c(n_1784), .d(FE_OFN336_n_4860), .o(n_19512) );
oa22f80 g550176 ( .a(n_18982), .b(n_23813), .c(n_1556), .d(FE_OFN102_n_27449), .o(n_18983) );
oa22f80 g550177 ( .a(n_19113), .b(FE_OFN402_n_28303), .c(n_1934), .d(FE_OFN134_n_27449), .o(n_20176) );
na02f80 g550230 ( .a(n_19274), .b(x_in_2_4), .o(n_20221) );
in01f80 g550231 ( .a(n_19510), .o(n_19511) );
no02f80 g550232 ( .a(n_19274), .b(x_in_2_4), .o(n_19510) );
no02f80 g550233 ( .a(n_19824), .b(n_19823), .o(n_19825) );
no02f80 g550234 ( .a(n_18980), .b(n_18979), .o(n_18981) );
in01f80 g550235 ( .a(n_19508), .o(n_19509) );
no02f80 g550236 ( .a(n_19266), .b(x_in_34_4), .o(n_19508) );
in01f80 g550237 ( .a(n_19272), .o(n_19273) );
no02f80 g550238 ( .a(n_18961), .b(x_in_56_6), .o(n_19272) );
no02f80 g550239 ( .a(n_19821), .b(n_19820), .o(n_19822) );
in01f80 g550240 ( .a(n_20491), .o(n_20492) );
na02f80 g550241 ( .a(n_20175), .b(n_19418), .o(n_20491) );
na02f80 g550242 ( .a(n_19271), .b(x_in_20_4), .o(n_20220) );
na02f80 g550243 ( .a(n_18978), .b(x_in_18_4), .o(n_19883) );
in01f80 g550244 ( .a(n_19269), .o(n_19270) );
no02f80 g550245 ( .a(n_18978), .b(x_in_18_4), .o(n_19269) );
no02f80 g550246 ( .a(n_19282), .b(n_18976), .o(n_18977) );
no02f80 g550247 ( .a(n_20173), .b(n_20172), .o(n_20174) );
na02f80 g550248 ( .a(n_18975), .b(x_in_50_4), .o(n_19872) );
in01f80 g550249 ( .a(n_19267), .o(n_19268) );
no02f80 g550250 ( .a(n_18975), .b(x_in_50_4), .o(n_19267) );
no02f80 g550251 ( .a(n_18657), .b(n_18366), .o(n_18367) );
na02f80 g550252 ( .a(n_18644), .b(x_in_6_4), .o(n_19554) );
in01f80 g550253 ( .a(n_18973), .o(n_18974) );
no02f80 g550254 ( .a(n_18644), .b(x_in_6_4), .o(n_18973) );
no02f80 g550255 ( .a(n_20170), .b(n_20169), .o(n_20171) );
in01f80 g550256 ( .a(n_18971), .o(n_18972) );
no02f80 g550257 ( .a(n_18626), .b(x_in_10_4), .o(n_18971) );
na02f80 g550258 ( .a(n_19499), .b(x_in_62_4), .o(n_20520) );
no02f80 g550259 ( .a(n_19818), .b(n_19817), .o(n_19819) );
na02f80 g550260 ( .a(n_18643), .b(x_in_42_4), .o(n_19555) );
in01f80 g550261 ( .a(n_18969), .o(n_18970) );
no02f80 g550262 ( .a(n_18643), .b(x_in_42_4), .o(n_18969) );
na02f80 g550263 ( .a(n_19266), .b(x_in_34_4), .o(n_20208) );
na02f80 g550264 ( .a(n_18389), .b(n_18085), .o(n_18086) );
na02f80 g550265 ( .a(n_18656), .b(n_18364), .o(n_18365) );
in01f80 g550266 ( .a(n_19506), .o(n_19507) );
no02f80 g550267 ( .a(n_19227), .b(x_in_26_4), .o(n_19506) );
no02f80 g550268 ( .a(n_19815), .b(n_19814), .o(n_19816) );
na02f80 g550269 ( .a(n_18642), .b(x_in_58_4), .o(n_19553) );
in01f80 g550270 ( .a(n_18967), .o(n_18968) );
no02f80 g550271 ( .a(n_18642), .b(x_in_58_4), .o(n_18967) );
na02f80 g550272 ( .a(n_19505), .b(x_in_6_3), .o(n_20526) );
in01f80 g550273 ( .a(n_19812), .o(n_19813) );
no02f80 g550274 ( .a(n_19505), .b(x_in_6_3), .o(n_19812) );
no02f80 g550275 ( .a(n_20167), .b(n_20166), .o(n_20168) );
in01f80 g550276 ( .a(n_19503), .o(n_19504) );
na02f80 g550277 ( .a(n_19265), .b(n_18568), .o(n_19503) );
in01f80 g550278 ( .a(n_20489), .o(n_20490) );
na02f80 g550279 ( .a(n_20165), .b(n_19428), .o(n_20489) );
na02f80 g550280 ( .a(n_19502), .b(x_in_22_4), .o(n_20530) );
in01f80 g550281 ( .a(n_19810), .o(n_19811) );
no02f80 g550282 ( .a(n_19502), .b(x_in_22_4), .o(n_19810) );
na02f80 g550283 ( .a(n_19501), .b(x_in_54_4), .o(n_20528) );
in01f80 g550284 ( .a(n_19808), .o(n_19809) );
no02f80 g550285 ( .a(n_19501), .b(x_in_54_4), .o(n_19808) );
na02f80 g550286 ( .a(n_18641), .b(x_in_2_5), .o(n_19551) );
in01f80 g550287 ( .a(n_18965), .o(n_18966) );
no02f80 g550288 ( .a(n_18641), .b(x_in_2_5), .o(n_18965) );
no02f80 g550289 ( .a(n_18091), .b(n_17807), .o(n_17808) );
na02f80 g550290 ( .a(n_18363), .b(x_in_52_4), .o(n_19316) );
in01f80 g550291 ( .a(n_18639), .o(n_18640) );
no02f80 g550292 ( .a(n_18363), .b(x_in_52_4), .o(n_18639) );
na02f80 g550293 ( .a(n_18655), .b(n_18361), .o(n_18362) );
na02f80 g550294 ( .a(n_18964), .b(x_in_22_5), .o(n_19885) );
in01f80 g550295 ( .a(n_19263), .o(n_19264) );
no02f80 g550296 ( .a(n_18964), .b(x_in_22_5), .o(n_19263) );
no02f80 g550297 ( .a(n_20163), .b(n_20162), .o(n_20164) );
na02f80 g550298 ( .a(n_18943), .b(x_in_40_4), .o(n_19888) );
no02f80 g550299 ( .a(n_19261), .b(n_19260), .o(n_19262) );
in01f80 g550300 ( .a(n_19806), .o(n_19807) );
no02f80 g550301 ( .a(n_19486), .b(x_in_14_4), .o(n_19806) );
no02f80 g550302 ( .a(n_19258), .b(n_19257), .o(n_19259) );
na02f80 g550303 ( .a(n_19500), .b(x_in_46_4), .o(n_20529) );
in01f80 g550304 ( .a(n_19804), .o(n_19805) );
no02f80 g550305 ( .a(n_19500), .b(x_in_46_4), .o(n_19804) );
in01f80 g550306 ( .a(n_19802), .o(n_19803) );
no02f80 g550307 ( .a(n_19492), .b(x_in_30_4), .o(n_19802) );
no02f80 g550308 ( .a(n_20160), .b(n_20159), .o(n_20161) );
na02f80 g550309 ( .a(n_18638), .b(x_in_54_5), .o(n_19550) );
in01f80 g550310 ( .a(n_18962), .o(n_18963) );
no02f80 g550311 ( .a(n_18638), .b(x_in_54_5), .o(n_18962) );
in01f80 g550312 ( .a(n_19800), .o(n_19801) );
no02f80 g550313 ( .a(n_19499), .b(x_in_62_4), .o(n_19800) );
no02f80 g550314 ( .a(n_20157), .b(n_20156), .o(n_20158) );
no02f80 g550315 ( .a(n_20154), .b(n_20153), .o(n_20155) );
no02f80 g550316 ( .a(n_18292), .b(n_18976), .o(n_19984) );
na02f80 g550317 ( .a(n_18961), .b(x_in_56_6), .o(n_19869) );
no02f80 g550318 ( .a(n_18382), .b(n_18083), .o(n_18084) );
in01f80 g550319 ( .a(n_19798), .o(n_19799) );
no02f80 g550320 ( .a(n_19485), .b(x_in_36_4), .o(n_19798) );
na02f80 g550321 ( .a(n_18387), .b(n_18081), .o(n_18082) );
na02f80 g550322 ( .a(n_18637), .b(x_in_14_5), .o(n_19549) );
in01f80 g550323 ( .a(n_18959), .o(n_18960) );
no02f80 g550324 ( .a(n_18637), .b(x_in_14_5), .o(n_18959) );
no02f80 g550325 ( .a(n_19255), .b(n_19254), .o(n_19256) );
na02f80 g550326 ( .a(n_18958), .b(x_in_34_5), .o(n_19884) );
in01f80 g550327 ( .a(n_19252), .o(n_19253) );
no02f80 g550328 ( .a(n_18958), .b(x_in_34_5), .o(n_19252) );
na02f80 g550329 ( .a(n_18386), .b(n_18079), .o(n_18080) );
na02f80 g550330 ( .a(n_18636), .b(x_in_46_5), .o(n_19548) );
in01f80 g550331 ( .a(n_18956), .o(n_18957) );
no02f80 g550332 ( .a(n_18636), .b(x_in_46_5), .o(n_18956) );
no02f80 g550333 ( .a(n_19250), .b(n_19249), .o(n_19251) );
no02f80 g550334 ( .a(n_18385), .b(n_18077), .o(n_18078) );
na02f80 g550335 ( .a(n_18635), .b(x_in_16_5), .o(n_19547) );
in01f80 g550336 ( .a(n_18954), .o(n_18955) );
no02f80 g550337 ( .a(n_18635), .b(x_in_16_5), .o(n_18954) );
no02f80 g550338 ( .a(n_19497), .b(n_19496), .o(n_19498) );
no02f80 g550339 ( .a(n_19494), .b(n_19493), .o(n_19495) );
no02f80 g550340 ( .a(n_19796), .b(n_19795), .o(n_19797) );
no02f80 g550341 ( .a(n_19247), .b(n_19246), .o(n_19248) );
na02f80 g550342 ( .a(n_18384), .b(n_18075), .o(n_18076) );
na02f80 g550343 ( .a(n_18634), .b(x_in_30_5), .o(n_19546) );
in01f80 g550344 ( .a(n_18952), .o(n_18953) );
no02f80 g550345 ( .a(n_18634), .b(x_in_30_5), .o(n_18952) );
na02f80 g550346 ( .a(n_18633), .b(x_in_18_5), .o(n_19544) );
in01f80 g550347 ( .a(n_18950), .o(n_18951) );
no02f80 g550348 ( .a(n_18633), .b(x_in_18_5), .o(n_18950) );
no02f80 g550349 ( .a(n_19244), .b(n_19243), .o(n_19245) );
na02f80 g550350 ( .a(n_18949), .b(x_in_12_5), .o(n_19882) );
in01f80 g550351 ( .a(n_19241), .o(n_19242) );
no02f80 g550352 ( .a(n_18949), .b(x_in_12_5), .o(n_19241) );
na02f80 g550353 ( .a(n_18383), .b(n_18073), .o(n_18074) );
na02f80 g550354 ( .a(n_18632), .b(x_in_62_5), .o(n_19545) );
in01f80 g550355 ( .a(n_18947), .o(n_18948) );
no02f80 g550356 ( .a(n_18632), .b(x_in_62_5), .o(n_18947) );
no02f80 g550357 ( .a(n_19239), .b(n_19238), .o(n_19240) );
na02f80 g550358 ( .a(n_19492), .b(x_in_30_4), .o(n_20531) );
no02f80 g550359 ( .a(n_18945), .b(n_18944), .o(n_18946) );
na02f80 g550360 ( .a(n_19491), .b(x_in_32_3), .o(n_20525) );
in01f80 g550361 ( .a(n_19793), .o(n_19794) );
no02f80 g550362 ( .a(n_19491), .b(x_in_32_3), .o(n_19793) );
in01f80 g550363 ( .a(n_19236), .o(n_19237) );
no02f80 g550364 ( .a(n_18943), .b(x_in_40_4), .o(n_19236) );
na02f80 g550365 ( .a(n_19235), .b(x_in_16_4), .o(n_20215) );
in01f80 g550366 ( .a(n_19489), .o(n_19490) );
no02f80 g550367 ( .a(n_19235), .b(x_in_16_4), .o(n_19489) );
no02f80 g550368 ( .a(n_19791), .b(n_19790), .o(n_19792) );
na02f80 g550369 ( .a(n_18631), .b(x_in_50_5), .o(n_19539) );
in01f80 g550370 ( .a(n_18941), .o(n_18942) );
no02f80 g550371 ( .a(n_18631), .b(x_in_50_5), .o(n_18941) );
no02f80 g550372 ( .a(n_20151), .b(n_20150), .o(n_20152) );
no02f80 g550373 ( .a(n_19233), .b(n_19232), .o(n_19234) );
no02f80 g550374 ( .a(n_19230), .b(n_19229), .o(n_19231) );
na02f80 g550375 ( .a(n_19228), .b(n_18563), .o(n_19863) );
na02f80 g550376 ( .a(n_19227), .b(x_in_26_4), .o(n_20209) );
in01f80 g550377 ( .a(n_18939), .o(n_18940) );
no02f80 g550378 ( .a(n_18630), .b(x_in_58_5), .o(n_18939) );
na02f80 g550379 ( .a(n_18938), .b(x_in_8_6), .o(n_19881) );
in01f80 g550380 ( .a(n_19225), .o(n_19226) );
no02f80 g550381 ( .a(n_18938), .b(x_in_8_6), .o(n_19225) );
no02f80 g550382 ( .a(n_18654), .b(n_18359), .o(n_18360) );
na02f80 g550383 ( .a(n_18630), .b(x_in_58_5), .o(n_19552) );
no02f80 g550384 ( .a(n_19223), .b(n_19222), .o(n_19224) );
na02f80 g550385 ( .a(n_19471), .b(x_in_44_6), .o(n_20212) );
na02f80 g550386 ( .a(n_18937), .b(x_in_40_3), .o(n_19880) );
in01f80 g550387 ( .a(n_19487), .o(n_19488) );
no02f80 g550388 ( .a(n_19471), .b(x_in_44_6), .o(n_19487) );
in01f80 g550389 ( .a(n_19220), .o(n_19221) );
no02f80 g550390 ( .a(n_18937), .b(x_in_40_3), .o(n_19220) );
na02f80 g550391 ( .a(n_18629), .b(x_in_32_4), .o(n_19538) );
in01f80 g550392 ( .a(n_18935), .o(n_18936) );
no02f80 g550393 ( .a(n_18629), .b(x_in_32_4), .o(n_18935) );
na02f80 g550394 ( .a(n_19486), .b(x_in_14_4), .o(n_20524) );
no02f80 g550395 ( .a(n_19788), .b(n_19787), .o(n_19789) );
no02f80 g550396 ( .a(n_19785), .b(n_19784), .o(n_19786) );
in01f80 g550397 ( .a(n_20148), .o(n_20149) );
na02f80 g550398 ( .a(n_19783), .b(n_19138), .o(n_20148) );
in01f80 g550399 ( .a(n_19218), .o(n_19219) );
na02f80 g550400 ( .a(n_18934), .b(n_18308), .o(n_19218) );
no02f80 g550401 ( .a(n_18381), .b(n_18071), .o(n_18072) );
no02f80 g550402 ( .a(n_18018), .b(n_18620), .o(n_19613) );
na02f80 g550403 ( .a(n_18628), .b(x_in_56_5), .o(n_19535) );
in01f80 g550404 ( .a(n_18932), .o(n_18933) );
no02f80 g550405 ( .a(n_18628), .b(x_in_56_5), .o(n_18932) );
no02f80 g550406 ( .a(n_19216), .b(n_19215), .o(n_19217) );
na02f80 g550407 ( .a(n_18627), .b(x_in_10_5), .o(n_19534) );
in01f80 g550408 ( .a(n_18930), .o(n_18931) );
no02f80 g550409 ( .a(n_18627), .b(x_in_10_5), .o(n_18930) );
na02f80 g550410 ( .a(n_18929), .b(x_in_48_4), .o(n_19874) );
in01f80 g550411 ( .a(n_19213), .o(n_19214) );
no02f80 g550412 ( .a(n_18929), .b(x_in_48_4), .o(n_19213) );
na02f80 g550413 ( .a(n_19485), .b(x_in_36_4), .o(n_20527) );
no02f80 g550414 ( .a(n_19211), .b(n_19210), .o(n_19212) );
no02f80 g550415 ( .a(n_19301), .b(n_18927), .o(n_18928) );
na02f80 g550416 ( .a(n_19209), .b(n_18558), .o(n_19876) );
in01f80 g550417 ( .a(n_19483), .o(n_19484) );
no02f80 g550418 ( .a(n_19271), .b(x_in_20_4), .o(n_19483) );
na02f80 g550419 ( .a(n_19775), .b(x_in_60_3), .o(n_20907) );
no02f80 g550420 ( .a(n_19781), .b(n_19780), .o(n_19782) );
na02f80 g550421 ( .a(n_18626), .b(x_in_10_4), .o(n_19556) );
na02f80 g550422 ( .a(n_18625), .b(x_in_42_5), .o(n_19533) );
in01f80 g550423 ( .a(n_18925), .o(n_18926) );
no02f80 g550424 ( .a(n_18625), .b(x_in_42_5), .o(n_18925) );
no02f80 g550425 ( .a(n_19300), .b(n_18923), .o(n_18924) );
na02f80 g550426 ( .a(n_19779), .b(x_in_36_3), .o(n_20906) );
in01f80 g550427 ( .a(n_20146), .o(n_20147) );
no02f80 g550428 ( .a(n_19779), .b(x_in_36_3), .o(n_20146) );
no02f80 g550429 ( .a(n_19207), .b(n_19206), .o(n_19208) );
in01f80 g550430 ( .a(n_20144), .o(n_20145) );
na02f80 g550431 ( .a(n_19778), .b(n_19134), .o(n_20144) );
no02f80 g550432 ( .a(n_18988), .b(n_18623), .o(n_18624) );
no02f80 g550433 ( .a(n_18388), .b(n_18069), .o(n_18070) );
no02f80 g550434 ( .a(n_18019), .b(n_18623), .o(n_19617) );
in01f80 g550435 ( .a(n_19204), .o(n_19205) );
na02f80 g550436 ( .a(n_18922), .b(n_18306), .o(n_19204) );
na02f80 g550437 ( .a(n_20143), .b(x_in_20_3), .o(n_21195) );
in01f80 g550438 ( .a(n_20487), .o(n_20488) );
no02f80 g550439 ( .a(n_20143), .b(x_in_20_3), .o(n_20487) );
na02f80 g550440 ( .a(n_18622), .b(x_in_26_5), .o(n_19532) );
in01f80 g550441 ( .a(n_18920), .o(n_18921) );
no02f80 g550442 ( .a(n_18622), .b(x_in_26_5), .o(n_18920) );
no02f80 g550443 ( .a(n_18982), .b(n_18620), .o(n_18621) );
no02f80 g550444 ( .a(n_19481), .b(n_19480), .o(n_19482) );
na02f80 g550445 ( .a(n_19203), .b(x_in_52_3), .o(n_20207) );
in01f80 g550446 ( .a(n_19478), .o(n_19479) );
no02f80 g550447 ( .a(n_19203), .b(x_in_52_3), .o(n_19478) );
in01f80 g550448 ( .a(n_18618), .o(n_18619) );
na02f80 g550449 ( .a(n_18358), .b(n_17796), .o(n_18618) );
no02f80 g550450 ( .a(n_19201), .b(n_19200), .o(n_19202) );
na02f80 g550451 ( .a(n_19477), .b(x_in_12_4), .o(n_20521) );
in01f80 g550452 ( .a(n_19776), .o(n_19777) );
no02f80 g550453 ( .a(n_19477), .b(x_in_12_4), .o(n_19776) );
no02f80 g550454 ( .a(n_19198), .b(n_19197), .o(n_19199) );
no02f80 g550455 ( .a(n_20141), .b(n_20140), .o(n_20142) );
na02f80 g550456 ( .a(n_18919), .b(x_in_8_7), .o(n_19886) );
no02f80 g550457 ( .a(n_19195), .b(n_19194), .o(n_19196) );
no02f80 g550458 ( .a(n_20138), .b(n_20137), .o(n_20139) );
in01f80 g550459 ( .a(n_19192), .o(n_19193) );
no02f80 g550460 ( .a(n_18919), .b(x_in_8_7), .o(n_19192) );
in01f80 g550461 ( .a(n_20135), .o(n_20136) );
no02f80 g550462 ( .a(n_19775), .b(x_in_60_3), .o(n_20135) );
na02f80 g550463 ( .a(n_18918), .b(x_in_60_4), .o(n_19873) );
in01f80 g550464 ( .a(n_19190), .o(n_19191) );
no02f80 g550465 ( .a(n_18918), .b(x_in_60_4), .o(n_19190) );
na02f80 g550466 ( .a(n_18653), .b(n_18356), .o(n_18357) );
na02f80 g550467 ( .a(n_18090), .b(n_17805), .o(n_17806) );
no02f80 g550468 ( .a(n_18380), .b(n_18067), .o(n_18068) );
no02f80 g550469 ( .a(n_19001), .b(n_18616), .o(n_18617) );
no02f80 g550470 ( .a(n_18652), .b(n_18354), .o(n_18355) );
no02f80 g550471 ( .a(n_19299), .b(n_18916), .o(n_18917) );
no02f80 g550472 ( .a(n_18651), .b(n_18352), .o(n_18353) );
na02f80 g550473 ( .a(n_18379), .b(n_18065), .o(n_18066) );
no02f80 g550474 ( .a(n_19298), .b(n_18914), .o(n_18915) );
no02f80 g550475 ( .a(n_18378), .b(n_18063), .o(n_18064) );
no02f80 g550476 ( .a(n_18650), .b(n_18350), .o(n_18351) );
na02f80 g550477 ( .a(n_18089), .b(n_17803), .o(n_17804) );
na02f80 g550478 ( .a(n_18912), .b(n_18911), .o(n_18913) );
no02f80 g550479 ( .a(n_18964), .b(n_18910), .o(n_19931) );
na02f80 g550480 ( .a(n_18908), .b(n_18910), .o(n_18909) );
no02f80 g550481 ( .a(n_18638), .b(n_18911), .o(n_19603) );
no02f80 g550482 ( .a(n_18637), .b(n_18907), .o(n_19602) );
na02f80 g550483 ( .a(n_18905), .b(n_18907), .o(n_18906) );
no02f80 g550484 ( .a(n_18636), .b(n_18904), .o(n_19601) );
na02f80 g550485 ( .a(n_18902), .b(n_18904), .o(n_18903) );
no02f80 g550486 ( .a(n_18634), .b(n_18901), .o(n_19605) );
na02f80 g550487 ( .a(n_18899), .b(n_18901), .o(n_18900) );
no02f80 g550488 ( .a(n_18632), .b(n_18898), .o(n_19606) );
na02f80 g550489 ( .a(n_18896), .b(n_18898), .o(n_18897) );
no02f80 g550490 ( .a(n_18919), .b(n_18895), .o(n_20253) );
na02f80 g550491 ( .a(n_18614), .b(n_18895), .o(n_18615) );
no02f80 g550492 ( .a(n_18949), .b(n_18894), .o(n_19930) );
na02f80 g550493 ( .a(n_18892), .b(n_18894), .o(n_18893) );
no02f80 g550494 ( .a(n_19000), .b(n_18612), .o(n_18613) );
no02f80 g550495 ( .a(n_18377), .b(n_18061), .o(n_18062) );
no02f80 g550496 ( .a(n_18376), .b(n_18059), .o(n_18060) );
no02f80 g550497 ( .a(n_19835), .b(n_19475), .o(n_19476) );
no02f80 g550498 ( .a(n_18812), .b(n_19475), .o(n_20561) );
na02f80 g550499 ( .a(n_19474), .b(n_19473), .o(n_20560) );
na02f80 g550500 ( .a(n_19474), .b(n_19471), .o(n_19472) );
no02f80 g550501 ( .a(n_18649), .b(n_18348), .o(n_18349) );
no02f80 g550502 ( .a(n_18375), .b(n_18057), .o(n_18058) );
no02f80 g550503 ( .a(n_18374), .b(n_18055), .o(n_18056) );
no02f80 g550504 ( .a(n_18373), .b(n_18053), .o(n_18054) );
no02f80 g550505 ( .a(n_18289), .b(n_18890), .o(n_19927) );
no02f80 g550506 ( .a(n_19278), .b(n_18890), .o(n_18891) );
na02f80 g550507 ( .a(n_18372), .b(n_18051), .o(n_18052) );
no02f80 g550508 ( .a(n_18346), .b(n_18345), .o(n_18347) );
na02f80 g550509 ( .a(n_18050), .b(n_18345), .o(n_19339) );
no02f80 g550510 ( .a(n_18087), .b(n_17801), .o(n_17802) );
no02f80 g550511 ( .a(n_17158), .b(n_17801), .o(n_18663) );
no02f80 g550512 ( .a(n_18371), .b(n_18048), .o(n_18049) );
no02f80 g550513 ( .a(n_20485), .b(n_20484), .o(n_20486) );
no02f80 g550514 ( .a(n_20133), .b(n_20132), .o(n_20134) );
no02f80 g550515 ( .a(n_19469), .b(n_19468), .o(n_19470) );
no02f80 g550516 ( .a(n_19466), .b(n_19465), .o(n_19467) );
no02f80 g550517 ( .a(n_20482), .b(n_20481), .o(n_20483) );
no02f80 g550518 ( .a(n_20880), .b(n_20879), .o(n_20881) );
no02f80 g550519 ( .a(n_19463), .b(n_19462), .o(n_19464) );
no02f80 g550520 ( .a(n_18888), .b(n_18887), .o(n_18889) );
na02f80 g550521 ( .a(n_18885), .b(n_18187), .o(n_19585) );
na02f80 g550522 ( .a(n_18885), .b(n_18884), .o(n_18886) );
na02f80 g550523 ( .a(n_18882), .b(n_18881), .o(n_18883) );
na02f80 g550524 ( .a(n_18343), .b(n_18596), .o(n_18344) );
in01f80 g550525 ( .a(n_18880), .o(n_19582) );
no02f80 g550526 ( .a(n_18631), .b(n_18611), .o(n_18880) );
na02f80 g550527 ( .a(n_18341), .b(n_18611), .o(n_18342) );
in01f80 g550528 ( .a(n_18879), .o(n_19586) );
na02f80 g550529 ( .a(FE_OFN1059_n_18610), .b(n_18887), .o(n_18879) );
na02f80 g550530 ( .a(n_18609), .b(n_17953), .o(n_19581) );
na02f80 g550531 ( .a(n_18609), .b(n_18339), .o(n_18340) );
na02f80 g550532 ( .a(n_18597), .b(n_18337), .o(n_18338) );
na02f80 g550533 ( .a(n_18877), .b(n_18876), .o(n_18878) );
na02f80 g550534 ( .a(n_18335), .b(n_18605), .o(n_18336) );
na02f80 g550535 ( .a(n_19773), .b(n_19460), .o(n_19461) );
na02f80 g550536 ( .a(n_18877), .b(n_18185), .o(n_19579) );
no02f80 g550537 ( .a(n_18608), .b(n_17950), .o(n_19916) );
no02f80 g550538 ( .a(n_18608), .b(n_18606), .o(n_18607) );
na02f80 g550539 ( .a(n_18533), .b(n_19189), .o(n_20242) );
ao12f80 g550540 ( .a(n_10837), .b(n_18334), .c(n_12062), .o(n_19322) );
in01f80 g550541 ( .a(n_19459), .o(n_20247) );
no02f80 g550542 ( .a(n_18629), .b(n_19188), .o(n_19459) );
na02f80 g550543 ( .a(n_19186), .b(n_19188), .o(n_19187) );
in01f80 g550544 ( .a(n_21237), .o(n_19185) );
oa12f80 g550545 ( .a(n_18837), .b(n_18252), .c(n_17620), .o(n_21237) );
no02f80 g550546 ( .a(n_18332), .b(n_18331), .o(n_18333) );
in01f80 g550547 ( .a(n_18330), .o(n_19018) );
na02f80 g550548 ( .a(n_18047), .b(n_18331), .o(n_18330) );
ao12f80 g550549 ( .a(n_5794), .b(n_16886), .c(n_6646), .o(n_17810) );
in01f80 g550550 ( .a(n_19184), .o(n_19913) );
no02f80 g550551 ( .a(n_18635), .b(n_18875), .o(n_19184) );
na02f80 g550552 ( .a(n_18873), .b(n_18875), .o(n_18874) );
in01f80 g550553 ( .a(n_18872), .o(n_19576) );
no02f80 g550554 ( .a(n_18630), .b(n_18605), .o(n_18872) );
in01f80 g550555 ( .a(n_19183), .o(n_19910) );
no02f80 g550556 ( .a(n_18871), .b(n_18929), .o(n_19183) );
na02f80 g550557 ( .a(n_18871), .b(n_18869), .o(n_18870) );
na02f80 g550558 ( .a(n_18918), .b(n_19189), .o(n_18868) );
no02f80 g550559 ( .a(n_18603), .b(n_18602), .o(n_18604) );
no02f80 g550560 ( .a(n_18603), .b(n_17945), .o(n_19570) );
na02f80 g550561 ( .a(n_18644), .b(n_18862), .o(n_18601) );
in01f80 g550562 ( .a(n_21246), .o(n_19774) );
oa12f80 g550563 ( .a(n_19433), .b(n_18785), .c(n_18172), .o(n_21246) );
in01f80 g550564 ( .a(n_19182), .o(n_19907) );
no02f80 g550565 ( .a(n_18943), .b(n_18867), .o(n_19182) );
na02f80 g550566 ( .a(n_18599), .b(n_18867), .o(n_18600) );
in01f80 g550567 ( .a(n_20590), .o(n_19181) );
oa12f80 g550568 ( .a(n_18830), .b(n_18247), .c(n_17862), .o(n_20590) );
in01f80 g550569 ( .a(n_21596), .o(n_20131) );
oa12f80 g550570 ( .a(n_19745), .b(n_19078), .c(n_18420), .o(n_21596) );
in01f80 g550571 ( .a(n_19290), .o(n_18598) );
na02f80 g550572 ( .a(n_17779), .b(n_12170), .o(n_19290) );
na02f80 g550573 ( .a(n_18882), .b(n_18186), .o(n_19923) );
na02f80 g550574 ( .a(n_18597), .b(n_17955), .o(n_19580) );
in01f80 g550575 ( .a(n_18866), .o(n_19563) );
no02f80 g550576 ( .a(n_18633), .b(n_18596), .o(n_18866) );
na02f80 g550577 ( .a(n_18595), .b(n_17943), .o(n_20245) );
na02f80 g550578 ( .a(n_18595), .b(n_18593), .o(n_18594) );
no02f80 g550579 ( .a(n_18591), .b(n_18590), .o(n_18592) );
in01f80 g550580 ( .a(n_18589), .o(n_19329) );
na02f80 g550581 ( .a(n_18329), .b(n_18590), .o(n_18589) );
in01f80 g550582 ( .a(n_21593), .o(n_20480) );
oa12f80 g550583 ( .a(n_19740), .b(n_19081), .c(n_19065), .o(n_21593) );
in01f80 g550584 ( .a(n_18588), .o(n_19325) );
na02f80 g550585 ( .a(n_18328), .b(n_18585), .o(n_18588) );
na02f80 g550586 ( .a(n_19271), .b(n_19458), .o(n_19180) );
na02f80 g550587 ( .a(n_19773), .b(n_19066), .o(n_20558) );
in01f80 g550588 ( .a(n_20243), .o(n_19772) );
na02f80 g550589 ( .a(n_18805), .b(n_19458), .o(n_20243) );
in01f80 g550590 ( .a(n_21984), .o(n_20479) );
oa12f80 g550591 ( .a(n_20108), .b(n_19398), .c(n_18693), .o(n_21984) );
in01f80 g550592 ( .a(n_19179), .o(n_19902) );
no02f80 g550593 ( .a(n_18865), .b(n_18363), .o(n_19179) );
na02f80 g550594 ( .a(n_18865), .b(n_18863), .o(n_18864) );
in01f80 g550595 ( .a(n_20926), .o(n_19178) );
oa12f80 g550596 ( .a(n_18832), .b(n_18234), .c(n_17617), .o(n_20926) );
no02f80 g550597 ( .a(n_18586), .b(n_18585), .o(n_18587) );
in01f80 g550598 ( .a(n_19566), .o(n_19177) );
na02f80 g550599 ( .a(n_18294), .b(n_18862), .o(n_19566) );
in01f80 g550600 ( .a(n_20953), .o(n_20130) );
oa12f80 g550601 ( .a(n_19147), .b(n_18716), .c(n_18517), .o(n_20953) );
in01f80 g550602 ( .a(n_20619), .o(n_20129) );
oa12f80 g550603 ( .a(n_18312), .b(n_17767), .c(n_18706), .o(n_20619) );
in01f80 g550604 ( .a(n_20649), .o(n_20128) );
oa12f80 g550605 ( .a(n_19435), .b(n_18714), .c(n_18789), .o(n_20649) );
in01f80 g550606 ( .a(n_20947), .o(n_20127) );
oa12f80 g550607 ( .a(n_19148), .b(n_18515), .c(n_18715), .o(n_20947) );
in01f80 g550608 ( .a(n_20646), .o(n_20126) );
oa12f80 g550609 ( .a(n_19423), .b(n_18787), .c(n_18713), .o(n_20646) );
in01f80 g550610 ( .a(n_20308), .o(n_19771) );
oa12f80 g550611 ( .a(n_19146), .b(n_18444), .c(n_18511), .o(n_20308) );
in01f80 g550612 ( .a(n_20295), .o(n_19770) );
oa12f80 g550613 ( .a(n_19145), .b(n_18443), .c(n_18509), .o(n_20295) );
oa12f80 g550614 ( .a(n_12434), .b(n_18046), .c(n_13627), .o(n_19017) );
in01f80 g550615 ( .a(n_20278), .o(n_19769) );
oa12f80 g550616 ( .a(n_19144), .b(n_18440), .c(n_18507), .o(n_20278) );
in01f80 g550617 ( .a(n_19768), .o(n_20912) );
oa12f80 g550618 ( .a(n_17349), .b(n_19448), .c(n_16746), .o(n_19768) );
in01f80 g550619 ( .a(n_19457), .o(n_20553) );
oa12f80 g550620 ( .a(n_18781), .b(n_19176), .c(n_18135), .o(n_19457) );
in01f80 g550621 ( .a(n_21260), .o(n_19767) );
oa12f80 g550622 ( .a(n_19432), .b(n_18439), .c(n_18767), .o(n_21260) );
in01f80 g550623 ( .a(n_21255), .o(n_19766) );
oa12f80 g550624 ( .a(n_19425), .b(n_18438), .c(n_18779), .o(n_21255) );
in01f80 g550625 ( .a(n_21252), .o(n_19765) );
oa12f80 g550626 ( .a(n_19430), .b(n_18441), .c(n_18775), .o(n_21252) );
in01f80 g550627 ( .a(n_20290), .o(n_19764) );
oa12f80 g550628 ( .a(n_18840), .b(n_18437), .c(n_18263), .o(n_20290) );
in01f80 g550629 ( .a(n_20628), .o(n_20125) );
oa12f80 g550630 ( .a(n_18566), .b(n_18000), .c(n_18704), .o(n_20628) );
in01f80 g550631 ( .a(n_20643), .o(n_20124) );
oa12f80 g550632 ( .a(n_18560), .b(n_18004), .c(n_18712), .o(n_20643) );
in01f80 g550633 ( .a(n_20633), .o(n_20123) );
oa12f80 g550634 ( .a(n_18569), .b(n_17996), .c(n_18711), .o(n_20633) );
in01f80 g550635 ( .a(n_21249), .o(n_19763) );
oa12f80 g550636 ( .a(n_19424), .b(n_18435), .c(n_18773), .o(n_21249) );
in01f80 g550637 ( .a(n_21224), .o(n_19762) );
oa12f80 g550638 ( .a(n_19420), .b(n_18434), .c(n_18763), .o(n_21224) );
in01f80 g550639 ( .a(n_19456), .o(n_20545) );
oa12f80 g550640 ( .a(n_17745), .b(n_19170), .c(n_17112), .o(n_19456) );
in01f80 g550641 ( .a(n_18861), .o(n_19897) );
oa12f80 g550642 ( .a(n_2874), .b(n_18580), .c(n_2194), .o(n_18861) );
in01f80 g550643 ( .a(n_21234), .o(n_20478) );
oa12f80 g550644 ( .a(n_19426), .b(n_18771), .c(n_19068), .o(n_21234) );
in01f80 g550645 ( .a(n_20616), .o(n_20122) );
oa12f80 g550646 ( .a(n_18318), .b(n_17765), .c(n_18703), .o(n_20616) );
in01f80 g550647 ( .a(n_21243), .o(n_20878) );
oa12f80 g550648 ( .a(n_18839), .b(n_18259), .c(n_19397), .o(n_21243) );
in01f80 g550649 ( .a(n_20613), .o(n_20121) );
oa12f80 g550650 ( .a(n_18317), .b(n_17763), .c(n_18702), .o(n_20613) );
in01f80 g550651 ( .a(n_20287), .o(n_19761) );
oa12f80 g550652 ( .a(n_18564), .b(n_17993), .c(n_18426), .o(n_20287) );
in01f80 g550653 ( .a(n_20610), .o(n_20120) );
oa12f80 g550654 ( .a(n_18316), .b(n_17759), .c(n_18701), .o(n_20610) );
in01f80 g550655 ( .a(n_20284), .o(n_19760) );
oa12f80 g550656 ( .a(n_18314), .b(n_17757), .c(n_18425), .o(n_20284) );
in01f80 g550657 ( .a(n_21240), .o(n_19759) );
oa12f80 g550658 ( .a(n_19431), .b(n_18436), .c(n_18777), .o(n_21240) );
in01f80 g550659 ( .a(n_20597), .o(n_20119) );
oa12f80 g550660 ( .a(n_18561), .b(n_17991), .c(n_18700), .o(n_20597) );
in01f80 g550661 ( .a(n_20607), .o(n_20118) );
oa12f80 g550662 ( .a(n_18315), .b(n_17755), .c(n_18699), .o(n_20607) );
in01f80 g550663 ( .a(n_20652), .o(n_20117) );
oa12f80 g550664 ( .a(n_18559), .b(n_17998), .c(n_18705), .o(n_20652) );
in01f80 g550665 ( .a(n_19175), .o(n_20234) );
oa12f80 g550666 ( .a(n_15275), .b(n_18856), .c(n_14505), .o(n_19175) );
in01f80 g550667 ( .a(n_20944), .o(n_19758) );
oa12f80 g550668 ( .a(n_19135), .b(n_18442), .c(n_18504), .o(n_20944) );
in01f80 g550669 ( .a(n_20936), .o(n_19455) );
oa12f80 g550670 ( .a(n_19140), .b(n_18481), .c(n_18182), .o(n_20936) );
in01f80 g550671 ( .a(n_18860), .o(n_19895) );
oa12f80 g550672 ( .a(n_3254), .b(n_18578), .c(n_2257), .o(n_18860) );
in01f80 g550673 ( .a(n_20594), .o(n_20116) );
oa12f80 g550674 ( .a(n_18311), .b(n_17753), .c(n_18698), .o(n_20594) );
ao12f80 g550675 ( .a(n_9425), .b(n_18584), .c(n_9424), .o(n_19568) );
in01f80 g550676 ( .a(n_19757), .o(n_20917) );
oa12f80 g550677 ( .a(n_18474), .b(n_19454), .c(n_17899), .o(n_19757) );
in01f80 g550678 ( .a(n_20267), .o(n_19756) );
oa12f80 g550679 ( .a(n_19136), .b(n_18475), .c(n_18432), .o(n_20267) );
in01f80 g550680 ( .a(n_18859), .o(n_19900) );
oa12f80 g550681 ( .a(n_18245), .b(n_18583), .c(n_17690), .o(n_18859) );
oa12f80 g550682 ( .a(n_13130), .b(n_18327), .c(n_14277), .o(n_19321) );
in01f80 g550683 ( .a(n_20582), .o(n_20115) );
oa12f80 g550684 ( .a(n_18303), .b(n_18696), .c(n_17748), .o(n_20582) );
in01f80 g550685 ( .a(n_19453), .o(n_20540) );
oa12f80 g550686 ( .a(n_17044), .b(n_19165), .c(n_16542), .o(n_19453) );
in01f80 g550687 ( .a(n_20950), .o(n_20477) );
oa12f80 g550688 ( .a(n_18836), .b(n_18240), .c(n_19067), .o(n_20950) );
in01f80 g550689 ( .a(n_19174), .o(n_20229) );
oa12f80 g550690 ( .a(n_15108), .b(n_18854), .c(n_14500), .o(n_19174) );
in01f80 g550691 ( .a(n_20578), .o(n_20114) );
oa12f80 g550692 ( .a(n_18302), .b(n_18695), .c(n_17746), .o(n_20578) );
in01f80 g550693 ( .a(n_20568), .o(n_20113) );
oa12f80 g550694 ( .a(n_18555), .b(n_18697), .c(n_17966), .o(n_20568) );
in01f80 g550695 ( .a(n_21229), .o(n_19755) );
oa12f80 g550696 ( .a(n_19419), .b(n_18765), .c(n_18428), .o(n_21229) );
in01f80 g550697 ( .a(n_19452), .o(n_20548) );
oa12f80 g550698 ( .a(n_18556), .b(n_18181), .c(n_17968), .o(n_19452) );
in01f80 g550699 ( .a(n_19451), .o(n_20547) );
oa12f80 g550700 ( .a(n_18784), .b(n_19173), .c(n_18120), .o(n_19451) );
in01f80 g550701 ( .a(n_20258), .o(n_19754) );
oa12f80 g550702 ( .a(n_18321), .b(n_18423), .c(n_17736), .o(n_20258) );
in01f80 g550703 ( .a(n_20640), .o(n_20112) );
oa12f80 g550704 ( .a(n_18843), .b(n_18273), .c(n_18717), .o(n_20640) );
oa12f80 g550705 ( .a(n_12280), .b(n_18326), .c(n_12499), .o(n_19336) );
oa12f80 g550706 ( .a(n_12273), .b(n_17800), .c(n_12944), .o(n_18676) );
in01f80 g550707 ( .a(n_18045), .o(n_19016) );
ao12f80 g550708 ( .a(n_7215), .b(n_17799), .c(n_5113), .o(n_18045) );
oa22f80 g550709 ( .a(n_18156), .b(n_8760), .c(n_6637), .d(n_6775), .o(n_20238) );
oa12f80 g550710 ( .a(n_12041), .b(n_18044), .c(n_13112), .o(n_19014) );
ao12f80 g550711 ( .a(n_19131), .b(n_19130), .c(n_19129), .o(n_19753) );
ao12f80 g550712 ( .a(n_18553), .b(n_18851), .c(n_18552), .o(n_19172) );
in01f80 g550713 ( .a(n_18660), .o(n_18325) );
oa12f80 g550714 ( .a(n_17490), .b(n_17800), .c(n_17489), .o(n_18660) );
in01f80 g550715 ( .a(n_19304), .o(n_18582) );
oa12f80 g550716 ( .a(n_17794), .b(n_18046), .c(n_17793), .o(n_19304) );
ao12f80 g550717 ( .a(n_18824), .b(n_18823), .c(n_18822), .o(n_19450) );
oa12f80 g550718 ( .a(n_18546), .b(n_18545), .c(n_18547), .o(n_19887) );
ao22s80 g550719 ( .a(n_19448), .b(n_17586), .c(n_18427), .d(n_17585), .o(n_19449) );
ao22s80 g550720 ( .a(n_19105), .b(n_19176), .c(n_19104), .d(n_18176), .o(n_20111) );
in01f80 g550721 ( .a(n_19309), .o(n_19530) );
ao12f80 g550722 ( .a(n_18040), .b(n_18326), .c(n_18039), .o(n_19309) );
ao22s80 g550723 ( .a(n_17972), .b(n_19170), .c(n_17971), .d(n_18175), .o(n_19171) );
ao22s80 g550724 ( .a(n_18580), .b(n_3407), .c(n_17710), .d(n_3406), .o(n_18581) );
in01f80 g550725 ( .a(n_18858), .o(n_19891) );
oa12f80 g550726 ( .a(n_18038), .b(n_18334), .c(n_18037), .o(n_18858) );
ao22s80 g550727 ( .a(n_18856), .b(n_15676), .c(n_17939), .d(n_15675), .o(n_18857) );
ao12f80 g550728 ( .a(n_18835), .b(n_18834), .c(n_18833), .o(n_19447) );
in01f80 g550729 ( .a(n_17809), .o(n_18096) );
ao12f80 g550730 ( .a(n_16640), .b(n_16886), .c(n_16639), .o(n_17809) );
oa12f80 g550731 ( .a(n_18033), .b(n_18301), .c(n_18032), .o(n_19315) );
ao22s80 g550732 ( .a(n_18578), .b(n_4127), .c(n_17709), .d(n_4126), .o(n_18579) );
ao12f80 g550733 ( .a(n_18828), .b(n_18827), .c(n_18826), .o(n_19446) );
in01f80 g550734 ( .a(n_19169), .o(n_20226) );
oa12f80 g550735 ( .a(n_18310), .b(n_18584), .c(n_18309), .o(n_19169) );
in01f80 g550736 ( .a(n_18390), .o(n_18664) );
ao22s80 g550737 ( .a(n_17799), .b(n_7423), .c(n_16879), .d(n_7422), .o(n_18390) );
ao12f80 g550738 ( .a(n_11826), .b(FE_OFN672_n_17494), .c(n_10699), .o(n_18093) );
in01f80 g550739 ( .a(n_19343), .o(n_18043) );
oa12f80 g550740 ( .a(n_17163), .b(FE_OFN672_n_17494), .c(n_17162), .o(n_19343) );
in01f80 g550741 ( .a(n_18391), .o(n_18672) );
ao12f80 g550742 ( .a(n_17166), .b(n_17165), .c(n_17164), .o(n_18391) );
oa12f80 g550743 ( .a(n_17488), .b(n_17491), .c(n_17792), .o(n_18667) );
ao12f80 g550744 ( .a(n_18541), .b(n_18849), .c(n_18540), .o(n_19168) );
in01f80 g550745 ( .a(n_19302), .o(n_19526) );
ao12f80 g550746 ( .a(n_18035), .b(n_18327), .c(n_18034), .o(n_19302) );
ao22s80 g550747 ( .a(n_18762), .b(n_19454), .c(n_18761), .d(n_18424), .o(n_19752) );
ao22s80 g550748 ( .a(n_18473), .b(n_18583), .c(n_18472), .d(n_17708), .o(n_19445) );
in01f80 g550749 ( .a(n_19307), .o(n_19310) );
ao12f80 g550750 ( .a(n_17791), .b(n_18044), .c(n_17790), .o(n_19307) );
ao12f80 g550751 ( .a(n_18544), .b(n_18543), .c(n_18542), .o(n_19167) );
ao22s80 g550752 ( .a(n_18854), .b(n_15339), .c(n_17937), .d(n_15338), .o(n_18855) );
ao12f80 g550753 ( .a(n_19739), .b(n_19738), .c(n_19737), .o(n_20476) );
ao22s80 g550754 ( .a(n_19165), .b(n_17324), .c(n_18174), .d(n_17323), .o(n_19166) );
ao12f80 g550755 ( .a(n_18030), .b(n_18029), .c(n_18028), .o(n_18577) );
ao12f80 g550756 ( .a(n_17168), .b(n_17492), .c(n_17167), .o(n_17798) );
ao12f80 g550757 ( .a(n_19416), .b(n_19415), .c(n_19414), .o(n_20110) );
in01f80 g550758 ( .a(n_19871), .o(n_19444) );
oa12f80 g550759 ( .a(n_18551), .b(n_18846), .c(n_18825), .o(n_19871) );
oa12f80 g550760 ( .a(n_18550), .b(n_18549), .c(n_18548), .o(n_19870) );
ao22s80 g550761 ( .a(n_19107), .b(n_19173), .c(n_19106), .d(n_18173), .o(n_20109) );
oa22f80 g550762 ( .a(n_18692), .b(FE_OFN309_n_3069), .c(n_1371), .d(FE_OFN128_n_27449), .o(n_19751) );
oa22f80 g550763 ( .a(n_18170), .b(FE_OFN208_n_29661), .c(n_907), .d(FE_OFN122_n_27449), .o(n_19164) );
oa22f80 g550764 ( .a(n_17789), .b(FE_OFN300_n_3069), .c(n_528), .d(FE_OFN329_n_4860), .o(n_18042) );
oa22f80 g550765 ( .a(n_18691), .b(FE_OFN313_n_3069), .c(n_1397), .d(FE_OFN139_n_27449), .o(n_19750) );
oa22f80 g550766 ( .a(n_18554), .b(FE_OFN295_n_3069), .c(n_866), .d(FE_OFN127_n_27449), .o(n_18853) );
oa22f80 g550767 ( .a(n_18418), .b(FE_OFN417_n_28303), .c(n_1437), .d(FE_OFN131_n_27449), .o(n_19443) );
oa22f80 g550768 ( .a(n_18417), .b(FE_OFN308_n_3069), .c(n_1195), .d(FE_OFN1114_rst), .o(n_19442) );
oa22f80 g550769 ( .a(n_18169), .b(FE_OFN299_n_3069), .c(n_1715), .d(FE_OFN136_n_27449), .o(n_19163) );
oa22f80 g550770 ( .a(n_18416), .b(FE_OFN268_n_4280), .c(n_1958), .d(FE_OFN93_n_27449), .o(n_19441) );
oa22f80 g550771 ( .a(n_18168), .b(n_22960), .c(n_787), .d(FE_OFN347_n_4860), .o(n_19162) );
oa22f80 g550772 ( .a(n_18167), .b(FE_OFN256_n_4280), .c(n_211), .d(FE_OFN122_n_27449), .o(n_19161) );
oa22f80 g550773 ( .a(n_18415), .b(FE_OFN204_n_28771), .c(n_623), .d(FE_OFN105_n_27449), .o(n_19440) );
oa22f80 g550774 ( .a(n_18166), .b(FE_OFN248_n_4162), .c(n_548), .d(FE_OFN92_n_27449), .o(n_19160) );
oa22f80 g550775 ( .a(n_17428), .b(n_23813), .c(n_441), .d(FE_OFN89_n_27449), .o(n_18324) );
oa22f80 g550776 ( .a(n_18851), .b(n_22615), .c(n_183), .d(FE_OFN1182_rst), .o(n_18852) );
oa22f80 g550777 ( .a(n_18165), .b(FE_OFN257_n_4280), .c(n_743), .d(FE_OFN336_n_4860), .o(n_19159) );
oa22f80 g550778 ( .a(n_18163), .b(FE_OFN239_n_4162), .c(n_1224), .d(FE_OFN136_n_27449), .o(n_19158) );
oa22f80 g550779 ( .a(n_18157), .b(FE_OFN257_n_4280), .c(n_1607), .d(FE_OFN101_n_27449), .o(n_19157) );
oa22f80 g550780 ( .a(n_18162), .b(FE_OFN236_n_4162), .c(n_283), .d(FE_OFN76_n_27012), .o(n_19156) );
oa22f80 g550781 ( .a(n_18161), .b(FE_OFN236_n_4162), .c(n_279), .d(FE_OFN93_n_27449), .o(n_19155) );
oa22f80 g550782 ( .a(n_18160), .b(FE_OFN1152_n_3069), .c(n_1509), .d(FE_OFN335_n_4860), .o(n_19154) );
oa22f80 g550783 ( .a(n_18159), .b(n_21988), .c(n_379), .d(FE_OFN324_n_4860), .o(n_19153) );
oa22f80 g550784 ( .a(n_18849), .b(n_27933), .c(n_1829), .d(FE_OFN1106_rst), .o(n_18850) );
oa22f80 g550785 ( .a(n_17932), .b(FE_OFN268_n_4280), .c(n_683), .d(FE_OFN93_n_27449), .o(n_18848) );
oa22f80 g550786 ( .a(n_17427), .b(FE_OFN308_n_3069), .c(n_1285), .d(n_27449), .o(n_18323) );
oa22f80 g550787 ( .a(n_18690), .b(FE_OFN307_n_3069), .c(n_141), .d(FE_OFN99_n_27449), .o(n_19749) );
oa22f80 g550788 ( .a(n_18575), .b(FE_OFN297_n_3069), .c(n_1011), .d(FE_OFN141_n_27449), .o(n_18576) );
oa22f80 g550789 ( .a(FE_OFN428_n_17707), .b(n_22960), .c(n_1888), .d(n_27449), .o(n_18574) );
oa22f80 g550790 ( .a(n_18158), .b(FE_OFN240_n_4162), .c(n_9), .d(FE_OFN1119_rst), .o(n_19152) );
oa22f80 g550791 ( .a(n_18689), .b(FE_OFN413_n_28303), .c(n_1110), .d(FE_OFN352_n_4860), .o(n_19748) );
oa22f80 g550792 ( .a(n_17492), .b(FE_OFN235_n_4162), .c(n_1033), .d(FE_OFN335_n_4860), .o(n_17493) );
oa22f80 g550793 ( .a(n_17425), .b(FE_OFN410_n_28303), .c(n_1060), .d(FE_OFN76_n_27012), .o(n_18322) );
oa22f80 g550794 ( .a(FE_OFN494_n_18414), .b(n_22019), .c(n_657), .d(FE_OFN324_n_4860), .o(n_19439) );
oa22f80 g550795 ( .a(n_18688), .b(FE_OFN154_n_22615), .c(n_1438), .d(FE_OFN355_n_4860), .o(n_19747) );
oa22f80 g550796 ( .a(n_17117), .b(n_22615), .c(n_650), .d(FE_OFN329_n_4860), .o(n_18041) );
oa22f80 g550797 ( .a(n_18846), .b(FE_OFN251_n_4162), .c(n_393), .d(FE_OFN124_n_27449), .o(n_18847) );
oa22f80 g550798 ( .a(n_18413), .b(FE_OFN251_n_4162), .c(n_871), .d(FE_OFN1111_rst), .o(n_19438) );
oa22f80 g550799 ( .a(n_18412), .b(FE_OFN310_n_3069), .c(n_377), .d(FE_OFN1113_rst), .o(n_19437) );
oa22f80 g550800 ( .a(n_17704), .b(FE_OFN150_n_25677), .c(n_215), .d(FE_OFN347_n_4860), .o(n_18573) );
oa22f80 g550801 ( .a(FE_OFN682_n_18155), .b(n_23813), .c(n_342), .d(FE_OFN102_n_27449), .o(n_19151) );
oa22f80 g550802 ( .a(n_18154), .b(FE_OFN235_n_4162), .c(n_888), .d(FE_OFN129_n_27449), .o(n_19150) );
oa22f80 g550803 ( .a(n_16876), .b(FE_OFN199_n_29637), .c(n_415), .d(FE_OFN335_n_4860), .o(n_17797) );
oa22f80 g550804 ( .a(n_18153), .b(FE_OFN314_n_3069), .c(n_763), .d(FE_OFN65_n_27012), .o(n_19149) );
oa22f80 g550805 ( .a(n_18419), .b(FE_OFN314_n_3069), .c(n_1154), .d(FE_OFN124_n_27449), .o(n_19436) );
oa22f80 g550806 ( .a(n_18687), .b(FE_OFN296_n_3069), .c(n_139), .d(n_28362), .o(n_19746) );
na02f80 g550851 ( .a(n_19745), .b(n_19079), .o(n_20485) );
na02f80 g550852 ( .a(n_17491), .b(x_in_24_6), .o(n_18358) );
na02f80 g550853 ( .a(n_19148), .b(n_18516), .o(n_19821) );
na02f80 g550854 ( .a(n_18321), .b(n_17737), .o(n_18980) );
in01f80 g550855 ( .a(n_18571), .o(n_18572) );
na02f80 g550856 ( .a(n_18320), .b(n_17772), .o(n_18571) );
na02f80 g550857 ( .a(n_19435), .b(n_18790), .o(n_20173) );
in01f80 g550858 ( .a(n_18844), .o(n_18845) );
na02f80 g550859 ( .a(n_18570), .b(n_17978), .o(n_18844) );
na02f80 g550860 ( .a(n_18569), .b(n_17997), .o(n_19261) );
na02f80 g550861 ( .a(n_19147), .b(n_18518), .o(n_19824) );
na02f80 g550862 ( .a(n_19146), .b(n_18512), .o(n_19818) );
na02f80 g550863 ( .a(n_19145), .b(n_18510), .o(n_19788) );
na02f80 g550864 ( .a(n_18843), .b(n_18274), .o(n_19481) );
in01f80 g550865 ( .a(n_19743), .o(n_19744) );
na02f80 g550866 ( .a(n_19434), .b(n_18759), .o(n_19743) );
in01f80 g550867 ( .a(n_18567), .o(n_18568) );
no02f80 g550868 ( .a(n_18319), .b(x_in_38_7), .o(n_18567) );
na02f80 g550869 ( .a(n_19144), .b(n_18508), .o(n_19781) );
na02f80 g550870 ( .a(n_19433), .b(n_18786), .o(n_20133) );
na02f80 g550871 ( .a(n_19143), .b(x_in_38_6), .o(n_20165) );
na02f80 g550872 ( .a(n_19132), .b(x_in_28_6), .o(n_20175) );
na02f80 g550873 ( .a(n_19432), .b(n_18768), .o(n_20154) );
na02f80 g550874 ( .a(n_18566), .b(n_18001), .o(n_19258) );
na02f80 g550875 ( .a(n_19431), .b(n_18778), .o(n_20151) );
na02f80 g550876 ( .a(n_19430), .b(n_18776), .o(n_20157) );
in01f80 g550877 ( .a(n_19741), .o(n_19742) );
na02f80 g550878 ( .a(n_19429), .b(n_18783), .o(n_19741) );
in01f80 g550879 ( .a(n_17795), .o(n_17796) );
no02f80 g550880 ( .a(n_17491), .b(x_in_24_6), .o(n_17795) );
no02f80 g550881 ( .a(n_18326), .b(n_18039), .o(n_18040) );
in01f80 g550882 ( .a(n_19427), .o(n_19428) );
no02f80 g550883 ( .a(n_19143), .b(x_in_38_6), .o(n_19427) );
in01f80 g550884 ( .a(n_18841), .o(n_18842) );
na02f80 g550885 ( .a(n_18565), .b(n_17987), .o(n_18841) );
na02f80 g550886 ( .a(n_19426), .b(n_18772), .o(n_20167) );
na02f80 g550887 ( .a(n_18318), .b(n_17766), .o(n_19255) );
na02f80 g550888 ( .a(n_18317), .b(n_17764), .o(n_19250) );
na02f80 g550889 ( .a(n_18840), .b(n_18264), .o(n_19497) );
na02f80 g550890 ( .a(n_19425), .b(n_18780), .o(n_20163) );
na02f80 g550891 ( .a(n_18839), .b(n_18260), .o(n_19796) );
na02f80 g550892 ( .a(n_18334), .b(n_18037), .o(n_18038) );
na02f80 g550893 ( .a(n_18564), .b(n_17994), .o(n_19247) );
na02f80 g550894 ( .a(n_18316), .b(n_17760), .o(n_19244) );
no02f80 g550895 ( .a(n_16635), .b(n_17167), .o(n_18095) );
na02f80 g550896 ( .a(n_19424), .b(n_18774), .o(n_20160) );
na02f80 g550897 ( .a(n_18315), .b(n_17756), .o(n_19239) );
in01f80 g550898 ( .a(n_19141), .o(n_19142) );
na02f80 g550899 ( .a(n_18838), .b(n_18258), .o(n_19141) );
na02f80 g550900 ( .a(n_18314), .b(n_17758), .o(n_18945) );
na02f80 g550901 ( .a(n_18319), .b(x_in_38_7), .o(n_19265) );
na02f80 g550902 ( .a(n_18837), .b(n_18253), .o(n_19469) );
na02f80 g550903 ( .a(n_18836), .b(n_18241), .o(n_19494) );
no02f80 g550904 ( .a(n_18834), .b(n_18833), .o(n_18835) );
na02f80 g550905 ( .a(n_18575), .b(n_18833), .o(n_19542) );
na02f80 g550906 ( .a(n_18046), .b(n_17793), .o(n_17794) );
na02f80 g550907 ( .a(n_19140), .b(n_18482), .o(n_19791) );
na02f80 g550908 ( .a(n_18313), .b(x_in_48_2), .o(n_19228) );
in01f80 g550909 ( .a(n_18562), .o(n_18563) );
no02f80 g550910 ( .a(n_18313), .b(x_in_48_2), .o(n_18562) );
na02f80 g550911 ( .a(n_18561), .b(n_17992), .o(n_19233) );
na02f80 g550912 ( .a(n_18312), .b(n_17768), .o(n_19216) );
na02f80 g550913 ( .a(n_18832), .b(n_18235), .o(n_19463) );
na02f80 g550914 ( .a(n_19423), .b(n_18788), .o(n_20170) );
na02f80 g550915 ( .a(n_18311), .b(n_17754), .o(n_19223) );
na02f80 g550916 ( .a(n_18584), .b(n_18309), .o(n_18310) );
na02f80 g550917 ( .a(n_18560), .b(n_18005), .o(n_19230) );
in01f80 g550918 ( .a(n_19421), .o(n_19422) );
na02f80 g550919 ( .a(n_19139), .b(n_18479), .o(n_19421) );
na02f80 g550920 ( .a(n_18831), .b(x_in_44_5), .o(n_19783) );
in01f80 g550921 ( .a(n_19137), .o(n_19138) );
no02f80 g550922 ( .a(n_18831), .b(x_in_44_5), .o(n_19137) );
na02f80 g550923 ( .a(n_18830), .b(n_18248), .o(n_19466) );
na02f80 g550924 ( .a(n_20108), .b(n_19399), .o(n_20880) );
na02f80 g550925 ( .a(n_18036), .b(x_in_24_5), .o(n_18934) );
in01f80 g550926 ( .a(n_18307), .o(n_18308) );
no02f80 g550927 ( .a(n_18036), .b(x_in_24_5), .o(n_18307) );
no02f80 g550928 ( .a(n_18327), .b(n_18034), .o(n_18035) );
na02f80 g550929 ( .a(n_19136), .b(n_18476), .o(n_19785) );
na02f80 g550930 ( .a(n_18559), .b(n_17999), .o(n_19201) );
na02f80 g550931 ( .a(n_18549), .b(x_in_28_7), .o(n_18922) );
in01f80 g550932 ( .a(n_18305), .o(n_18306) );
no02f80 g550933 ( .a(n_18549), .b(x_in_28_7), .o(n_18305) );
na02f80 g550934 ( .a(n_18304), .b(x_in_48_3), .o(n_19209) );
in01f80 g550935 ( .a(n_18557), .o(n_18558) );
no02f80 g550936 ( .a(n_18304), .b(x_in_48_3), .o(n_18557) );
na02f80 g550937 ( .a(n_18303), .b(n_17749), .o(n_19211) );
na02f80 g550938 ( .a(n_18302), .b(n_17747), .o(n_19207) );
na02f80 g550939 ( .a(n_19740), .b(n_19082), .o(n_20482) );
na02f80 g550940 ( .a(n_18556), .b(n_17969), .o(n_19195) );
na02f80 g550941 ( .a(n_19135), .b(n_18505), .o(n_19815) );
na02f80 g550942 ( .a(n_19420), .b(n_18764), .o(n_20138) );
na02f80 g550943 ( .a(n_18555), .b(n_17967), .o(n_19198) );
no02f80 g550944 ( .a(n_17492), .b(n_17167), .o(n_17168) );
na02f80 g550945 ( .a(n_19419), .b(n_18766), .o(n_20141) );
na02f80 g550946 ( .a(n_18829), .b(x_in_44_4), .o(n_19778) );
in01f80 g550947 ( .a(n_19133), .o(n_19134) );
no02f80 g550948 ( .a(n_18829), .b(x_in_44_4), .o(n_19133) );
in01f80 g550949 ( .a(n_19417), .o(n_19418) );
no02f80 g550950 ( .a(n_19132), .b(x_in_28_6), .o(n_19417) );
no02f80 g550951 ( .a(n_16886), .b(n_16639), .o(n_16640) );
no02f80 g550952 ( .a(n_17165), .b(n_17164), .o(n_17166) );
na02f80 g550953 ( .a(n_17800), .b(n_17489), .o(n_17490) );
no02f80 g550954 ( .a(n_18827), .b(n_18826), .o(n_18828) );
na02f80 g550955 ( .a(n_18554), .b(n_18826), .o(n_19867) );
no02f80 g550956 ( .a(n_17933), .b(n_18552), .o(n_19529) );
no02f80 g550957 ( .a(n_18851), .b(n_18552), .o(n_18553) );
na02f80 g550958 ( .a(n_17116), .b(n_17792), .o(n_18666) );
na02f80 g550959 ( .a(n_17491), .b(n_17792), .o(n_17488) );
no02f80 g550960 ( .a(n_18831), .b(n_18825), .o(n_19474) );
na02f80 g550961 ( .a(n_18846), .b(n_18825), .o(n_18551) );
no02f80 g550962 ( .a(n_19130), .b(n_19129), .o(n_19131) );
no02f80 g550963 ( .a(n_18823), .b(n_18822), .o(n_18824) );
no02f80 g550964 ( .a(n_19738), .b(n_19737), .o(n_19739) );
no02f80 g550965 ( .a(n_19415), .b(n_19414), .o(n_19416) );
na02f80 g550966 ( .a(n_18549), .b(n_18548), .o(n_18550) );
na02f80 g550967 ( .a(n_17705), .b(n_18548), .o(n_19306) );
no02f80 g550968 ( .a(n_18044), .b(n_17790), .o(n_17791) );
no02f80 g550969 ( .a(n_18319), .b(n_18547), .o(n_19303) );
na02f80 g550970 ( .a(n_18545), .b(n_18547), .o(n_18546) );
no02f80 g550971 ( .a(n_18543), .b(n_18542), .o(n_18544) );
na02f80 g550972 ( .a(n_18301), .b(n_17626), .o(n_18871) );
na02f80 g550973 ( .a(n_18301), .b(n_18032), .o(n_18033) );
in01f80 g550974 ( .a(n_18031), .o(n_18658) );
na02f80 g550975 ( .a(n_17789), .b(n_18028), .o(n_18031) );
na02f80 g550976 ( .a(FE_OFN672_n_17494), .b(n_17162), .o(n_17163) );
no02f80 g550977 ( .a(n_18849), .b(n_18540), .o(n_18541) );
no02f80 g550978 ( .a(n_17930), .b(n_18540), .o(n_19525) );
in01f80 g550979 ( .a(n_19875), .o(n_18821) );
oa12f80 g550980 ( .a(n_17988), .b(n_17415), .c(n_17506), .o(n_19875) );
no02f80 g550981 ( .a(n_18029), .b(n_18028), .o(n_18030) );
in01f80 g550982 ( .a(n_19413), .o(n_20515) );
oa12f80 g550983 ( .a(n_17412), .b(n_19125), .c(n_16842), .o(n_19413) );
ao12f80 g550984 ( .a(n_15567), .b(n_17788), .c(n_16264), .o(n_18657) );
ao12f80 g550985 ( .a(n_13667), .b(n_17787), .c(n_14787), .o(n_18656) );
oa12f80 g550986 ( .a(n_15551), .b(n_17161), .c(n_16265), .o(n_18091) );
oa12f80 g550987 ( .a(n_14634), .b(n_17786), .c(n_15345), .o(n_18655) );
oa12f80 g550988 ( .a(n_14784), .b(n_17487), .c(n_15426), .o(n_18389) );
in01f80 g550989 ( .a(n_18820), .o(n_19854) );
oa12f80 g550990 ( .a(n_17698), .b(n_18539), .c(n_17072), .o(n_18820) );
oa12f80 g550991 ( .a(n_14757), .b(n_17486), .c(n_15405), .o(n_18387) );
oa12f80 g550992 ( .a(n_14737), .b(n_17485), .c(n_15395), .o(n_18386) );
ao12f80 g550993 ( .a(n_14376), .b(n_17484), .c(n_15140), .o(n_18385) );
oa12f80 g550994 ( .a(n_14709), .b(n_17483), .c(n_15383), .o(n_18384) );
oa12f80 g550995 ( .a(n_14683), .b(n_17482), .c(n_15365), .o(n_18383) );
ao12f80 g550996 ( .a(n_13148), .b(n_17785), .c(n_14319), .o(n_18654) );
in01f80 g550997 ( .a(n_18300), .o(n_19292) );
ao12f80 g550998 ( .a(n_12300), .b(n_18023), .c(n_12952), .o(n_18300) );
in01f80 g550999 ( .a(n_19128), .o(n_20199) );
oa12f80 g551000 ( .a(n_18399), .b(n_18819), .c(n_17822), .o(n_19128) );
oa12f80 g551001 ( .a(n_15509), .b(n_18299), .c(n_16253), .o(n_19301) );
in01f80 g551002 ( .a(n_18298), .o(n_19289) );
ao12f80 g551003 ( .a(n_11014), .b(n_18022), .c(n_12134), .o(n_18298) );
in01f80 g551004 ( .a(n_18818), .o(n_19848) );
oa12f80 g551005 ( .a(n_17911), .b(n_18538), .c(n_17329), .o(n_18818) );
ao12f80 g551006 ( .a(n_11487), .b(n_17481), .c(n_12475), .o(n_18382) );
oa12f80 g551007 ( .a(n_16095), .b(n_18297), .c(n_16683), .o(n_19300) );
ao12f80 g551008 ( .a(n_11432), .b(n_17480), .c(n_12438), .o(n_18388) );
ao12f80 g551009 ( .a(n_13868), .b(n_17479), .c(n_14918), .o(n_18381) );
ao12f80 g551010 ( .a(n_14697), .b(n_17784), .c(n_15370), .o(n_18653) );
oa12f80 g551011 ( .a(n_11499), .b(n_17160), .c(n_12486), .o(n_18090) );
ao12f80 g551012 ( .a(n_14343), .b(n_17478), .c(n_15129), .o(n_18380) );
ao12f80 g551013 ( .a(n_15484), .b(n_18027), .c(n_16245), .o(n_19001) );
oa12f80 g551014 ( .a(n_8269), .b(n_17783), .c(n_9464), .o(n_18652) );
oa12f80 g551015 ( .a(n_14657), .b(n_18296), .c(n_15351), .o(n_19299) );
ao12f80 g551016 ( .a(n_14300), .b(n_17782), .c(n_15111), .o(n_18651) );
oa12f80 g551017 ( .a(n_13203), .b(n_17477), .c(n_14413), .o(n_18379) );
ao12f80 g551018 ( .a(n_13178), .b(n_18295), .c(n_14369), .o(n_19298) );
oa12f80 g551019 ( .a(n_14440), .b(n_17476), .c(n_15107), .o(n_18378) );
ao12f80 g551020 ( .a(n_13273), .b(n_18025), .c(n_14486), .o(n_19000) );
oa12f80 g551021 ( .a(n_14411), .b(n_17781), .c(n_15153), .o(n_18650) );
oa12f80 g551022 ( .a(n_10759), .b(n_17159), .c(n_11792), .o(n_18089) );
ao12f80 g551023 ( .a(n_14253), .b(n_17475), .c(n_15095), .o(n_18377) );
ao12f80 g551024 ( .a(n_14246), .b(n_17474), .c(n_15093), .o(n_18376) );
ao12f80 g551025 ( .a(n_12272), .b(n_17780), .c(n_12489), .o(n_18649) );
ao12f80 g551026 ( .a(n_15518), .b(n_17473), .c(n_16256), .o(n_18375) );
ao12f80 g551027 ( .a(n_14234), .b(n_17472), .c(n_15172), .o(n_18374) );
oa12f80 g551028 ( .a(n_13955), .b(n_17471), .c(n_14931), .o(n_18373) );
ao12f80 g551029 ( .a(n_10671), .b(n_17470), .c(n_12015), .o(n_18372) );
in01f80 g551030 ( .a(n_17158), .o(n_18087) );
oa22f80 g551031 ( .a(n_16638), .b(n_5104), .c(n_15990), .d(n_16637), .o(n_17158) );
oa12f80 g551032 ( .a(n_8276), .b(n_17469), .c(n_9466), .o(n_18371) );
ao12f80 g551033 ( .a(n_18190), .b(n_18189), .c(n_18188), .o(n_18817) );
oa12f80 g551034 ( .a(n_17941), .b(n_17940), .c(n_17957), .o(n_19274) );
ao12f80 g551035 ( .a(n_19077), .b(n_19076), .c(n_19075), .o(n_19736) );
ao12f80 g551036 ( .a(n_18756), .b(n_18755), .c(n_18754), .o(n_19412) );
oa12f80 g551037 ( .a(n_17952), .b(n_17951), .c(n_17956), .o(n_19266) );
ao12f80 g551038 ( .a(n_18463), .b(n_18462), .c(n_18461), .o(n_19127) );
ao12f80 g551039 ( .a(n_18270), .b(n_18269), .c(n_18268), .o(n_18816) );
ao12f80 g551040 ( .a(n_18753), .b(n_18752), .c(n_18751), .o(n_19411) );
ao22s80 g551041 ( .a(n_19125), .b(n_17688), .c(n_18108), .d(n_17687), .o(n_19126) );
oa12f80 g551042 ( .a(n_17729), .b(n_17728), .c(n_17730), .o(n_18978) );
in01f80 g551043 ( .a(n_18912), .o(n_18638) );
ao12f80 g551044 ( .a(n_17157), .b(n_17487), .c(n_17156), .o(n_18912) );
ao12f80 g551045 ( .a(n_18008), .b(n_18007), .c(n_18006), .o(n_18537) );
ao12f80 g551046 ( .a(n_19074), .b(n_19073), .c(n_19072), .o(n_19735) );
in01f80 g551047 ( .a(n_18644), .o(n_18294) );
oa12f80 g551048 ( .a(n_17468), .b(n_17788), .c(n_17467), .o(n_18644) );
ao12f80 g551049 ( .a(n_19071), .b(n_19070), .c(n_19069), .o(n_19734) );
oa12f80 g551050 ( .a(n_17431), .b(n_17460), .c(n_17723), .o(n_18626) );
ao12f80 g551051 ( .a(n_18750), .b(n_18749), .c(n_18748), .o(n_19410) );
oa12f80 g551052 ( .a(n_17442), .b(n_17459), .c(n_17724), .o(n_18643) );
in01f80 g551053 ( .a(FE_OFN1059_n_18610), .o(n_18888) );
ao12f80 g551054 ( .a(n_17466), .b(n_17787), .c(n_17465), .o(n_18610) );
ao12f80 g551055 ( .a(n_18744), .b(n_18743), .c(n_18742), .o(n_19409) );
ao12f80 g551056 ( .a(n_18202), .b(n_18201), .c(n_18200), .o(n_18815) );
oa12f80 g551057 ( .a(n_17949), .b(n_17948), .c(n_17954), .o(n_19227) );
ao12f80 g551058 ( .a(n_18457), .b(n_18456), .c(n_18455), .o(n_19124) );
oa12f80 g551059 ( .a(n_17443), .b(n_17456), .c(n_17722), .o(n_18642) );
ao12f80 g551060 ( .a(n_18747), .b(n_18746), .c(n_18745), .o(n_19408) );
oa12f80 g551061 ( .a(n_18180), .b(n_18179), .c(n_18178), .o(n_19505) );
ao12f80 g551062 ( .a(n_18499), .b(n_18498), .c(n_18497), .o(n_19123) );
ao12f80 g551063 ( .a(n_18741), .b(n_18740), .c(n_18739), .o(n_19407) );
oa12f80 g551064 ( .a(n_18224), .b(n_18223), .c(n_18222), .o(n_19501) );
in01f80 g551065 ( .a(n_18885), .o(n_18641) );
ao12f80 g551066 ( .a(n_17135), .b(n_17476), .c(n_17134), .o(n_18885) );
in01f80 g551067 ( .a(n_18863), .o(n_18363) );
ao12f80 g551068 ( .a(n_16885), .b(n_17161), .c(n_16884), .o(n_18863) );
in01f80 g551069 ( .a(n_18908), .o(n_18964) );
ao12f80 g551070 ( .a(n_17464), .b(n_17786), .c(n_17463), .o(n_18908) );
ao12f80 g551071 ( .a(n_18735), .b(n_18734), .c(n_18733), .o(n_19406) );
ao12f80 g551072 ( .a(n_18199), .b(n_18198), .c(n_18197), .o(n_18814) );
oa12f80 g551073 ( .a(n_18233), .b(n_18232), .c(n_18231), .o(n_19486) );
ao12f80 g551074 ( .a(n_19103), .b(n_19102), .c(n_19101), .o(n_19733) );
ao12f80 g551075 ( .a(n_18738), .b(n_18737), .c(n_18736), .o(n_19405) );
oa12f80 g551076 ( .a(n_18220), .b(n_18219), .c(n_18218), .o(n_19500) );
ao12f80 g551077 ( .a(n_18732), .b(n_18731), .c(n_18730), .o(n_19404) );
oa12f80 g551078 ( .a(n_18217), .b(n_18216), .c(n_18221), .o(n_19492) );
ao12f80 g551079 ( .a(n_18729), .b(n_18728), .c(n_18727), .o(n_19403) );
oa12f80 g551080 ( .a(n_18230), .b(n_18229), .c(n_18228), .o(n_19499) );
ao12f80 g551081 ( .a(n_18726), .b(n_18725), .c(n_18724), .o(n_19402) );
ao12f80 g551082 ( .a(n_17721), .b(n_18011), .c(n_17720), .o(n_18293) );
ao12f80 g551083 ( .a(n_19100), .b(n_19099), .c(n_19098), .o(n_19732) );
ao12f80 g551084 ( .a(n_18723), .b(n_18722), .c(n_18721), .o(n_19401) );
in01f80 g551085 ( .a(n_18328), .o(n_18586) );
ao12f80 g551086 ( .a(n_17137), .b(n_17477), .c(n_17136), .o(n_18328) );
in01f80 g551087 ( .a(n_18905), .o(n_18637) );
ao12f80 g551088 ( .a(n_17153), .b(n_17486), .c(n_17152), .o(n_18905) );
ao12f80 g551089 ( .a(n_19097), .b(n_19096), .c(n_19095), .o(n_19731) );
in01f80 g551090 ( .a(n_18882), .o(n_18958) );
ao12f80 g551091 ( .a(n_17449), .b(n_17781), .c(n_17448), .o(n_18882) );
in01f80 g551092 ( .a(n_18902), .o(n_18636) );
ao12f80 g551093 ( .a(n_17151), .b(n_17485), .c(n_17150), .o(n_18902) );
ao12f80 g551094 ( .a(n_19094), .b(n_19093), .c(n_19092), .o(n_19730) );
ao12f80 g551095 ( .a(n_18196), .b(n_18195), .c(n_18194), .o(n_18813) );
in01f80 g551096 ( .a(n_18873), .o(n_18635) );
ao12f80 g551097 ( .a(n_17149), .b(n_17484), .c(n_17148), .o(n_18873) );
in01f80 g551098 ( .a(n_18812), .o(n_19835) );
oa12f80 g551099 ( .a(n_17963), .b(n_18295), .c(n_17962), .o(n_18812) );
ao12f80 g551100 ( .a(n_18489), .b(n_18488), .c(n_18487), .o(n_19122) );
ao12f80 g551101 ( .a(n_18486), .b(n_18485), .c(n_18484), .o(n_19121) );
in01f80 g551102 ( .a(n_18899), .o(n_18634) );
ao12f80 g551103 ( .a(n_17147), .b(n_17483), .c(n_17146), .o(n_18899) );
in01f80 g551104 ( .a(n_18343), .o(n_18633) );
ao12f80 g551105 ( .a(n_17139), .b(n_17478), .c(n_17138), .o(n_18343) );
ao12f80 g551106 ( .a(n_19091), .b(n_19090), .c(n_19089), .o(n_19729) );
ao12f80 g551107 ( .a(n_18454), .b(n_18453), .c(n_18452), .o(n_19120) );
in01f80 g551108 ( .a(n_18892), .o(n_18949) );
ao12f80 g551109 ( .a(n_17455), .b(n_17784), .c(n_17454), .o(n_18892) );
in01f80 g551110 ( .a(n_18896), .o(n_18632) );
ao12f80 g551111 ( .a(n_17145), .b(n_17482), .c(n_17144), .o(n_18896) );
ao12f80 g551112 ( .a(n_19088), .b(n_19087), .c(n_19086), .o(n_19728) );
in01f80 g551113 ( .a(n_18292), .o(n_19282) );
oa12f80 g551114 ( .a(n_17447), .b(n_17780), .c(n_17446), .o(n_18292) );
ao12f80 g551115 ( .a(n_18256), .b(n_18255), .c(n_18254), .o(n_18811) );
oa12f80 g551116 ( .a(n_18184), .b(n_18246), .c(n_18433), .o(n_19491) );
ao12f80 g551117 ( .a(n_18208), .b(n_18207), .c(n_18206), .o(n_18810) );
ao12f80 g551118 ( .a(n_17439), .b(FE_OFN722_n_17438), .c(n_17437), .o(n_18026) );
oa12f80 g551119 ( .a(n_17947), .b(n_18183), .c(n_17946), .o(n_19235) );
ao12f80 g551120 ( .a(n_18451), .b(n_18450), .c(n_18449), .o(n_19119) );
in01f80 g551121 ( .a(n_18341), .o(n_18631) );
ao12f80 g551122 ( .a(n_17125), .b(n_17471), .c(n_17124), .o(n_18341) );
in01f80 g551123 ( .a(n_18869), .o(n_18929) );
ao22s80 g551124 ( .a(n_18025), .b(n_14816), .c(n_17106), .d(n_14817), .o(n_18869) );
ao12f80 g551125 ( .a(n_19085), .b(n_19084), .c(n_19083), .o(n_19727) );
ao12f80 g551126 ( .a(n_18493), .b(n_18492), .c(n_18491), .o(n_19118) );
ao12f80 g551127 ( .a(n_18205), .b(n_18204), .c(n_18203), .o(n_18809) );
ao12f80 g551128 ( .a(n_17719), .b(n_17718), .c(n_17717), .o(n_18291) );
in01f80 g551129 ( .a(n_18603), .o(n_18024) );
oa12f80 g551130 ( .a(n_17121), .b(n_17469), .c(n_17120), .o(n_18603) );
in01f80 g551131 ( .a(n_18614), .o(n_18919) );
ao22s80 g551132 ( .a(n_17102), .b(n_13503), .c(n_18023), .d(n_13502), .o(n_18614) );
oa12f80 g551133 ( .a(n_17732), .b(n_17731), .c(n_17733), .o(n_18938) );
in01f80 g551134 ( .a(n_18608), .o(n_18290) );
oa12f80 g551135 ( .a(n_17462), .b(n_17785), .c(n_17461), .o(n_18608) );
ao12f80 g551136 ( .a(n_17985), .b(n_17984), .c(n_17983), .o(n_18536) );
ao22s80 g551137 ( .a(n_18685), .b(n_18819), .c(n_18684), .d(n_17864), .o(n_19726) );
in01f80 g551138 ( .a(n_19471), .o(n_19473) );
oa12f80 g551139 ( .a(n_17965), .b(n_18296), .c(n_17964), .o(n_19471) );
in01f80 g551140 ( .a(n_18599), .o(n_18943) );
ao12f80 g551141 ( .a(n_17451), .b(n_17782), .c(n_17450), .o(n_18599) );
oa12f80 g551142 ( .a(n_17714), .b(n_17769), .c(n_17944), .o(n_18937) );
in01f80 g551143 ( .a(n_19186), .o(n_18629) );
ao12f80 g551144 ( .a(n_17129), .b(n_17473), .c(n_17128), .o(n_19186) );
ao12f80 g551145 ( .a(n_18460), .b(n_18459), .c(n_18458), .o(n_19117) );
na03f80 g551146 ( .a(n_12316), .b(n_16878), .c(n_10698), .o(n_17779) );
in01f80 g551147 ( .a(n_18047), .o(n_18332) );
ao12f80 g551148 ( .a(n_16883), .b(n_17160), .c(n_16882), .o(n_18047) );
in01f80 g551149 ( .a(n_18335), .o(n_18630) );
ao12f80 g551150 ( .a(n_17141), .b(n_17479), .c(n_17140), .o(n_18335) );
ao12f80 g551151 ( .a(n_18193), .b(n_18192), .c(n_18191), .o(n_18808) );
ao12f80 g551152 ( .a(n_17981), .b(n_17980), .c(n_17979), .o(n_18535) );
ao22s80 g551153 ( .a(n_17909), .b(n_18539), .c(n_17908), .d(n_17623), .o(n_18807) );
in01f80 g551154 ( .a(n_18595), .o(n_18961) );
ao22s80 g551155 ( .a(n_17101), .b(n_12560), .c(n_18022), .d(n_12559), .o(n_18595) );
oa12f80 g551156 ( .a(n_17436), .b(n_17435), .c(n_17713), .o(n_18628) );
in01f80 g551157 ( .a(n_18609), .o(n_18627) );
ao12f80 g551158 ( .a(n_17133), .b(n_17475), .c(n_17132), .o(n_18609) );
ao12f80 g551159 ( .a(n_17434), .b(FE_OFN1017_n_17433), .c(n_17432), .o(n_18021) );
in01f80 g551160 ( .a(n_18329), .o(n_18591) );
ao12f80 g551161 ( .a(n_17123), .b(n_17470), .c(n_17122), .o(n_18329) );
ao22s80 g551162 ( .a(n_18140), .b(n_18538), .c(n_18139), .d(n_17625), .o(n_19116) );
oa12f80 g551163 ( .a(n_18226), .b(n_18225), .c(n_18227), .o(n_19502) );
ao12f80 g551164 ( .a(n_18244), .b(n_18243), .c(n_18242), .o(n_18806) );
in01f80 g551165 ( .a(n_19271), .o(n_18805) );
oa12f80 g551166 ( .a(n_17976), .b(n_18299), .c(n_17975), .o(n_19271) );
ao12f80 g551167 ( .a(n_17445), .b(n_17777), .c(n_17444), .o(n_18020) );
in01f80 g551168 ( .a(n_18050), .o(n_18346) );
ao12f80 g551169 ( .a(n_16881), .b(n_17159), .c(n_16880), .o(n_18050) );
in01f80 g551170 ( .a(n_18597), .o(n_18625) );
ao12f80 g551171 ( .a(n_17131), .b(n_17474), .c(n_17130), .o(n_18597) );
in01f80 g551172 ( .a(n_18289), .o(n_19278) );
oa12f80 g551173 ( .a(n_17453), .b(n_17783), .c(n_17452), .o(n_18289) );
in01f80 g551174 ( .a(n_19773), .o(n_19485) );
ao12f80 g551175 ( .a(n_17974), .b(n_18297), .c(n_17973), .o(n_19773) );
oa12f80 g551176 ( .a(n_18445), .b(n_18490), .c(n_18710), .o(n_19779) );
ao12f80 g551177 ( .a(n_18239), .b(n_18238), .c(n_18237), .o(n_18804) );
ao12f80 g551178 ( .a(n_17744), .b(n_17743), .c(n_17742), .o(n_18288) );
in01f80 g551179 ( .a(n_18019), .o(n_18988) );
oa12f80 g551180 ( .a(n_17143), .b(n_17480), .c(n_17142), .o(n_18019) );
oa12f80 g551181 ( .a(n_18709), .b(n_18708), .c(n_18707), .o(n_20143) );
in01f80 g551182 ( .a(n_18877), .o(n_18622) );
ao12f80 g551183 ( .a(n_17127), .b(n_17472), .c(n_17126), .o(n_18877) );
ao12f80 g551184 ( .a(n_17741), .b(n_17740), .c(n_17739), .o(n_18287) );
oa12f80 g551185 ( .a(n_17726), .b(n_17725), .c(n_17727), .o(n_18975) );
oa12f80 g551186 ( .a(n_17942), .b(n_18003), .c(n_18177), .o(n_19203) );
ao12f80 g551187 ( .a(n_18211), .b(n_18210), .c(n_18209), .o(n_18803) );
ao12f80 g551188 ( .a(n_17712), .b(n_18015), .c(n_17711), .o(n_18286) );
oa12f80 g551189 ( .a(n_18214), .b(n_18213), .c(n_18215), .o(n_19477) );
ao12f80 g551190 ( .a(n_18467), .b(n_18466), .c(n_18465), .o(n_19115) );
ao12f80 g551191 ( .a(n_18720), .b(n_18719), .c(n_18718), .o(n_19400) );
ao12f80 g551192 ( .a(n_18448), .b(n_18447), .c(n_18446), .o(n_19114) );
ao12f80 g551193 ( .a(n_17959), .b(n_17958), .c(n_17960), .o(n_18534) );
in01f80 g551194 ( .a(n_18018), .o(n_18982) );
oa12f80 g551195 ( .a(n_17155), .b(n_17481), .c(n_17154), .o(n_18018) );
ao12f80 g551196 ( .a(n_18502), .b(n_18501), .c(n_18500), .o(n_19113) );
oa12f80 g551197 ( .a(n_18431), .b(n_18430), .c(n_18429), .o(n_19775) );
in01f80 g551198 ( .a(n_18918), .o(n_18533) );
oa12f80 g551199 ( .a(n_17735), .b(n_18027), .c(n_17734), .o(n_18918) );
oa22f80 g551200 ( .a(n_18107), .b(FE_OFN314_n_3069), .c(n_1789), .d(rst), .o(n_19112) );
oa22f80 g551201 ( .a(n_17616), .b(FE_OFN411_n_28303), .c(n_934), .d(FE_OFN1182_rst), .o(n_18532) );
oa22f80 g551202 ( .a(n_18106), .b(FE_OFN313_n_3069), .c(n_1834), .d(FE_OFN361_n_4860), .o(n_19111) );
oa22f80 g551203 ( .a(n_17855), .b(FE_OFN264_n_4280), .c(n_1336), .d(FE_OFN1110_rst), .o(n_18802) );
oa22f80 g551204 ( .a(n_17861), .b(FE_OFN406_n_28303), .c(n_1725), .d(FE_OFN1112_rst), .o(n_18801) );
oa22f80 g551205 ( .a(FE_OFN598_n_17615), .b(n_23291), .c(n_928), .d(FE_OFN63_n_27012), .o(n_18531) );
oa22f80 g551206 ( .a(n_17390), .b(FE_OFN198_n_29637), .c(n_59), .d(FE_OFN65_n_27012), .o(n_18285) );
oa22f80 g551207 ( .a(n_18105), .b(FE_OFN292_n_3069), .c(n_1567), .d(FE_OFN1115_rst), .o(n_19110) );
oa22f80 g551208 ( .a(n_17613), .b(FE_OFN1160_n_26184), .c(n_660), .d(FE_OFN65_n_27012), .o(n_18530) );
oa22f80 g551209 ( .a(n_17606), .b(n_26184), .c(n_1414), .d(FE_OFN128_n_27449), .o(n_18529) );
oa22f80 g551210 ( .a(n_17612), .b(FE_OFN239_n_4162), .c(n_151), .d(FE_OFN74_n_27012), .o(n_18528) );
oa22f80 g551211 ( .a(n_17607), .b(n_28303), .c(n_936), .d(FE_OFN1117_rst), .o(n_18527) );
oa22f80 g551212 ( .a(n_17089), .b(n_29698), .c(n_375), .d(FE_OFN1118_rst), .o(n_18017) );
oa22f80 g551213 ( .a(n_17605), .b(FE_OFN414_n_28303), .c(n_1396), .d(FE_OFN115_n_27449), .o(n_18526) );
oa22f80 g551214 ( .a(n_17777), .b(FE_OFN267_n_4280), .c(n_1883), .d(FE_OFN92_n_27449), .o(n_17778) );
oa22f80 g551215 ( .a(n_18015), .b(FE_OFN187_n_29496), .c(n_438), .d(FE_OFN135_n_27449), .o(n_18016) );
oa22f80 g551216 ( .a(n_17458), .b(FE_OFN406_n_28303), .c(n_1521), .d(FE_OFN99_n_27449), .o(n_17776) );
oa22f80 g551217 ( .a(n_17611), .b(FE_OFN409_n_28303), .c(n_863), .d(FE_OFN355_n_4860), .o(n_18524) );
oa22f80 g551218 ( .a(n_17859), .b(FE_OFN186_n_29496), .c(n_1605), .d(FE_OFN189_n_28362), .o(n_18800) );
oa22f80 g551219 ( .a(n_18212), .b(FE_OFN254_n_4280), .c(n_1768), .d(FE_OFN77_n_27012), .o(n_18523) );
oa22f80 g551220 ( .a(n_17858), .b(FE_OFN244_n_4162), .c(n_956), .d(FE_OFN139_n_27449), .o(n_18799) );
oa22f80 g551221 ( .a(n_17857), .b(FE_OFN187_n_29496), .c(n_401), .d(FE_OFN350_n_4860), .o(n_18798) );
oa22f80 g551222 ( .a(n_18104), .b(FE_OFN265_n_4280), .c(n_356), .d(FE_OFN129_n_27449), .o(n_19109) );
oa22f80 g551223 ( .a(n_17389), .b(FE_OFN410_n_28303), .c(n_925), .d(FE_OFN130_n_27449), .o(n_18284) );
oa22f80 g551224 ( .a(n_17610), .b(FE_OFN300_n_3069), .c(n_1385), .d(FE_OFN324_n_4860), .o(n_18522) );
oa22f80 g551225 ( .a(FE_OFN602_n_17761), .b(n_29698), .c(n_1086), .d(FE_OFN336_n_4860), .o(n_18014) );
oa22f80 g551226 ( .a(n_17856), .b(FE_OFN214_n_29687), .c(n_673), .d(FE_OFN361_n_4860), .o(n_18797) );
oa22f80 g551227 ( .a(n_17090), .b(FE_OFN258_n_4280), .c(n_461), .d(FE_OFN358_n_4860), .o(n_18013) );
oa22f80 g551228 ( .a(FE_OFN584_n_18103), .b(n_23291), .c(n_839), .d(FE_OFN63_n_27012), .o(n_19108) );
oa22f80 g551229 ( .a(n_17387), .b(FE_OFN309_n_3069), .c(n_1426), .d(FE_OFN134_n_27449), .o(n_18283) );
oa22f80 g551230 ( .a(n_17854), .b(FE_OFN198_n_29637), .c(n_901), .d(FE_OFN352_n_4860), .o(n_18796) );
oa22f80 g551231 ( .a(n_18011), .b(FE_OFN269_n_4280), .c(n_982), .d(FE_OFN1114_rst), .o(n_18012) );
oa22f80 g551232 ( .a(n_17609), .b(FE_OFN235_n_4162), .c(n_824), .d(FE_OFN1114_rst), .o(n_18520) );
oa22f80 g551233 ( .a(n_17608), .b(FE_OFN295_n_3069), .c(n_58), .d(FE_OFN1112_rst), .o(n_18519) );
oa22f80 g551234 ( .a(n_17384), .b(FE_OFN258_n_4280), .c(n_1916), .d(FE_OFN358_n_4860), .o(n_18282) );
oa22f80 g551235 ( .a(n_16850), .b(n_23813), .c(n_1141), .d(FE_OFN102_n_27449), .o(n_17775) );
oa22f80 g551236 ( .a(n_17383), .b(FE_OFN314_n_3069), .c(n_1456), .d(FE_OFN124_n_27449), .o(n_18281) );
oa22f80 g551237 ( .a(n_17382), .b(FE_OFN314_n_3069), .c(n_1721), .d(FE_OFN98_n_27449), .o(n_18280) );
oa22f80 g551238 ( .a(n_17381), .b(FE_OFN310_n_3069), .c(n_1933), .d(FE_OFN1143_n_27012), .o(n_18279) );
oa22f80 g551239 ( .a(n_17852), .b(FE_OFN152_n_22615), .c(n_261), .d(FE_OFN1119_rst), .o(n_18795) );
oa22f80 g551240 ( .a(n_17380), .b(FE_OFN158_n_28014), .c(n_1564), .d(FE_OFN1121_rst), .o(n_18278) );
oa22f80 g551241 ( .a(n_17716), .b(FE_OFN297_n_3069), .c(n_1793), .d(FE_OFN1121_rst), .o(n_17774) );
oa22f80 g551242 ( .a(n_17085), .b(n_29698), .c(n_574), .d(FE_OFN89_n_27449), .o(n_18010) );
oa22f80 g551243 ( .a(n_17961), .b(FE_OFN149_n_25677), .c(n_1551), .d(FE_OFN336_n_4860), .o(n_18009) );
oa22f80 g551244 ( .a(n_17851), .b(n_29698), .c(n_577), .d(FE_OFN56_n_27012), .o(n_18794) );
oa22f80 g551245 ( .a(FE_OFN769_n_17379), .b(n_28303), .c(n_586), .d(n_25680), .o(n_18277) );
oa22f80 g551246 ( .a(n_17850), .b(FE_OFN247_n_4162), .c(n_1627), .d(FE_OFN69_n_27012), .o(n_18793) );
oa22f80 g551247 ( .a(FE_OFN624_n_17378), .b(n_28608), .c(n_539), .d(n_27709), .o(n_18276) );
oa22f80 g551248 ( .a(n_17849), .b(n_28303), .c(n_813), .d(FE_OFN1109_rst), .o(n_18792) );
oa22f80 g551249 ( .a(n_17377), .b(FE_OFN314_n_3069), .c(n_1680), .d(FE_OFN124_n_27449), .o(n_18275) );
oa22f80 g551250 ( .a(n_17848), .b(n_29496), .c(n_1646), .d(FE_OFN1108_rst), .o(n_18791) );
oa22f80 g551251 ( .a(n_17457), .b(FE_OFN311_n_3069), .c(n_1303), .d(FE_OFN134_n_27449), .o(n_17773) );
in01f80 g551300 ( .a(n_18273), .o(n_18274) );
no02f80 g551301 ( .a(n_18430), .b(x_in_60_3), .o(n_18273) );
na02f80 g551302 ( .a(n_18266), .b(x_in_42_3), .o(n_19145) );
na02f80 g551303 ( .a(n_18272), .b(x_in_2_3), .o(n_19147) );
in01f80 g551304 ( .a(n_18517), .o(n_18518) );
no02f80 g551305 ( .a(n_18272), .b(x_in_2_3), .o(n_18517) );
na02f80 g551306 ( .a(n_17752), .b(x_in_56_5), .o(n_18565) );
in01f80 g551307 ( .a(n_18515), .o(n_18516) );
no02f80 g551308 ( .a(n_18271), .b(x_in_34_3), .o(n_18515) );
na02f80 g551309 ( .a(n_18271), .b(x_in_34_3), .o(n_19148) );
no02f80 g551310 ( .a(n_17487), .b(n_17156), .o(n_17157) );
no02f80 g551311 ( .a(n_18269), .b(n_18268), .o(n_18270) );
in01f80 g551312 ( .a(n_17771), .o(n_17772) );
no02f80 g551313 ( .a(n_17731), .b(x_in_8_6), .o(n_17771) );
na02f80 g551314 ( .a(n_17481), .b(n_17154), .o(n_17155) );
na02f80 g551315 ( .a(n_18514), .b(x_in_18_3), .o(n_19435) );
in01f80 g551316 ( .a(n_18789), .o(n_18790) );
no02f80 g551317 ( .a(n_18514), .b(x_in_18_3), .o(n_18789) );
no02f80 g551318 ( .a(n_18007), .b(n_18006), .o(n_18008) );
na02f80 g551319 ( .a(n_18513), .b(x_in_50_3), .o(n_19423) );
in01f80 g551320 ( .a(n_18787), .o(n_18788) );
no02f80 g551321 ( .a(n_18513), .b(x_in_50_3), .o(n_18787) );
na02f80 g551322 ( .a(n_17788), .b(n_17467), .o(n_17468) );
na02f80 g551323 ( .a(n_18179), .b(x_in_6_3), .o(n_18560) );
in01f80 g551324 ( .a(n_18004), .o(n_18005) );
no02f80 g551325 ( .a(n_18179), .b(x_in_6_3), .o(n_18004) );
na02f80 g551326 ( .a(n_18267), .b(x_in_10_3), .o(n_19146) );
in01f80 g551327 ( .a(n_18511), .o(n_18512) );
no02f80 g551328 ( .a(n_18267), .b(x_in_10_3), .o(n_18511) );
in01f80 g551329 ( .a(n_18509), .o(n_18510) );
no02f80 g551330 ( .a(n_18266), .b(x_in_42_3), .o(n_18509) );
no02f80 g551331 ( .a(n_17787), .b(n_17465), .o(n_17466) );
na02f80 g551332 ( .a(n_18265), .b(x_in_58_3), .o(n_19144) );
in01f80 g551333 ( .a(n_18507), .o(n_18508) );
no02f80 g551334 ( .a(n_18265), .b(x_in_58_3), .o(n_18507) );
na02f80 g551335 ( .a(n_18506), .b(x_in_6_2), .o(n_19433) );
in01f80 g551336 ( .a(n_18785), .o(n_18786) );
no02f80 g551337 ( .a(n_18506), .b(x_in_6_2), .o(n_18785) );
in01f80 g551338 ( .a(n_18504), .o(n_18505) );
no02f80 g551339 ( .a(n_18251), .b(x_in_26_3), .o(n_18504) );
in01f80 g551340 ( .a(n_18263), .o(n_18264) );
no02f80 g551341 ( .a(n_18003), .b(x_in_52_3), .o(n_18263) );
in01f80 g551342 ( .a(n_19106), .o(n_19107) );
na02f80 g551343 ( .a(n_18784), .b(n_18121), .o(n_19106) );
na02f80 g551344 ( .a(n_18503), .b(x_in_38_5), .o(n_19429) );
in01f80 g551345 ( .a(n_18782), .o(n_18783) );
no02f80 g551346 ( .a(n_18503), .b(x_in_38_5), .o(n_18782) );
in01f80 g551347 ( .a(n_18261), .o(n_18262) );
na02f80 g551348 ( .a(n_18002), .b(n_17419), .o(n_18261) );
no02f80 g551349 ( .a(n_18501), .b(n_18500), .o(n_18502) );
na02f80 g551350 ( .a(n_17731), .b(x_in_8_6), .o(n_18320) );
no02f80 g551351 ( .a(n_18498), .b(n_18497), .o(n_18499) );
in01f80 g551352 ( .a(n_19104), .o(n_19105) );
na02f80 g551353 ( .a(n_18781), .b(n_18136), .o(n_19104) );
na02f80 g551354 ( .a(n_18480), .b(x_in_22_3), .o(n_19432) );
in01f80 g551355 ( .a(n_18779), .o(n_18780) );
no02f80 g551356 ( .a(n_18468), .b(x_in_54_3), .o(n_18779) );
na02f80 g551357 ( .a(n_17770), .b(x_in_2_4), .o(n_18559) );
no02f80 g551358 ( .a(n_17786), .b(n_17463), .o(n_17464) );
no02f80 g551359 ( .a(n_17161), .b(n_16884), .o(n_16885) );
na02f80 g551360 ( .a(n_18003), .b(x_in_52_3), .o(n_18840) );
in01f80 g551361 ( .a(n_18000), .o(n_18001) );
no02f80 g551362 ( .a(n_18225), .b(x_in_22_4), .o(n_18000) );
na02f80 g551363 ( .a(n_17769), .b(x_in_40_3), .o(n_18569) );
na02f80 g551364 ( .a(n_18496), .b(x_in_14_3), .o(n_19431) );
in01f80 g551365 ( .a(n_18777), .o(n_18778) );
no02f80 g551366 ( .a(n_18496), .b(x_in_14_3), .o(n_18777) );
no02f80 g551367 ( .a(n_19102), .b(n_19101), .o(n_19103) );
in01f80 g551368 ( .a(n_17998), .o(n_17999) );
no02f80 g551369 ( .a(n_17770), .b(x_in_2_4), .o(n_17998) );
na02f80 g551370 ( .a(n_18495), .b(x_in_46_3), .o(n_19430) );
in01f80 g551371 ( .a(n_18775), .o(n_18776) );
no02f80 g551372 ( .a(n_18495), .b(x_in_46_3), .o(n_18775) );
na02f80 g551373 ( .a(n_18494), .b(x_in_30_3), .o(n_19424) );
in01f80 g551374 ( .a(n_18773), .o(n_18774) );
no02f80 g551375 ( .a(n_18494), .b(x_in_30_3), .o(n_18773) );
na02f80 g551376 ( .a(n_18223), .b(x_in_54_4), .o(n_18312) );
in01f80 g551377 ( .a(n_17767), .o(n_17768) );
no02f80 g551378 ( .a(n_18223), .b(x_in_54_4), .o(n_17767) );
na02f80 g551379 ( .a(n_18477), .b(x_in_62_3), .o(n_19420) );
in01f80 g551380 ( .a(n_17996), .o(n_17997) );
no02f80 g551381 ( .a(n_17769), .b(x_in_40_3), .o(n_17996) );
no02f80 g551382 ( .a(n_19099), .b(n_19098), .o(n_19100) );
no02f80 g551383 ( .a(n_18492), .b(n_18491), .o(n_18493) );
na02f80 g551384 ( .a(n_18490), .b(x_in_36_3), .o(n_19426) );
in01f80 g551385 ( .a(n_18771), .o(n_18772) );
no02f80 g551386 ( .a(n_18490), .b(x_in_36_3), .o(n_18771) );
no02f80 g551387 ( .a(n_17486), .b(n_17152), .o(n_17153) );
na02f80 g551388 ( .a(n_18232), .b(x_in_14_4), .o(n_18318) );
in01f80 g551389 ( .a(n_17765), .o(n_17766) );
no02f80 g551390 ( .a(n_18232), .b(x_in_14_4), .o(n_17765) );
no02f80 g551391 ( .a(n_19096), .b(n_19095), .o(n_19097) );
na02f80 g551392 ( .a(n_17995), .b(x_in_34_4), .o(n_18839) );
in01f80 g551393 ( .a(n_18259), .o(n_18260) );
no02f80 g551394 ( .a(n_17995), .b(x_in_34_4), .o(n_18259) );
no02f80 g551395 ( .a(n_17485), .b(n_17150), .o(n_17151) );
na02f80 g551396 ( .a(n_18219), .b(x_in_46_4), .o(n_18317) );
in01f80 g551397 ( .a(n_17763), .o(n_17764) );
no02f80 g551398 ( .a(n_18219), .b(x_in_46_4), .o(n_17763) );
no02f80 g551399 ( .a(n_19093), .b(n_19092), .o(n_19094) );
no02f80 g551400 ( .a(n_17484), .b(n_17148), .o(n_17149) );
na02f80 g551401 ( .a(n_17762), .b(x_in_16_4), .o(n_18564) );
in01f80 g551402 ( .a(n_17993), .o(n_17994) );
no02f80 g551403 ( .a(n_17762), .b(x_in_16_4), .o(n_17993) );
no02f80 g551404 ( .a(n_18488), .b(n_18487), .o(n_18489) );
na02f80 g551405 ( .a(FE_OFN602_n_17761), .b(n_18006), .o(n_18976) );
no02f80 g551406 ( .a(n_18485), .b(n_18484), .o(n_18486) );
no02f80 g551407 ( .a(n_17483), .b(n_17146), .o(n_17147) );
na02f80 g551408 ( .a(n_18216), .b(x_in_30_4), .o(n_18316) );
in01f80 g551409 ( .a(n_17759), .o(n_17760) );
no02f80 g551410 ( .a(n_18216), .b(x_in_30_4), .o(n_17759) );
na02f80 g551411 ( .a(n_17728), .b(x_in_18_4), .o(n_18314) );
in01f80 g551412 ( .a(n_17757), .o(n_17758) );
no02f80 g551413 ( .a(n_17728), .b(x_in_18_4), .o(n_17757) );
no02f80 g551414 ( .a(n_19090), .b(n_19089), .o(n_19091) );
na02f80 g551415 ( .a(n_18213), .b(x_in_12_4), .o(n_18561) );
in01f80 g551416 ( .a(n_17991), .o(n_17992) );
no02f80 g551417 ( .a(n_18213), .b(x_in_12_4), .o(n_17991) );
no02f80 g551418 ( .a(n_17482), .b(n_17144), .o(n_17145) );
na02f80 g551419 ( .a(n_18229), .b(x_in_62_4), .o(n_18315) );
in01f80 g551420 ( .a(n_17755), .o(n_17756) );
no02f80 g551421 ( .a(n_18229), .b(x_in_62_4), .o(n_17755) );
no02f80 g551422 ( .a(n_19087), .b(n_19086), .o(n_19088) );
in01f80 g551423 ( .a(n_18769), .o(n_18770) );
na02f80 g551424 ( .a(n_18483), .b(n_17903), .o(n_18769) );
na02f80 g551425 ( .a(n_17990), .b(x_in_0_14), .o(n_18838) );
in01f80 g551426 ( .a(n_18257), .o(n_18258) );
no02f80 g551427 ( .a(n_17990), .b(x_in_0_14), .o(n_18257) );
no02f80 g551428 ( .a(n_18255), .b(n_18254), .o(n_18256) );
na02f80 g551429 ( .a(n_17989), .b(x_in_32_2), .o(n_18837) );
in01f80 g551430 ( .a(n_18252), .o(n_18253) );
no02f80 g551431 ( .a(n_17989), .b(x_in_32_2), .o(n_18252) );
na02f80 g551432 ( .a(n_18251), .b(x_in_26_3), .o(n_19135) );
na02f80 g551433 ( .a(n_18250), .b(x_in_16_3), .o(n_19140) );
in01f80 g551434 ( .a(n_18481), .o(n_18482) );
no02f80 g551435 ( .a(n_18250), .b(x_in_16_3), .o(n_18481) );
na02f80 g551436 ( .a(n_17988), .b(n_17416), .o(n_18543) );
na02f80 g551437 ( .a(n_17725), .b(x_in_50_4), .o(n_18311) );
in01f80 g551438 ( .a(n_17753), .o(n_17754) );
no02f80 g551439 ( .a(n_17725), .b(x_in_50_4), .o(n_17753) );
in01f80 g551440 ( .a(n_18767), .o(n_18768) );
no02f80 g551441 ( .a(n_18480), .b(x_in_22_3), .o(n_18767) );
in01f80 g551442 ( .a(n_18765), .o(n_18766) );
no02f80 g551443 ( .a(n_18471), .b(x_in_12_3), .o(n_18765) );
no02f80 g551444 ( .a(n_19084), .b(n_19083), .o(n_19085) );
in01f80 g551445 ( .a(n_17986), .o(n_17987) );
no02f80 g551446 ( .a(n_17752), .b(x_in_56_5), .o(n_17986) );
na02f80 g551447 ( .a(n_18249), .b(x_in_8_5), .o(n_19139) );
in01f80 g551448 ( .a(n_18478), .o(n_18479) );
no02f80 g551449 ( .a(n_18249), .b(x_in_8_5), .o(n_18478) );
na02f80 g551450 ( .a(n_17785), .b(n_17461), .o(n_17462) );
in01f80 g551451 ( .a(n_18763), .o(n_18764) );
no02f80 g551452 ( .a(n_18477), .b(x_in_62_3), .o(n_18763) );
no02f80 g551453 ( .a(n_17984), .b(n_17983), .o(n_17985) );
na02f80 g551454 ( .a(n_17982), .b(x_in_40_2), .o(n_18830) );
in01f80 g551455 ( .a(n_18247), .o(n_18248) );
no02f80 g551456 ( .a(n_17982), .b(x_in_40_2), .o(n_18247) );
na02f80 g551457 ( .a(n_18246), .b(x_in_32_3), .o(n_19136) );
in01f80 g551458 ( .a(n_18475), .o(n_18476) );
no02f80 g551459 ( .a(n_18246), .b(x_in_32_3), .o(n_18475) );
na02f80 g551460 ( .a(n_19080), .b(x_in_20_2), .o(n_20108) );
no02f80 g551461 ( .a(n_17160), .b(n_16882), .o(n_16883) );
na02f80 g551462 ( .a(n_17751), .b(x_in_26_4), .o(n_18555) );
no02f80 g551463 ( .a(n_17980), .b(n_17979), .o(n_17981) );
in01f80 g551464 ( .a(n_18761), .o(n_18762) );
na02f80 g551465 ( .a(n_18474), .b(n_17900), .o(n_18761) );
in01f80 g551466 ( .a(n_18472), .o(n_18473) );
na02f80 g551467 ( .a(n_18245), .b(n_17691), .o(n_18472) );
in01f80 g551468 ( .a(n_17977), .o(n_17978) );
no02f80 g551469 ( .a(n_17750), .b(x_in_56_4), .o(n_17977) );
na02f80 g551470 ( .a(n_17750), .b(x_in_56_4), .o(n_18570) );
in01f80 g551471 ( .a(n_17748), .o(n_17749) );
no02f80 g551472 ( .a(n_17460), .b(x_in_10_4), .o(n_17748) );
na02f80 g551473 ( .a(n_17460), .b(x_in_10_4), .o(n_18303) );
na02f80 g551474 ( .a(n_18225), .b(x_in_22_4), .o(n_18566) );
no02f80 g551475 ( .a(n_18243), .b(n_18242), .o(n_18244) );
na02f80 g551476 ( .a(n_18471), .b(x_in_12_3), .o(n_19419) );
na02f80 g551477 ( .a(n_18299), .b(n_17975), .o(n_17976) );
na02f80 g551478 ( .a(n_18708), .b(x_in_20_3), .o(n_18836) );
in01f80 g551479 ( .a(n_18240), .o(n_18241) );
no02f80 g551480 ( .a(n_18708), .b(x_in_20_3), .o(n_18240) );
na02f80 g551481 ( .a(n_17459), .b(x_in_42_4), .o(n_18302) );
in01f80 g551482 ( .a(n_17746), .o(n_17747) );
no02f80 g551483 ( .a(n_17459), .b(x_in_42_4), .o(n_17746) );
no02f80 g551484 ( .a(n_18297), .b(n_17973), .o(n_17974) );
na02f80 g551485 ( .a(n_18760), .b(x_in_36_2), .o(n_19740) );
in01f80 g551486 ( .a(n_19081), .o(n_19082) );
no02f80 g551487 ( .a(n_18760), .b(x_in_36_2), .o(n_19081) );
no02f80 g551488 ( .a(n_18238), .b(n_18237), .o(n_18239) );
in01f80 g551489 ( .a(n_17971), .o(n_17972) );
na02f80 g551490 ( .a(n_17745), .b(n_17113), .o(n_17971) );
no02f80 g551491 ( .a(n_17743), .b(n_17742), .o(n_17744) );
na02f80 g551492 ( .a(n_17480), .b(n_17142), .o(n_17143) );
na02f80 g551493 ( .a(n_17458), .b(n_17742), .o(n_18623) );
in01f80 g551494 ( .a(n_18469), .o(n_18470) );
na02f80 g551495 ( .a(n_18236), .b(n_17686), .o(n_18469) );
na02f80 g551496 ( .a(n_17457), .b(n_17739), .o(n_18620) );
in01f80 g551497 ( .a(n_19398), .o(n_19399) );
no02f80 g551498 ( .a(n_19080), .b(x_in_20_2), .o(n_19398) );
no02f80 g551499 ( .a(n_17740), .b(n_17739), .o(n_17741) );
na02f80 g551500 ( .a(n_18468), .b(x_in_54_3), .o(n_19425) );
na02f80 g551501 ( .a(n_17970), .b(x_in_52_2), .o(n_18832) );
in01f80 g551502 ( .a(n_18234), .o(n_18235) );
no02f80 g551503 ( .a(n_17970), .b(x_in_52_2), .o(n_18234) );
no02f80 g551504 ( .a(n_18466), .b(n_18465), .o(n_18467) );
na02f80 g551505 ( .a(n_17738), .b(x_in_44_3), .o(n_18556) );
in01f80 g551506 ( .a(n_17968), .o(n_17969) );
no02f80 g551507 ( .a(n_17738), .b(x_in_44_3), .o(n_17968) );
na02f80 g551508 ( .a(n_18464), .b(x_in_28_5), .o(n_19434) );
in01f80 g551509 ( .a(n_18758), .o(n_18759) );
no02f80 g551510 ( .a(n_18464), .b(x_in_28_5), .o(n_18758) );
in01f80 g551511 ( .a(n_17966), .o(n_17967) );
no02f80 g551512 ( .a(n_17751), .b(x_in_26_4), .o(n_17966) );
no02f80 g551513 ( .a(n_17479), .b(n_17140), .o(n_17141) );
na02f80 g551514 ( .a(n_17456), .b(x_in_58_4), .o(n_18321) );
in01f80 g551515 ( .a(n_17736), .o(n_17737) );
no02f80 g551516 ( .a(n_17456), .b(x_in_58_4), .o(n_17736) );
na02f80 g551517 ( .a(n_18757), .b(x_in_60_2), .o(n_19745) );
in01f80 g551518 ( .a(n_19078), .o(n_19079) );
no02f80 g551519 ( .a(n_18757), .b(x_in_60_2), .o(n_19078) );
na02f80 g551520 ( .a(n_18430), .b(x_in_60_3), .o(n_18843) );
no02f80 g551521 ( .a(n_17784), .b(n_17454), .o(n_17455) );
no02f80 g551522 ( .a(n_17478), .b(n_17138), .o(n_17139) );
na02f80 g551523 ( .a(n_18027), .b(n_17734), .o(n_17735) );
na02f80 g551524 ( .a(n_17783), .b(n_17452), .o(n_17453) );
na02f80 g551525 ( .a(n_18296), .b(n_17964), .o(n_17965) );
no02f80 g551526 ( .a(n_17782), .b(n_17450), .o(n_17451) );
no02f80 g551527 ( .a(n_17477), .b(n_17136), .o(n_17137) );
na02f80 g551528 ( .a(n_18295), .b(n_17962), .o(n_17963) );
no02f80 g551529 ( .a(n_17476), .b(n_17134), .o(n_17135) );
no02f80 g551530 ( .a(n_17781), .b(n_17448), .o(n_17449) );
no02f80 g551531 ( .a(n_17159), .b(n_16880), .o(n_16881) );
na02f80 g551532 ( .a(n_18232), .b(n_18231), .o(n_18233) );
na02f80 g551533 ( .a(n_18229), .b(n_18228), .o(n_18230) );
na02f80 g551534 ( .a(n_17385), .b(n_18227), .o(n_18910) );
na02f80 g551535 ( .a(n_18225), .b(n_18227), .o(n_18226) );
na02f80 g551536 ( .a(n_18223), .b(n_18222), .o(n_18224) );
na02f80 g551537 ( .a(n_17093), .b(n_18221), .o(n_18901) );
na02f80 g551538 ( .a(n_17095), .b(n_18231), .o(n_18907) );
na02f80 g551539 ( .a(n_18219), .b(n_18218), .o(n_18220) );
na02f80 g551540 ( .a(n_18216), .b(n_18221), .o(n_18217) );
na02f80 g551541 ( .a(n_17091), .b(n_18228), .o(n_18898) );
na02f80 g551542 ( .a(n_17097), .b(n_18222), .o(n_18911) );
na02f80 g551543 ( .a(n_17087), .b(n_17733), .o(n_18895) );
na02f80 g551544 ( .a(n_17731), .b(n_17733), .o(n_17732) );
na02f80 g551545 ( .a(n_17094), .b(n_18218), .o(n_18904) );
na02f80 g551546 ( .a(n_17388), .b(n_18215), .o(n_18894) );
na02f80 g551547 ( .a(n_18213), .b(n_18215), .o(n_18214) );
no02f80 g551548 ( .a(n_17475), .b(n_17132), .o(n_17133) );
no02f80 g551549 ( .a(n_17474), .b(n_17130), .o(n_17131) );
no02f80 g551550 ( .a(n_18462), .b(n_18461), .o(n_18463) );
na02f80 g551551 ( .a(n_18212), .b(n_18461), .o(n_19475) );
na02f80 g551552 ( .a(n_17780), .b(n_17446), .o(n_17447) );
no02f80 g551553 ( .a(n_18210), .b(n_18209), .o(n_18211) );
no02f80 g551554 ( .a(n_18207), .b(n_18206), .o(n_18208) );
no02f80 g551555 ( .a(n_18204), .b(n_18203), .o(n_18205) );
no02f80 g551556 ( .a(n_18459), .b(n_18458), .o(n_18460) );
no02f80 g551557 ( .a(n_17473), .b(n_17128), .o(n_17129) );
no02f80 g551558 ( .a(n_17472), .b(n_17126), .o(n_17127) );
no02f80 g551559 ( .a(n_17471), .b(n_17124), .o(n_17125) );
na02f80 g551560 ( .a(n_17961), .b(n_17960), .o(n_18890) );
no02f80 g551561 ( .a(n_17958), .b(n_17960), .o(n_17959) );
no02f80 g551562 ( .a(n_17470), .b(n_17122), .o(n_17123) );
no02f80 g551563 ( .a(n_17777), .b(n_17444), .o(n_17445) );
no02f80 g551564 ( .a(n_16848), .b(n_17444), .o(n_18345) );
in01f80 g551565 ( .a(n_16879), .o(n_17799) );
na02f80 g551566 ( .a(n_16638), .b(n_16637), .o(n_16879) );
na02f80 g551567 ( .a(n_17469), .b(n_17120), .o(n_17121) );
no02f80 g551568 ( .a(n_19076), .b(n_19075), .o(n_19077) );
no02f80 g551569 ( .a(n_18755), .b(n_18754), .o(n_18756) );
no02f80 g551570 ( .a(n_18752), .b(n_18751), .o(n_18753) );
no02f80 g551571 ( .a(n_19073), .b(n_19072), .o(n_19074) );
no02f80 g551572 ( .a(n_19070), .b(n_19069), .o(n_19071) );
no02f80 g551573 ( .a(n_18749), .b(n_18748), .o(n_18750) );
no02f80 g551574 ( .a(n_18746), .b(n_18745), .o(n_18747) );
no02f80 g551575 ( .a(n_18743), .b(n_18742), .o(n_18744) );
no02f80 g551576 ( .a(n_18201), .b(n_18200), .o(n_18202) );
no02f80 g551577 ( .a(n_18456), .b(n_18455), .o(n_18457) );
no02f80 g551578 ( .a(n_18453), .b(n_18452), .o(n_18454) );
no02f80 g551579 ( .a(n_18740), .b(n_18739), .o(n_18741) );
no02f80 g551580 ( .a(n_18737), .b(n_18736), .o(n_18738) );
no02f80 g551581 ( .a(n_18734), .b(n_18733), .o(n_18735) );
no02f80 g551582 ( .a(n_18198), .b(n_18197), .o(n_18199) );
no02f80 g551583 ( .a(n_18731), .b(n_18730), .o(n_18732) );
no02f80 g551584 ( .a(n_18728), .b(n_18727), .o(n_18729) );
no02f80 g551585 ( .a(n_18725), .b(n_18724), .o(n_18726) );
no02f80 g551586 ( .a(n_18722), .b(n_18721), .o(n_18723) );
no02f80 g551587 ( .a(n_18195), .b(n_18194), .o(n_18196) );
no02f80 g551588 ( .a(n_18450), .b(n_18449), .o(n_18451) );
no02f80 g551589 ( .a(n_18192), .b(n_18191), .o(n_18193) );
no02f80 g551590 ( .a(n_18719), .b(n_18718), .o(n_18720) );
no02f80 g551591 ( .a(n_18447), .b(n_18446), .o(n_18448) );
in01f80 g551592 ( .a(n_19480), .o(n_18717) );
oa12f80 g551593 ( .a(n_17910), .b(n_17514), .c(n_17360), .o(n_19480) );
no02f80 g551594 ( .a(n_18189), .b(n_18188), .o(n_18190) );
na02f80 g551595 ( .a(n_17456), .b(n_17722), .o(n_17443) );
in01f80 g551596 ( .a(n_18187), .o(n_18884) );
no02f80 g551597 ( .a(n_17770), .b(n_17957), .o(n_18187) );
in01f80 g551598 ( .a(n_19823), .o(n_18716) );
oa12f80 g551599 ( .a(n_18134), .b(n_17598), .c(n_17513), .o(n_19823) );
na02f80 g551600 ( .a(n_18490), .b(n_18710), .o(n_18445) );
in01f80 g551601 ( .a(n_18186), .o(n_18881) );
no02f80 g551602 ( .a(n_17995), .b(n_17956), .o(n_18186) );
in01f80 g551603 ( .a(n_19820), .o(n_18715) );
oa12f80 g551604 ( .a(n_18142), .b(n_17596), .c(n_17512), .o(n_19820) );
na02f80 g551605 ( .a(n_17092), .b(n_17730), .o(n_18596) );
na02f80 g551606 ( .a(n_17728), .b(n_17730), .o(n_17729) );
in01f80 g551607 ( .a(n_20172), .o(n_18714) );
oa12f80 g551608 ( .a(n_18398), .b(n_17840), .c(n_17212), .o(n_20172) );
na02f80 g551609 ( .a(n_17088), .b(n_17727), .o(n_18611) );
na02f80 g551610 ( .a(n_17725), .b(n_17727), .o(n_17726) );
in01f80 g551611 ( .a(n_20169), .o(n_18713) );
oa12f80 g551612 ( .a(n_18407), .b(n_17838), .c(n_17211), .o(n_20169) );
in01f80 g551613 ( .a(n_19229), .o(n_18712) );
oa12f80 g551614 ( .a(n_17699), .b(n_17511), .c(n_17068), .o(n_19229) );
no02f80 g551615 ( .a(n_18189), .b(n_17532), .o(n_18887) );
in01f80 g551616 ( .a(n_19817), .o(n_18444) );
oa12f80 g551617 ( .a(n_18141), .b(n_17592), .c(n_16965), .o(n_19817) );
in01f80 g551618 ( .a(n_18337), .o(n_17955) );
na02f80 g551619 ( .a(n_17084), .b(n_17724), .o(n_18337) );
na02f80 g551620 ( .a(n_17459), .b(n_17724), .o(n_17442) );
in01f80 g551621 ( .a(n_19787), .o(n_18443) );
oa12f80 g551622 ( .a(n_18138), .b(n_17590), .c(n_16964), .o(n_19787) );
in01f80 g551623 ( .a(n_18185), .o(n_18876) );
no02f80 g551624 ( .a(n_17751), .b(n_17954), .o(n_18185) );
in01f80 g551625 ( .a(n_19814), .o(n_18442) );
oa12f80 g551626 ( .a(n_17895), .b(n_17354), .c(n_17208), .o(n_19814) );
in01f80 g551627 ( .a(n_18339), .o(n_17953) );
na02f80 g551628 ( .a(n_17086), .b(n_17723), .o(n_18339) );
in01f80 g551629 ( .a(n_20156), .o(n_18441) );
oa12f80 g551630 ( .a(n_18130), .b(n_17553), .c(n_16959), .o(n_20156) );
na02f80 g551631 ( .a(n_17083), .b(n_17722), .o(n_18605) );
na02f80 g551632 ( .a(n_17951), .b(n_17956), .o(n_17952) );
in01f80 g551633 ( .a(n_19780), .o(n_18440) );
oa12f80 g551634 ( .a(n_18137), .b(n_17572), .c(n_16962), .o(n_19780) );
no02f80 g551635 ( .a(n_18179), .b(n_17517), .o(n_18862) );
in01f80 g551636 ( .a(n_20153), .o(n_18439) );
oa12f80 g551637 ( .a(n_18122), .b(n_17583), .c(n_16961), .o(n_20153) );
in01f80 g551638 ( .a(n_20162), .o(n_18438) );
oa12f80 g551639 ( .a(n_18123), .b(n_17581), .c(n_16960), .o(n_20162) );
in01f80 g551640 ( .a(n_19260), .o(n_18711) );
oa12f80 g551641 ( .a(n_17693), .b(n_17047), .c(n_17507), .o(n_19260) );
in01f80 g551642 ( .a(n_19496), .o(n_18437) );
oa12f80 g551643 ( .a(n_17697), .b(n_17064), .c(n_17202), .o(n_19496) );
in01f80 g551644 ( .a(n_20150), .o(n_18436) );
oa12f80 g551645 ( .a(n_18132), .b(n_17578), .c(n_16952), .o(n_20150) );
in01f80 g551646 ( .a(n_17950), .o(n_18606) );
na02f80 g551647 ( .a(n_18011), .b(n_17000), .o(n_17950) );
in01f80 g551648 ( .a(n_20159), .o(n_18435) );
oa12f80 g551649 ( .a(n_18133), .b(n_17576), .c(n_16958), .o(n_20159) );
ao12f80 g551650 ( .a(n_11573), .b(n_17441), .c(n_12510), .o(n_18326) );
in01f80 g551651 ( .a(n_20137), .o(n_18434) );
oa12f80 g551652 ( .a(n_18119), .b(n_17574), .c(n_16957), .o(n_20137) );
no02f80 g551653 ( .a(n_18011), .b(n_17720), .o(n_17721) );
in01f80 g551654 ( .a(n_20166), .o(n_19068) );
oa12f80 g551655 ( .a(n_18143), .b(n_17814), .c(n_17570), .o(n_20166) );
na02f80 g551656 ( .a(n_17948), .b(n_17954), .o(n_17949) );
oa12f80 g551657 ( .a(n_10783), .b(n_17440), .c(n_12046), .o(n_18334) );
na02f80 g551658 ( .a(n_17853), .b(n_18433), .o(n_19188) );
na02f80 g551659 ( .a(n_18246), .b(n_18433), .o(n_18184) );
no02f80 g551660 ( .a(FE_OFN722_n_17438), .b(n_17437), .o(n_17439) );
no02f80 g551661 ( .a(FE_OFN722_n_17438), .b(n_16791), .o(n_18331) );
na02f80 g551662 ( .a(n_18183), .b(n_17529), .o(n_18875) );
na02f80 g551663 ( .a(n_18183), .b(n_17946), .o(n_17947) );
in01f80 g551664 ( .a(n_19790), .o(n_18182) );
oa12f80 g551665 ( .a(n_17901), .b(n_17332), .c(n_16956), .o(n_19790) );
in01f80 g551666 ( .a(n_19194), .o(n_18181) );
oa12f80 g551667 ( .a(n_17912), .b(n_17320), .c(n_16949), .o(n_19194) );
no02f80 g551668 ( .a(n_17718), .b(n_17717), .o(n_17719) );
in01f80 g551669 ( .a(n_17945), .o(n_18602) );
na02f80 g551670 ( .a(n_17716), .b(n_17717), .o(n_17945) );
ao12f80 g551671 ( .a(n_8314), .b(n_17715), .c(n_9528), .o(n_18584) );
na02f80 g551672 ( .a(n_18179), .b(n_18178), .o(n_18180) );
na02f80 g551673 ( .a(n_17386), .b(n_17944), .o(n_18867) );
na02f80 g551674 ( .a(n_17769), .b(n_17944), .o(n_17714) );
in01f80 g551675 ( .a(n_19784), .o(n_18432) );
oa12f80 g551676 ( .a(n_17689), .b(n_17207), .c(n_17052), .o(n_19784) );
in01f80 g551677 ( .a(FE_OFN672_n_17494), .o(n_16878) );
ao22s80 g551678 ( .a(n_16636), .b(n_11126), .c(n_11128), .d(n_11687), .o(n_17494) );
na02f80 g551679 ( .a(n_18430), .b(n_18429), .o(n_18431) );
in01f80 g551680 ( .a(n_17943), .o(n_18593) );
no02f80 g551681 ( .a(n_17752), .b(n_17713), .o(n_17943) );
na02f80 g551682 ( .a(n_17435), .b(n_17713), .o(n_17436) );
no02f80 g551683 ( .a(FE_OFN1017_n_17433), .b(n_17432), .o(n_17434) );
no02f80 g551684 ( .a(FE_OFN1017_n_17433), .b(n_16781), .o(n_18590) );
in01f80 g551685 ( .a(n_19493), .o(n_19067) );
oa12f80 g551686 ( .a(n_18408), .b(n_17813), .c(n_17820), .o(n_19493) );
na02f80 g551687 ( .a(n_17460), .b(n_17723), .o(n_17431) );
in01f80 g551688 ( .a(n_19460), .o(n_19066) );
na02f80 g551689 ( .a(n_18102), .b(n_18710), .o(n_19460) );
na02f80 g551690 ( .a(n_18708), .b(n_18707), .o(n_18709) );
na02f80 g551691 ( .a(n_17614), .b(n_18177), .o(n_18865) );
na02f80 g551692 ( .a(n_18003), .b(n_18177), .o(n_17942) );
no02f80 g551693 ( .a(n_18015), .b(n_17711), .o(n_17712) );
na02f80 g551694 ( .a(n_17940), .b(n_17957), .o(n_17941) );
no02f80 g551695 ( .a(n_17096), .b(n_17711), .o(n_18585) );
in01f80 g551696 ( .a(n_20140), .o(n_18428) );
oa12f80 g551697 ( .a(n_18131), .b(n_17551), .c(n_16953), .o(n_20140) );
no02f80 g551698 ( .a(n_18708), .b(n_18100), .o(n_19458) );
no02f80 g551699 ( .a(n_18430), .b(n_17815), .o(n_19189) );
in01f80 g551700 ( .a(n_19215), .o(n_18706) );
oa12f80 g551701 ( .a(n_18405), .b(n_17836), .c(n_16988), .o(n_19215) );
in01f80 g551702 ( .a(n_18427), .o(n_19448) );
oa12f80 g551703 ( .a(n_16920), .b(n_18164), .c(n_16406), .o(n_18427) );
ao12f80 g551704 ( .a(n_12451), .b(n_17119), .c(n_13640), .o(n_18046) );
in01f80 g551705 ( .a(n_18176), .o(n_19176) );
oa12f80 g551706 ( .a(n_17897), .b(n_17350), .c(n_15353), .o(n_18176) );
in01f80 g551707 ( .a(n_19200), .o(n_18705) );
oa12f80 g551708 ( .a(n_17896), .b(n_17345), .c(n_17531), .o(n_19200) );
in01f80 g551709 ( .a(n_19257), .o(n_18704) );
oa12f80 g551710 ( .a(n_18406), .b(n_17834), .c(n_16990), .o(n_19257) );
in01f80 g551711 ( .a(n_18175), .o(n_19170) );
oa12f80 g551712 ( .a(n_16592), .b(n_17931), .c(n_15975), .o(n_18175) );
in01f80 g551713 ( .a(n_17710), .o(n_18580) );
oa12f80 g551714 ( .a(n_3272), .b(n_17426), .c(n_2190), .o(n_17710) );
in01f80 g551715 ( .a(n_19254), .o(n_18703) );
oa12f80 g551716 ( .a(n_18404), .b(n_17832), .c(n_16986), .o(n_19254) );
in01f80 g551717 ( .a(n_19795), .o(n_19397) );
oa12f80 g551718 ( .a(n_17907), .b(n_17337), .c(n_18101), .o(n_19795) );
in01f80 g551719 ( .a(n_19249), .o(n_18702) );
oa12f80 g551720 ( .a(n_18403), .b(n_17830), .c(n_16985), .o(n_19249) );
in01f80 g551721 ( .a(n_19246), .o(n_18426) );
oa12f80 g551722 ( .a(n_17906), .b(n_17335), .c(n_17256), .o(n_19246) );
in01f80 g551723 ( .a(n_19243), .o(n_18701) );
oa12f80 g551724 ( .a(n_18402), .b(n_17828), .c(n_17253), .o(n_19243) );
in01f80 g551725 ( .a(n_18944), .o(n_18425) );
oa12f80 g551726 ( .a(n_17694), .b(n_17057), .c(n_17252), .o(n_18944) );
in01f80 g551727 ( .a(n_19232), .o(n_18700) );
oa12f80 g551728 ( .a(n_18400), .b(n_17824), .c(n_16982), .o(n_19232) );
in01f80 g551729 ( .a(n_19238), .o(n_18699) );
oa12f80 g551730 ( .a(n_18401), .b(n_17826), .c(n_16983), .o(n_19238) );
in01f80 g551731 ( .a(n_17939), .o(n_18856) );
oa12f80 g551732 ( .a(n_14837), .b(n_17706), .c(n_13744), .o(n_17939) );
in01f80 g551733 ( .a(n_17709), .o(n_18578) );
oa12f80 g551734 ( .a(n_3258), .b(n_17424), .c(n_2183), .o(n_17709) );
in01f80 g551735 ( .a(n_19222), .o(n_18698) );
oa12f80 g551736 ( .a(n_17417), .b(n_16834), .c(n_17528), .o(n_19222) );
in01f80 g551737 ( .a(n_19197), .o(n_18697) );
oa12f80 g551738 ( .a(n_17894), .b(n_17520), .c(n_17339), .o(n_19197) );
in01f80 g551739 ( .a(n_18424), .o(n_19454) );
oa12f80 g551740 ( .a(n_17413), .b(n_17241), .c(n_16832), .o(n_18424) );
in01f80 g551741 ( .a(n_18174), .o(n_19165) );
oa12f80 g551742 ( .a(n_16910), .b(n_17938), .c(n_16412), .o(n_18174) );
in01f80 g551743 ( .a(n_17708), .o(n_18583) );
oa12f80 g551744 ( .a(n_17331), .b(n_17430), .c(n_16744), .o(n_17708) );
ao12f80 g551745 ( .a(n_13625), .b(n_17429), .c(n_14650), .o(n_18327) );
in01f80 g551746 ( .a(n_19210), .o(n_18696) );
oa12f80 g551747 ( .a(n_17684), .b(n_17524), .c(n_17049), .o(n_19210) );
in01f80 g551748 ( .a(n_17937), .o(n_18854) );
oa12f80 g551749 ( .a(n_14499), .b(n_17703), .c(n_13299), .o(n_17937) );
in01f80 g551750 ( .a(n_19206), .o(n_18695) );
oa12f80 g551751 ( .a(n_17683), .b(n_17530), .c(n_17045), .o(n_19206) );
in01f80 g551752 ( .a(n_18173), .o(n_19173) );
oa12f80 g551753 ( .a(n_17892), .b(n_17317), .c(n_14210), .o(n_18173) );
in01f80 g551754 ( .a(n_18979), .o(n_18423) );
oa12f80 g551755 ( .a(n_17700), .b(n_17231), .c(n_17040), .o(n_18979) );
oa12f80 g551756 ( .a(n_17843), .b(n_17395), .c(n_16800), .o(n_18422) );
oa12f80 g551757 ( .a(n_17363), .b(n_17621), .c(n_16043), .o(n_17936) );
oa12f80 g551758 ( .a(n_17362), .b(n_17397), .c(n_16038), .o(n_17935) );
ao12f80 g551759 ( .a(n_12366), .b(n_15993), .c(n_4929), .o(n_16886) );
oa12f80 g551760 ( .a(n_11825), .b(n_16636), .c(n_10697), .o(n_17165) );
ao12f80 g551761 ( .a(n_11506), .b(n_16877), .c(n_12490), .o(n_17800) );
ao12f80 g551762 ( .a(n_11810), .b(n_17118), .c(n_13111), .o(n_18044) );
in01f80 g551763 ( .a(n_20132), .o(n_18172) );
oa12f80 g551764 ( .a(n_17210), .b(n_17934), .c(n_17209), .o(n_20132) );
in01f80 g551765 ( .a(n_20481), .o(n_19065) );
oa12f80 g551766 ( .a(n_17510), .b(n_18694), .c(n_17509), .o(n_20481) );
in01f80 g551767 ( .a(n_20879), .o(n_18693) );
oa12f80 g551768 ( .a(n_17505), .b(n_18421), .c(n_17504), .o(n_20879) );
in01f80 g551769 ( .a(n_20484), .o(n_18420) );
oa12f80 g551770 ( .a(n_17216), .b(n_18171), .c(n_17215), .o(n_20484) );
ao22s80 g551771 ( .a(n_18171), .b(n_17191), .c(n_17501), .d(x_in_60_1), .o(n_19130) );
ao12f80 g551772 ( .a(n_18118), .b(n_18117), .c(n_18116), .o(n_18692) );
ao12f80 g551773 ( .a(n_17679), .b(n_17681), .c(n_17678), .o(n_18170) );
in01f80 g551774 ( .a(n_17789), .o(n_18029) );
ao12f80 g551775 ( .a(n_16633), .b(n_16877), .c(n_16632), .o(n_17789) );
ao12f80 g551776 ( .a(n_18115), .b(n_18114), .c(n_18113), .o(n_18691) );
in01f80 g551777 ( .a(n_18829), .o(n_18419) );
oa12f80 g551778 ( .a(n_17677), .b(n_17889), .c(n_17692), .o(n_18829) );
ao12f80 g551779 ( .a(n_17884), .b(n_17883), .c(n_17882), .o(n_18418) );
ao12f80 g551780 ( .a(n_17876), .b(n_17875), .c(n_17874), .o(n_18417) );
ao12f80 g551781 ( .a(n_17676), .b(n_17675), .c(n_17674), .o(n_18169) );
ao12f80 g551782 ( .a(n_17881), .b(n_17880), .c(n_19129), .o(n_18416) );
in01f80 g551783 ( .a(n_17933), .o(n_18851) );
oa12f80 g551784 ( .a(n_17105), .b(n_17441), .c(n_17104), .o(n_17933) );
ao12f80 g551785 ( .a(n_17673), .b(n_17672), .c(n_17671), .o(n_18168) );
ao12f80 g551786 ( .a(n_17670), .b(n_17669), .c(n_18822), .o(n_18167) );
ao12f80 g551787 ( .a(n_17879), .b(n_17878), .c(n_17877), .o(n_18415) );
ao12f80 g551788 ( .a(n_17668), .b(n_17667), .c(n_17666), .o(n_18166) );
ao12f80 g551789 ( .a(n_16861), .b(n_16862), .c(n_16860), .o(n_17428) );
in01f80 g551790 ( .a(n_18545), .o(n_18319) );
ao12f80 g551791 ( .a(n_16872), .b(n_17119), .c(n_16871), .o(n_18545) );
ao22s80 g551792 ( .a(n_17934), .b(n_16928), .c(n_17197), .d(x_in_6_1), .o(n_18823) );
oa12f80 g551793 ( .a(n_17869), .b(n_17870), .c(n_17868), .o(n_19143) );
ao22s80 g551794 ( .a(n_18164), .b(n_17180), .c(n_17230), .d(n_17179), .o(n_18165) );
ao12f80 g551795 ( .a(n_17665), .b(n_17664), .c(n_17663), .o(n_18163) );
ao12f80 g551796 ( .a(n_17659), .b(n_17658), .c(n_17657), .o(n_18162) );
ao12f80 g551797 ( .a(n_17656), .b(n_17655), .c(n_17654), .o(n_18161) );
ao12f80 g551798 ( .a(n_17653), .b(n_17652), .c(n_17651), .o(n_18160) );
ao12f80 g551799 ( .a(n_17650), .b(n_17649), .c(n_17648), .o(n_18159) );
ao22s80 g551800 ( .a(n_16827), .b(n_17931), .c(n_16826), .d(n_17002), .o(n_17932) );
ao22s80 g551801 ( .a(n_17426), .b(n_3705), .c(n_16568), .d(n_3704), .o(n_17427) );
ao12f80 g551802 ( .a(n_18112), .b(n_18111), .c(n_19737), .o(n_18690) );
in01f80 g551803 ( .a(n_18575), .o(n_18834) );
ao12f80 g551804 ( .a(n_17111), .b(n_17440), .c(n_17110), .o(n_18575) );
ao12f80 g551805 ( .a(n_17408), .b(n_17407), .c(n_26552), .o(n_26838) );
ao22s80 g551806 ( .a(n_17706), .b(n_15038), .c(n_16776), .d(n_15037), .o(n_17707) );
ao12f80 g551807 ( .a(n_17647), .b(n_17646), .c(n_17645), .o(n_18158) );
ao12f80 g551808 ( .a(n_18129), .b(n_18128), .c(n_18127), .o(n_18689) );
in01f80 g551809 ( .a(n_16635), .o(n_17492) );
oa12f80 g551810 ( .a(n_15652), .b(n_15993), .c(n_15651), .o(n_16635) );
in01f80 g551811 ( .a(n_18301), .o(n_18304) );
ao12f80 g551812 ( .a(n_16870), .b(n_16869), .c(n_16868), .o(n_18301) );
oa12f80 g551813 ( .a(n_17103), .b(n_17109), .c(n_17401), .o(n_18313) );
ao12f80 g551814 ( .a(n_17662), .b(n_17661), .c(n_17660), .o(n_18157) );
no03m80 g551815 ( .a(n_7567), .b(n_17405), .c(n_8891), .o(n_18156) );
ao22s80 g551816 ( .a(n_16567), .b(n_3700), .c(n_17424), .d(n_3701), .o(n_17425) );
ao12f80 g551817 ( .a(n_17891), .b(n_17890), .c(n_18151), .o(n_18414) );
in01f80 g551818 ( .a(n_18554), .o(n_18827) );
ao12f80 g551819 ( .a(n_17410), .b(n_17715), .c(n_17409), .o(n_18554) );
ao12f80 g551820 ( .a(n_18126), .b(n_18125), .c(n_18124), .o(n_18688) );
in01f80 g551821 ( .a(n_18846), .o(n_18831) );
ao12f80 g551822 ( .a(n_17403), .b(n_17404), .c(n_17402), .o(n_18846) );
ao12f80 g551823 ( .a(n_16631), .b(n_16630), .c(n_16629), .o(n_17117) );
in01f80 g551824 ( .a(n_17491), .o(n_17116) );
oa12f80 g551825 ( .a(n_16345), .b(n_16636), .c(n_16344), .o(n_17491) );
oa12f80 g551826 ( .a(n_16867), .b(n_16866), .c(n_16865), .o(n_18036) );
in01f80 g551827 ( .a(n_17930), .o(n_18849) );
oa12f80 g551828 ( .a(n_17108), .b(n_17429), .c(n_17107), .o(n_17930) );
ao22s80 g551829 ( .a(n_17557), .b(n_17430), .c(n_17556), .d(n_16574), .o(n_18413) );
ao12f80 g551830 ( .a(n_17867), .b(n_17866), .c(n_17865), .o(n_18412) );
in01f80 g551831 ( .a(n_18549), .o(n_17705) );
oa12f80 g551832 ( .a(n_16864), .b(n_17118), .c(n_16863), .o(n_18549) );
ao22s80 g551833 ( .a(n_16774), .b(n_14833), .c(n_17703), .d(n_14834), .o(n_17704) );
ao22s80 g551834 ( .a(n_18694), .b(n_17497), .c(n_18099), .d(x_in_36_1), .o(n_19738) );
ao22s80 g551835 ( .a(n_17938), .b(n_17176), .c(n_16970), .d(n_17175), .o(n_18155) );
ao22s80 g551836 ( .a(n_18421), .b(n_17498), .c(n_17811), .d(x_in_20_1), .o(n_19415) );
ao12f80 g551837 ( .a(n_17644), .b(n_17643), .c(n_17642), .o(n_18154) );
ao12f80 g551838 ( .a(n_16348), .b(n_16347), .c(n_16346), .o(n_16876) );
ao12f80 g551839 ( .a(n_17641), .b(n_17640), .c(n_17639), .o(n_18153) );
ao12f80 g551840 ( .a(n_18110), .b(n_18109), .c(n_19414), .o(n_18687) );
oa12f80 g551841 ( .a(n_17872), .b(n_17873), .c(n_17871), .o(n_19132) );
oa22f80 g551842 ( .a(n_16948), .b(FE_OFN248_n_4162), .c(n_330), .d(FE_OFN60_n_27012), .o(n_17929) );
oa22f80 g551843 ( .a(n_16561), .b(n_29046), .c(n_1577), .d(FE_OFN60_n_27012), .o(n_17423) );
oa22f80 g551844 ( .a(n_16947), .b(FE_OFN235_n_4162), .c(n_883), .d(FE_OFN364_n_4860), .o(n_17928) );
oa22f80 g551845 ( .a(n_18151), .b(FE_OFN260_n_4280), .c(n_1751), .d(FE_OFN1112_rst), .o(n_18152) );
oa22f80 g551846 ( .a(n_17812), .b(FE_OFN406_n_28303), .c(n_122), .d(FE_OFN360_n_4860), .o(n_18686) );
oa22f80 g551847 ( .a(n_16564), .b(FE_OFN219_n_23315), .c(n_1398), .d(FE_OFN113_n_27449), .o(n_17422) );
oa22f80 g551848 ( .a(n_16343), .b(FE_OFN148_n_25677), .c(n_991), .d(FE_OFN1111_rst), .o(n_16634) );
oa22f80 g551849 ( .a(n_17201), .b(FE_OFN162_n_26454), .c(n_99), .d(FE_OFN1146_n_4860), .o(n_18150) );
oa22f80 g551850 ( .a(FE_OFN450_n_17680), .b(n_29046), .c(n_890), .d(n_27449), .o(n_17702) );
oa22f80 g551851 ( .a(n_16945), .b(n_28303), .c(n_1349), .d(FE_OFN95_n_27449), .o(n_17927) );
oa22f80 g551852 ( .a(n_17503), .b(FE_OFN314_n_3069), .c(n_840), .d(FE_OFN72_n_27012), .o(n_18411) );
oa22f80 g551853 ( .a(FE_OFN1001_n_17200), .b(n_29691), .c(n_1301), .d(FE_OFN122_n_27449), .o(n_18149) );
oa22f80 g551854 ( .a(n_16300), .b(FE_OFN266_n_4280), .c(n_1471), .d(FE_OFN347_n_4860), .o(n_17115) );
oa22f80 g551855 ( .a(n_16944), .b(FE_OFN406_n_28303), .c(n_1634), .d(FE_OFN355_n_4860), .o(n_17926) );
oa22f80 g551856 ( .a(n_16943), .b(n_26454), .c(n_1926), .d(FE_OFN94_n_27449), .o(n_17925) );
oa22f80 g551857 ( .a(n_17199), .b(FE_OFN417_n_28303), .c(n_1880), .d(FE_OFN139_n_27449), .o(n_18148) );
oa22f80 g551858 ( .a(n_16757), .b(FE_OFN175_n_26184), .c(n_919), .d(FE_OFN350_n_4860), .o(n_17701) );
oa22f80 g551859 ( .a(n_18127), .b(FE_OFN240_n_4162), .c(n_6), .d(FE_OFN141_n_27449), .o(n_17924) );
oa22f80 g551860 ( .a(n_16941), .b(FE_OFN265_n_4280), .c(n_517), .d(FE_OFN129_n_27449), .o(n_17923) );
oa22f80 g551861 ( .a(n_16940), .b(FE_OFN249_n_4162), .c(n_68), .d(FE_OFN324_n_4860), .o(n_17922) );
oa22f80 g551862 ( .a(n_17198), .b(FE_OFN254_n_4280), .c(n_583), .d(FE_OFN361_n_4860), .o(n_18147) );
oa22f80 g551863 ( .a(n_16560), .b(FE_OFN295_n_3069), .c(n_95), .d(FE_OFN360_n_4860), .o(n_17421) );
oa22f80 g551864 ( .a(FE_OFN530_n_16938), .b(n_23291), .c(n_1811), .d(FE_OFN336_n_4860), .o(n_17921) );
oa22f80 g551865 ( .a(n_17502), .b(FE_OFN413_n_28303), .c(n_1740), .d(FE_OFN141_n_27449), .o(n_18410) );
oa22f80 g551866 ( .a(n_15991), .b(n_4162), .c(n_30), .d(FE_OFN129_n_27449), .o(n_16350) );
oa22f80 g551867 ( .a(n_16937), .b(FE_OFN158_n_28014), .c(n_1251), .d(FE_OFN104_n_27449), .o(n_17920) );
oa22f80 g551868 ( .a(n_17195), .b(FE_OFN269_n_4280), .c(n_1206), .d(FE_OFN335_n_4860), .o(n_18146) );
oa22f80 g551869 ( .a(FE_OFN424_n_16296), .b(FE_OFN234_n_4162), .c(n_1147), .d(n_28607), .o(n_17114) );
oa22f80 g551870 ( .a(n_16936), .b(FE_OFN260_n_4280), .c(n_160), .d(FE_OFN127_n_27449), .o(n_17919) );
oa22f80 g551871 ( .a(FE_OFN486_n_17500), .b(n_23813), .c(n_848), .d(FE_OFN357_n_4860), .o(n_18409) );
oa22f80 g551872 ( .a(FE_OFN813_n_15982), .b(FE_OFN400_n_28303), .c(n_832), .d(n_27709), .o(n_16875) );
oa22f80 g551873 ( .a(n_16935), .b(FE_OFN412_n_28303), .c(n_879), .d(FE_OFN65_n_27012), .o(n_17918) );
oa22f80 g551874 ( .a(n_17888), .b(n_21988), .c(n_1032), .d(n_27449), .o(n_18145) );
oa22f80 g551875 ( .a(FE_OFN993_n_16934), .b(n_21988), .c(n_1568), .d(n_29261), .o(n_17917) );
oa22f80 g551876 ( .a(n_16933), .b(FE_OFN239_n_4162), .c(n_688), .d(FE_OFN136_n_27449), .o(n_17916) );
oa22f80 g551877 ( .a(n_16563), .b(FE_OFN300_n_3069), .c(n_1544), .d(FE_OFN56_n_27012), .o(n_17420) );
oa22f80 g551878 ( .a(n_16946), .b(FE_OFN239_n_4162), .c(n_1461), .d(FE_OFN350_n_4860), .o(n_17915) );
oa22f80 g551879 ( .a(n_16931), .b(FE_OFN236_n_4162), .c(n_1917), .d(FE_OFN105_n_27449), .o(n_17914) );
oa22f80 g551880 ( .a(n_15981), .b(FE_OFN265_n_4280), .c(n_1038), .d(FE_OFN1113_rst), .o(n_16874) );
oa22f80 g551881 ( .a(n_17193), .b(FE_OFN402_n_28303), .c(n_1395), .d(FE_OFN1108_rst), .o(n_18144) );
oa22f80 g551882 ( .a(n_16932), .b(n_29683), .c(n_524), .d(FE_OFN89_n_27449), .o(n_17913) );
na02f80 g551959 ( .a(n_18408), .b(n_17821), .o(n_19076) );
na02f80 g551960 ( .a(n_18143), .b(n_17571), .o(n_18722) );
na02f80 g551961 ( .a(n_17700), .b(n_17041), .o(n_18269) );
na02f80 g551962 ( .a(n_17912), .b(n_17321), .o(n_18447) );
na02f80 g551963 ( .a(n_18407), .b(n_17839), .o(n_19070) );
na02f80 g551964 ( .a(n_16873), .b(x_in_24_5), .o(n_17745) );
in01f80 g551965 ( .a(n_17112), .o(n_17113) );
no02f80 g551966 ( .a(n_16873), .b(x_in_24_5), .o(n_17112) );
na02f80 g551967 ( .a(n_18142), .b(n_17597), .o(n_18752) );
na02f80 g551968 ( .a(n_18141), .b(n_17593), .o(n_18749) );
in01f80 g551969 ( .a(n_18139), .o(n_18140) );
na02f80 g551970 ( .a(n_17911), .b(n_17330), .o(n_18139) );
na02f80 g551971 ( .a(n_18138), .b(n_17591), .o(n_18743) );
na02f80 g551972 ( .a(n_17699), .b(n_17069), .o(n_18201) );
na02f80 g551973 ( .a(n_17910), .b(n_17361), .o(n_18456) );
na02f80 g551974 ( .a(n_17868), .b(x_in_38_6), .o(n_18002) );
na02f80 g551975 ( .a(n_18137), .b(n_17573), .o(n_18746) );
in01f80 g551976 ( .a(n_18135), .o(n_18136) );
no02f80 g551977 ( .a(n_17898), .b(x_in_38_4), .o(n_18135) );
na02f80 g551978 ( .a(n_18134), .b(n_17599), .o(n_18755) );
na02f80 g551979 ( .a(n_18406), .b(n_17835), .o(n_19102) );
na02f80 g551980 ( .a(n_18133), .b(n_17577), .o(n_18728) );
na02f80 g551981 ( .a(n_18405), .b(n_17837), .o(n_19099) );
in01f80 g551982 ( .a(n_17418), .o(n_17419) );
no02f80 g551983 ( .a(n_17868), .b(x_in_38_6), .o(n_17418) );
na02f80 g551984 ( .a(n_18132), .b(n_17579), .o(n_18737) );
no02f80 g551985 ( .a(n_17119), .b(n_16871), .o(n_16872) );
in01f80 g551986 ( .a(n_17908), .o(n_17909) );
na02f80 g551987 ( .a(n_17698), .b(n_17073), .o(n_17908) );
na02f80 g551988 ( .a(n_18404), .b(n_17833), .o(n_19096) );
na02f80 g551989 ( .a(n_18403), .b(n_17831), .o(n_19093) );
na02f80 g551990 ( .a(n_17697), .b(n_17065), .o(n_18195) );
na02f80 g551991 ( .a(n_17907), .b(n_17338), .o(n_18488) );
no02f80 g551992 ( .a(n_17440), .b(n_17110), .o(n_17111) );
na02f80 g551993 ( .a(n_17906), .b(n_17336), .o(n_18485) );
na02f80 g551994 ( .a(n_18402), .b(n_17829), .o(n_19090) );
na02f80 g551995 ( .a(n_18131), .b(n_17552), .o(n_18719) );
na02f80 g551996 ( .a(n_18401), .b(n_17827), .o(n_19087) );
in01f80 g551997 ( .a(n_17904), .o(n_17905) );
na02f80 g551998 ( .a(n_17696), .b(n_17056), .o(n_17904) );
na02f80 g551999 ( .a(n_17695), .b(x_in_0_13), .o(n_18483) );
in01f80 g552000 ( .a(n_17902), .o(n_17903) );
no02f80 g552001 ( .a(n_17695), .b(x_in_0_13), .o(n_17902) );
na02f80 g552002 ( .a(n_17694), .b(n_17058), .o(n_18255) );
na02f80 g552003 ( .a(n_18130), .b(n_17554), .o(n_18731) );
na02f80 g552004 ( .a(n_17693), .b(n_17048), .o(n_18198) );
no02f80 g552005 ( .a(n_18128), .b(n_18127), .o(n_18129) );
no02f80 g552006 ( .a(n_18128), .b(n_16942), .o(n_18833) );
na02f80 g552007 ( .a(n_17901), .b(n_17333), .o(n_18450) );
no02f80 g552008 ( .a(n_16869), .b(n_16868), .o(n_16870) );
na02f80 g552009 ( .a(n_18400), .b(n_17825), .o(n_19084) );
na02f80 g552010 ( .a(n_15991), .b(n_16346), .o(n_17167) );
na02f80 g552011 ( .a(n_17417), .b(n_16835), .o(n_17984) );
no02f80 g552012 ( .a(n_18125), .b(n_18124), .o(n_18126) );
in01f80 g552013 ( .a(n_18684), .o(n_18685) );
na02f80 g552014 ( .a(n_18399), .b(n_17823), .o(n_18684) );
na02f80 g552015 ( .a(n_17692), .b(x_in_44_4), .o(n_18474) );
in01f80 g552016 ( .a(n_17899), .o(n_17900) );
no02f80 g552017 ( .a(n_17692), .b(x_in_44_4), .o(n_17899) );
in01f80 g552018 ( .a(n_17415), .o(n_17416) );
no02f80 g552019 ( .a(n_17109), .b(x_in_48_2), .o(n_17415) );
na02f80 g552020 ( .a(n_17414), .b(x_in_24_4), .o(n_18245) );
in01f80 g552021 ( .a(n_17690), .o(n_17691) );
no02f80 g552022 ( .a(n_17414), .b(x_in_24_4), .o(n_17690) );
na02f80 g552023 ( .a(n_17898), .b(x_in_38_4), .o(n_18781) );
na02f80 g552024 ( .a(n_18123), .b(n_17582), .o(n_18734) );
na02f80 g552025 ( .a(n_17429), .b(n_17107), .o(n_17108) );
na02f80 g552026 ( .a(n_18398), .b(n_17841), .o(n_19073) );
na02f80 g552027 ( .a(n_17689), .b(n_17053), .o(n_18192) );
na02f80 g552028 ( .a(n_17413), .b(n_16833), .o(n_17980) );
in01f80 g552029 ( .a(n_17687), .o(n_17688) );
na02f80 g552030 ( .a(n_17412), .b(n_16843), .o(n_17687) );
na02f80 g552031 ( .a(n_18122), .b(n_17584), .o(n_18740) );
na02f80 g552032 ( .a(n_17411), .b(x_in_28_6), .o(n_18236) );
in01f80 g552033 ( .a(n_17685), .o(n_17686) );
no02f80 g552034 ( .a(n_17411), .b(x_in_28_6), .o(n_17685) );
na02f80 g552035 ( .a(n_17109), .b(x_in_48_2), .o(n_17988) );
na02f80 g552036 ( .a(n_17684), .b(n_17050), .o(n_18243) );
na02f80 g552037 ( .a(n_17897), .b(n_17351), .o(n_18498) );
na02f80 g552038 ( .a(n_17683), .b(n_17046), .o(n_18238) );
na02f80 g552039 ( .a(n_17896), .b(n_17346), .o(n_18492) );
na02f80 g552040 ( .a(n_17895), .b(n_17355), .o(n_18453) );
na02f80 g552041 ( .a(n_17894), .b(n_17340), .o(n_18466) );
no02f80 g552042 ( .a(n_16347), .b(n_16346), .o(n_16348) );
na02f80 g552043 ( .a(n_17893), .b(x_in_28_4), .o(n_18784) );
in01f80 g552044 ( .a(n_18120), .o(n_18121) );
no02f80 g552045 ( .a(n_17893), .b(x_in_28_4), .o(n_18120) );
na02f80 g552046 ( .a(n_17892), .b(n_17318), .o(n_18501) );
na02f80 g552047 ( .a(n_18119), .b(n_17575), .o(n_18725) );
na02f80 g552048 ( .a(n_16749), .b(n_17637), .o(n_17682) );
na02f80 g552049 ( .a(n_15993), .b(n_15651), .o(n_15652) );
na02f80 g552050 ( .a(n_16636), .b(n_16344), .o(n_16345) );
no02f80 g552051 ( .a(n_17715), .b(n_17409), .o(n_17410) );
no02f80 g552052 ( .a(n_16877), .b(n_16632), .o(n_16633) );
no02f80 g552053 ( .a(n_17890), .b(n_18151), .o(n_17891) );
no02f80 g552054 ( .a(n_17890), .b(n_17194), .o(n_18826) );
in01f80 g552055 ( .a(n_17106), .o(n_18025) );
na02f80 g552056 ( .a(n_16298), .b(n_14494), .o(n_17106) );
na02f80 g552057 ( .a(n_15990), .b(n_2739), .o(n_16638) );
na02f80 g552058 ( .a(n_17681), .b(FE_OFN450_n_17680), .o(n_18552) );
na02f80 g552059 ( .a(n_16866), .b(n_16865), .o(n_16867) );
no02f80 g552060 ( .a(n_17681), .b(n_17678), .o(n_17679) );
no02f80 g552061 ( .a(n_16873), .b(n_16865), .o(n_17792) );
na02f80 g552062 ( .a(n_17441), .b(n_17104), .o(n_17105) );
no02f80 g552063 ( .a(n_17407), .b(n_26552), .o(n_17408) );
na02f80 g552064 ( .a(n_17889), .b(n_17888), .o(n_18825) );
na02f80 g552065 ( .a(n_17889), .b(n_17692), .o(n_17677) );
na02f80 g552066 ( .a(n_17185), .b(n_17631), .o(n_17887) );
na02f80 g552067 ( .a(n_17188), .b(n_17628), .o(n_17886) );
na02f80 g552068 ( .a(n_17187), .b(n_17634), .o(n_17885) );
no02f80 g552069 ( .a(n_18117), .b(n_18116), .o(n_18118) );
no02f80 g552070 ( .a(n_18114), .b(n_18113), .o(n_18115) );
no02f80 g552071 ( .a(n_17883), .b(n_17882), .o(n_17884) );
no02f80 g552072 ( .a(n_17675), .b(n_17674), .o(n_17676) );
no02f80 g552073 ( .a(n_17880), .b(n_19129), .o(n_17881) );
no02f80 g552074 ( .a(n_17672), .b(n_17671), .o(n_17673) );
no02f80 g552075 ( .a(n_17669), .b(n_18822), .o(n_17670) );
no02f80 g552076 ( .a(n_17878), .b(n_17877), .o(n_17879) );
no02f80 g552077 ( .a(n_17667), .b(n_17666), .o(n_17668) );
no02f80 g552078 ( .a(n_17664), .b(n_17663), .o(n_17665) );
no02f80 g552079 ( .a(n_17661), .b(n_17660), .o(n_17662) );
no02f80 g552080 ( .a(n_17658), .b(n_17657), .o(n_17659) );
no02f80 g552081 ( .a(n_17655), .b(n_17654), .o(n_17656) );
no02f80 g552082 ( .a(n_17652), .b(n_17651), .o(n_17653) );
no02f80 g552083 ( .a(n_17649), .b(n_17648), .o(n_17650) );
no02f80 g552084 ( .a(n_17875), .b(n_17874), .o(n_17876) );
no02f80 g552085 ( .a(n_18111), .b(n_19737), .o(n_18112) );
no02f80 g552086 ( .a(n_17646), .b(n_17645), .o(n_17647) );
no02f80 g552087 ( .a(n_17643), .b(n_17642), .o(n_17644) );
no02f80 g552088 ( .a(n_17640), .b(n_17639), .o(n_17641) );
no02f80 g552089 ( .a(n_18109), .b(n_19414), .o(n_18110) );
na02f80 g552090 ( .a(n_16750), .b(FE_OFN48_n_17099), .o(n_17406) );
no02f80 g552091 ( .a(n_17873), .b(n_17411), .o(n_18548) );
na02f80 g552092 ( .a(n_17873), .b(n_17871), .o(n_17872) );
no02f80 g552093 ( .a(n_17404), .b(n_8892), .o(n_17405) );
no02f80 g552094 ( .a(n_17404), .b(n_17402), .o(n_17403) );
na02f80 g552095 ( .a(n_17118), .b(n_16863), .o(n_16864) );
na02f80 g552096 ( .a(n_17870), .b(n_16758), .o(n_18547) );
na02f80 g552097 ( .a(n_17870), .b(n_17868), .o(n_17869) );
no02f80 g552098 ( .a(n_17866), .b(n_17865), .o(n_17867) );
no02f80 g552099 ( .a(n_16862), .b(n_16246), .o(n_18028) );
ao12f80 g552100 ( .a(n_15573), .b(n_16838), .c(n_16269), .o(n_17161) );
oa12f80 g552101 ( .a(n_17637), .b(n_1024), .c(n_28928), .o(n_17638) );
oa12f80 g552102 ( .a(n_17637), .b(n_1791), .c(n_28607), .o(n_17636) );
oa12f80 g552103 ( .a(n_17634), .b(n_422), .c(FE_OFN352_n_4860), .o(n_17635) );
oa12f80 g552104 ( .a(n_17634), .b(n_21), .c(FE_OFN352_n_4860), .o(n_17633) );
oa12f80 g552105 ( .a(n_17631), .b(n_595), .c(FE_OFN122_n_27449), .o(n_17632) );
oa12f80 g552106 ( .a(n_17631), .b(n_1129), .c(FE_OFN1147_n_4860), .o(n_17630) );
oa12f80 g552107 ( .a(n_17628), .b(n_547), .c(FE_OFN350_n_4860), .o(n_17629) );
oa12f80 g552108 ( .a(n_17628), .b(n_1163), .c(FE_OFN350_n_4860), .o(n_17627) );
in01f80 g552109 ( .a(n_18032), .o(n_17626) );
na02f80 g552110 ( .a(n_16756), .b(n_17401), .o(n_18032) );
na02f80 g552111 ( .a(n_17109), .b(n_17401), .o(n_17103) );
no02f80 g552112 ( .a(n_16630), .b(n_16629), .o(n_16631) );
na02f80 g552113 ( .a(n_16343), .b(n_16629), .o(n_17801) );
in01f80 g552114 ( .a(n_17625), .o(n_18538) );
oa12f80 g552115 ( .a(n_17328), .b(n_16732), .c(n_15738), .o(n_17625) );
no02f80 g552116 ( .a(n_16862), .b(n_16860), .o(n_16861) );
oa12f80 g552117 ( .a(n_16759), .b(n_17254), .c(n_15284), .o(n_17624) );
in01f80 g552118 ( .a(n_18108), .o(n_19125) );
oa12f80 g552119 ( .a(n_16748), .b(n_17860), .c(n_16210), .o(n_18108) );
oa12f80 g552120 ( .a(n_13665), .b(n_16859), .c(n_14788), .o(n_17787) );
ao12f80 g552121 ( .a(n_14772), .b(n_16858), .c(n_15347), .o(n_17786) );
ao12f80 g552122 ( .a(n_14762), .b(n_16628), .c(n_15432), .o(n_17487) );
in01f80 g552123 ( .a(n_17623), .o(n_18539) );
oa12f80 g552124 ( .a(n_16540), .b(n_17400), .c(n_15894), .o(n_17623) );
ao12f80 g552125 ( .a(n_14641), .b(n_16627), .c(n_15404), .o(n_17486) );
ao12f80 g552126 ( .a(n_14735), .b(n_16626), .c(n_15394), .o(n_17485) );
oa12f80 g552127 ( .a(n_14374), .b(n_16625), .c(n_15139), .o(n_17484) );
ao12f80 g552128 ( .a(n_14705), .b(n_16624), .c(n_15382), .o(n_17483) );
ao12f80 g552129 ( .a(n_14681), .b(n_16623), .c(n_15364), .o(n_17482) );
ao12f80 g552130 ( .a(n_14320), .b(n_16857), .c(n_13146), .o(n_17785) );
in01f80 g552131 ( .a(n_17102), .o(n_18023) );
ao12f80 g552132 ( .a(n_12298), .b(n_16851), .c(n_12956), .o(n_17102) );
in01f80 g552133 ( .a(n_17864), .o(n_18819) );
oa12f80 g552134 ( .a(n_17558), .b(n_16914), .c(n_16684), .o(n_17864) );
ao12f80 g552135 ( .a(n_11452), .b(n_16342), .c(n_12445), .o(n_17160) );
in01f80 g552136 ( .a(n_17101), .o(n_18022) );
ao12f80 g552137 ( .a(n_11012), .b(n_16849), .c(n_12133), .o(n_17101) );
ao12f80 g552138 ( .a(n_16093), .b(n_17399), .c(n_16691), .o(n_18297) );
oa12f80 g552139 ( .a(n_12255), .b(n_16622), .c(n_12933), .o(n_17480) );
oa12f80 g552140 ( .a(n_11419), .b(n_16621), .c(n_12457), .o(n_17481) );
oa12f80 g552141 ( .a(n_13857), .b(FE_OFN1266_n_16620), .c(n_14904), .o(n_17479) );
oa12f80 g552142 ( .a(n_14800), .b(n_16856), .c(n_15433), .o(n_17784) );
oa12f80 g552143 ( .a(n_17189), .b(n_17227), .c(n_16686), .o(n_17863) );
oa12f80 g552144 ( .a(FE_OFN48_n_17099), .b(n_1966), .c(FE_OFN142_n_27449), .o(n_17100) );
oa12f80 g552145 ( .a(FE_OFN48_n_17099), .b(n_989), .c(FE_OFN142_n_27449), .o(n_17098) );
oa12f80 g552146 ( .a(n_17621), .b(n_971), .c(FE_OFN125_n_27449), .o(n_17622) );
oa12f80 g552147 ( .a(n_17397), .b(n_996), .c(FE_OFN135_n_27449), .o(n_17398) );
oa12f80 g552148 ( .a(FE_OFN1_n_17395), .b(n_976), .c(n_29261), .o(n_17396) );
oa12f80 g552149 ( .a(n_13972), .b(n_16619), .c(n_14946), .o(n_17478) );
ao12f80 g552150 ( .a(n_8294), .b(n_16855), .c(n_8936), .o(n_17783) );
ao22s80 g552151 ( .a(n_16465), .b(n_13023), .c(n_16272), .d(n_12895), .o(n_18296) );
oa12f80 g552152 ( .a(n_14458), .b(n_16854), .c(n_15011), .o(n_17782) );
oa12f80 g552153 ( .a(n_12287), .b(n_16853), .c(n_12504), .o(n_17780) );
ao12f80 g552154 ( .a(n_13652), .b(n_16618), .c(n_14749), .o(n_17477) );
oa12f80 g552155 ( .a(n_13176), .b(n_17394), .c(n_14370), .o(n_18295) );
ao12f80 g552156 ( .a(n_14438), .b(n_16617), .c(n_15164), .o(n_17476) );
ao12f80 g552157 ( .a(n_14409), .b(n_16852), .c(n_15152), .o(n_17781) );
ao12f80 g552158 ( .a(n_10657), .b(n_16341), .c(n_11793), .o(n_17159) );
oa12f80 g552159 ( .a(n_14251), .b(n_16616), .c(n_15098), .o(n_17475) );
oa12f80 g552160 ( .a(n_14244), .b(FE_OFN1236_n_16615), .c(n_15092), .o(n_17474) );
oa12f80 g552161 ( .a(n_15796), .b(n_17025), .c(n_16474), .o(n_17473) );
oa12f80 g552162 ( .a(n_14232), .b(n_16614), .c(n_15105), .o(n_17472) );
ao12f80 g552163 ( .a(n_14331), .b(n_16613), .c(n_15120), .o(n_17471) );
oa12f80 g552164 ( .a(n_10673), .b(n_16612), .c(n_11807), .o(n_17470) );
ao12f80 g552165 ( .a(n_8321), .b(n_16611), .c(n_8951), .o(n_17469) );
in01f80 g552166 ( .a(n_19468), .o(n_17620) );
oa12f80 g552167 ( .a(n_16955), .b(n_17393), .c(n_16954), .o(n_19468) );
in01f80 g552168 ( .a(n_19862), .o(n_17619) );
oa12f80 g552169 ( .a(n_17204), .b(n_17392), .c(n_17203), .o(n_19862) );
in01f80 g552170 ( .a(n_19465), .o(n_17862) );
oa12f80 g552171 ( .a(n_17206), .b(n_17618), .c(n_17205), .o(n_19465) );
in01f80 g552172 ( .a(n_19462), .o(n_17617) );
oa12f80 g552173 ( .a(n_16951), .b(n_17391), .c(n_16950), .o(n_19462) );
ao12f80 g552174 ( .a(n_17535), .b(n_17534), .c(n_17533), .o(n_18107) );
oa12f80 g552175 ( .a(n_17004), .b(n_17062), .c(n_17247), .o(n_18272) );
in01f80 g552176 ( .a(n_18223), .o(n_17097) );
oa12f80 g552177 ( .a(n_16340), .b(n_16628), .c(n_16339), .o(n_18223) );
ao12f80 g552178 ( .a(n_17034), .b(n_17033), .c(n_17032), .o(n_17616) );
ao12f80 g552179 ( .a(n_17543), .b(n_17845), .c(n_17542), .o(n_18106) );
oa12f80 g552180 ( .a(n_16996), .b(n_17266), .c(n_17061), .o(n_18251) );
ao22s80 g552181 ( .a(n_17860), .b(n_16923), .c(n_16898), .d(n_16922), .o(n_17861) );
ao12f80 g552182 ( .a(n_17071), .b(n_17374), .c(n_17070), .o(n_17615) );
oa12f80 g552183 ( .a(n_17240), .b(n_17239), .c(n_17238), .o(n_18513) );
oa12f80 g552184 ( .a(n_17003), .b(n_17060), .c(n_17242), .o(n_18271) );
oa12f80 g552185 ( .a(n_16999), .b(n_16998), .c(n_16997), .o(n_18266) );
oa12f80 g552186 ( .a(n_17313), .b(n_17312), .c(n_17546), .o(n_18495) );
in01f80 g552187 ( .a(n_18189), .o(n_17390) );
oa12f80 g552188 ( .a(n_16603), .b(n_16859), .c(n_16602), .o(n_18189) );
oa12f80 g552189 ( .a(n_17297), .b(n_17298), .c(n_17296), .o(n_18464) );
oa12f80 g552190 ( .a(n_16995), .b(n_16994), .c(n_16993), .o(n_18265) );
oa12f80 g552191 ( .a(n_17265), .b(n_17264), .c(n_17263), .o(n_18506) );
oa12f80 g552192 ( .a(n_16796), .b(n_16841), .c(n_16795), .o(n_17970) );
oa12f80 g552193 ( .a(n_17292), .b(n_17293), .c(n_17291), .o(n_18503) );
ao12f80 g552194 ( .a(n_17589), .b(n_17588), .c(n_17587), .o(n_18105) );
oa12f80 g552195 ( .a(n_17307), .b(n_17306), .c(n_17548), .o(n_18480) );
oa12f80 g552196 ( .a(n_16605), .b(n_16847), .c(n_16604), .o(n_18179) );
oa12f80 g552197 ( .a(n_17303), .b(n_17302), .c(n_17547), .o(n_18468) );
in01f80 g552198 ( .a(n_17940), .o(n_17770) );
ao12f80 g552199 ( .a(n_16318), .b(n_16617), .c(n_16317), .o(n_17940) );
in01f80 g552200 ( .a(n_18003), .o(n_17614) );
oa12f80 g552201 ( .a(n_16840), .b(n_16839), .c(n_16838), .o(n_18003) );
ao12f80 g552202 ( .a(n_17028), .b(n_17027), .c(n_18458), .o(n_17613) );
oa12f80 g552203 ( .a(n_17305), .b(n_17304), .c(n_17549), .o(n_18496) );
ao12f80 g552204 ( .a(n_17022), .b(n_17021), .c(n_17020), .o(n_17612) );
in01f80 g552205 ( .a(n_17948), .o(n_17751) );
ao12f80 g552206 ( .a(n_16312), .b(n_16614), .c(n_16311), .o(n_17948) );
ao12f80 g552207 ( .a(n_16816), .b(n_16815), .c(n_18209), .o(n_17389) );
in01f80 g552208 ( .a(n_17096), .o(n_18015) );
oa12f80 g552209 ( .a(n_16320), .b(n_16618), .c(n_16319), .o(n_17096) );
in01f80 g552210 ( .a(n_18232), .o(n_17095) );
oa12f80 g552211 ( .a(n_16338), .b(n_16627), .c(n_16337), .o(n_18232) );
ao12f80 g552212 ( .a(n_17019), .b(n_17018), .c(n_17017), .o(n_17611) );
in01f80 g552213 ( .a(n_17951), .o(n_17995) );
ao12f80 g552214 ( .a(n_16587), .b(n_16852), .c(n_16586), .o(n_17951) );
in01f80 g552215 ( .a(n_18219), .o(n_17094) );
oa12f80 g552216 ( .a(n_16336), .b(n_16626), .c(n_16335), .o(n_18219) );
ao12f80 g552217 ( .a(n_17290), .b(n_17289), .c(n_17288), .o(n_17859) );
in01f80 g552218 ( .a(n_18183), .o(n_17762) );
ao12f80 g552219 ( .a(n_16334), .b(n_16625), .c(n_16333), .o(n_18183) );
in01f80 g552220 ( .a(n_18212), .o(n_18462) );
ao12f80 g552221 ( .a(n_17036), .b(n_17394), .c(n_17035), .o(n_18212) );
ao12f80 g552222 ( .a(n_17287), .b(n_17286), .c(n_17285), .o(n_17858) );
ao12f80 g552223 ( .a(n_17284), .b(n_17283), .c(n_17282), .o(n_17857) );
in01f80 g552224 ( .a(n_18216), .o(n_17093) );
oa12f80 g552225 ( .a(n_16332), .b(n_16624), .c(n_16331), .o(n_18216) );
in01f80 g552226 ( .a(n_17728), .o(n_17092) );
oa12f80 g552227 ( .a(n_16322), .b(n_16619), .c(n_16321), .o(n_17728) );
ao12f80 g552228 ( .a(n_17538), .b(n_17537), .c(n_17536), .o(n_18104) );
in01f80 g552229 ( .a(n_18213), .o(n_17388) );
oa12f80 g552230 ( .a(n_16601), .b(n_16856), .c(n_16600), .o(n_18213) );
in01f80 g552231 ( .a(n_18229), .o(n_17091) );
oa12f80 g552232 ( .a(n_16330), .b(n_16623), .c(n_16329), .o(n_18229) );
ao12f80 g552233 ( .a(n_17016), .b(n_17015), .c(n_17014), .o(n_17610) );
oa12f80 g552234 ( .a(n_17251), .b(n_17250), .c(n_17249), .o(n_18514) );
in01f80 g552235 ( .a(FE_OFN602_n_17761), .o(n_18007) );
ao12f80 g552236 ( .a(n_16599), .b(n_16853), .c(n_16598), .o(n_17761) );
oa12f80 g552237 ( .a(n_16845), .b(n_16844), .c(x_in_1_14), .o(n_17990) );
ao12f80 g552238 ( .a(n_17281), .b(n_17280), .c(n_17279), .o(n_17856) );
oa12f80 g552239 ( .a(n_16793), .b(n_16831), .c(n_16792), .o(n_17989) );
ao22s80 g552240 ( .a(n_17393), .b(n_16224), .c(n_16666), .d(x_in_32_1), .o(n_18207) );
ao12f80 g552241 ( .a(n_16578), .b(n_16577), .c(n_16576), .o(n_17090) );
in01f80 g552242 ( .a(FE_OFN1017_n_17433), .o(n_17089) );
oa12f80 g552243 ( .a(n_16308), .b(n_16612), .c(n_16307), .o(n_17433) );
oa12f80 g552244 ( .a(n_16981), .b(n_17059), .c(n_17248), .o(n_18250) );
ao12f80 g552245 ( .a(n_17562), .b(n_17561), .c(n_17560), .o(n_18103) );
in01f80 g552246 ( .a(n_17725), .o(n_17088) );
oa12f80 g552247 ( .a(n_16310), .b(n_16613), .c(n_16309), .o(n_17725) );
ao12f80 g552248 ( .a(n_16812), .b(n_16811), .c(n_16810), .o(n_17387) );
ao12f80 g552249 ( .a(n_17278), .b(n_17277), .c(n_17276), .o(n_17855) );
ao22s80 g552250 ( .a(n_17392), .b(n_16221), .c(n_16664), .d(x_in_48_1), .o(n_18204) );
ao12f80 g552251 ( .a(n_17246), .b(n_17245), .c(n_17244), .o(n_17854) );
in01f80 g552252 ( .a(n_17716), .o(n_17718) );
ao12f80 g552253 ( .a(n_16305), .b(n_16611), .c(n_16304), .o(n_17716) );
in01f80 g552254 ( .a(n_17731), .o(n_17087) );
oa22f80 g552255 ( .a(n_16851), .b(n_13510), .c(n_15955), .d(n_13511), .o(n_17731) );
ao12f80 g552256 ( .a(n_16597), .b(n_16857), .c(n_16596), .o(n_18011) );
oa12f80 g552257 ( .a(n_17030), .b(n_17031), .c(n_17029), .o(n_18249) );
ao12f80 g552258 ( .a(n_17010), .b(n_17009), .c(n_17008), .o(n_17609) );
ao12f80 g552259 ( .a(n_17039), .b(n_17038), .c(n_17037), .o(n_17608) );
in01f80 g552260 ( .a(n_17769), .o(n_17386) );
oa12f80 g552261 ( .a(n_16589), .b(n_16854), .c(n_16588), .o(n_17769) );
oa12f80 g552262 ( .a(n_16788), .b(n_16837), .c(n_16787), .o(n_17982) );
in01f80 g552263 ( .a(n_18246), .o(n_17853) );
oa12f80 g552264 ( .a(n_17026), .b(n_17025), .c(n_17024), .o(n_18246) );
ao22s80 g552265 ( .a(n_17618), .b(n_16438), .c(n_16891), .d(x_in_40_1), .o(n_18459) );
in01f80 g552266 ( .a(n_18225), .o(n_17385) );
oa12f80 g552267 ( .a(n_16594), .b(n_16858), .c(n_16593), .o(n_18225) );
ao12f80 g552268 ( .a(n_17013), .b(n_17012), .c(n_17011), .o(n_17607) );
oa12f80 g552269 ( .a(n_16977), .b(n_16976), .c(n_16975), .o(n_18267) );
ao12f80 g552270 ( .a(n_16814), .b(n_16813), .c(n_18206), .o(n_17384) );
in01f80 g552271 ( .a(FE_OFN722_n_17438), .o(n_16850) );
oa12f80 g552272 ( .a(n_15987), .b(n_16342), .c(n_15986), .o(n_17438) );
oa12f80 g552273 ( .a(n_17527), .b(n_17526), .c(n_17525), .o(n_18757) );
ao12f80 g552274 ( .a(n_16809), .b(n_16808), .c(n_16807), .o(n_17383) );
oa12f80 g552275 ( .a(n_17311), .b(n_17310), .c(n_17545), .o(n_18494) );
ao12f80 g552276 ( .a(n_16806), .b(n_16805), .c(n_16804), .o(n_17382) );
in01f80 g552277 ( .a(n_17435), .o(n_17752) );
ao22s80 g552278 ( .a(n_15963), .b(n_12558), .c(n_16849), .d(n_12557), .o(n_17435) );
oa12f80 g552279 ( .a(n_16573), .b(n_16785), .c(n_16572), .o(n_17750) );
in01f80 g552280 ( .a(n_17460), .o(n_17086) );
oa12f80 g552281 ( .a(n_16316), .b(n_16616), .c(n_16315), .o(n_17460) );
ao12f80 g552282 ( .a(n_16784), .b(n_16783), .c(n_16782), .o(n_17381) );
ao12f80 g552283 ( .a(n_17275), .b(n_17274), .c(n_17273), .o(n_17852) );
ao12f80 g552284 ( .a(n_16818), .b(n_16817), .c(n_18203), .o(n_17380) );
oa12f80 g552285 ( .a(n_16829), .b(n_17369), .c(n_16828), .o(n_18708) );
ao12f80 g552286 ( .a(n_16583), .b(n_16582), .c(n_16581), .o(n_17085) );
in01f80 g552287 ( .a(n_16848), .o(n_17777) );
oa12f80 g552288 ( .a(n_15985), .b(n_16341), .c(n_15984), .o(n_16848) );
in01f80 g552289 ( .a(n_17459), .o(n_17084) );
oa12f80 g552290 ( .a(n_16314), .b(FE_OFN1236_n_16615), .c(n_16313), .o(n_17459) );
in01f80 g552291 ( .a(n_17961), .o(n_17958) );
ao12f80 g552292 ( .a(n_16591), .b(n_16855), .c(n_16590), .o(n_17961) );
in01f80 g552293 ( .a(n_18490), .o(n_18102) );
oa12f80 g552294 ( .a(n_17327), .b(n_17399), .c(n_17326), .o(n_18490) );
oa12f80 g552295 ( .a(n_17523), .b(n_17819), .c(n_17522), .o(n_18760) );
ao12f80 g552296 ( .a(n_17272), .b(n_17271), .c(n_17270), .o(n_17851) );
ao12f80 g552297 ( .a(n_17007), .b(n_17006), .c(n_17005), .o(n_17606) );
ao12f80 g552298 ( .a(n_16825), .b(n_17080), .c(n_16824), .o(n_17379) );
in01f80 g552299 ( .a(n_17458), .o(n_17743) );
ao12f80 g552300 ( .a(n_16328), .b(n_16622), .c(n_16327), .o(n_17458) );
ao12f80 g552301 ( .a(n_17359), .b(n_17358), .c(n_17357), .o(n_17850) );
oa12f80 g552302 ( .a(n_17817), .b(n_17818), .c(n_17816), .o(n_19080) );
ao12f80 g552303 ( .a(n_16823), .b(n_17075), .c(n_16822), .o(n_17378) );
ao22s80 g552304 ( .a(n_16728), .b(n_17400), .c(n_16727), .d(n_16489), .o(n_17605) );
ao22s80 g552305 ( .a(n_17391), .b(n_16227), .c(n_16661), .d(x_in_52_1), .o(n_18210) );
oa12f80 g552306 ( .a(n_17301), .b(n_17300), .c(n_17544), .o(n_18471) );
ao12f80 g552307 ( .a(n_17269), .b(n_17268), .c(n_17267), .o(n_17849) );
oa12f80 g552308 ( .a(n_17309), .b(n_17308), .c(n_17550), .o(n_18477) );
in01f80 g552309 ( .a(n_17738), .o(n_17377) );
oa12f80 g552310 ( .a(n_16585), .b(n_16584), .c(n_16607), .o(n_17738) );
ao12f80 g552311 ( .a(n_17294), .b(n_17366), .c(n_17295), .o(n_17848) );
in01f80 g552312 ( .a(n_17457), .o(n_17740) );
ao12f80 g552313 ( .a(n_16324), .b(n_16621), .c(n_16323), .o(n_17457) );
in01f80 g552314 ( .a(n_17456), .o(n_17083) );
oa12f80 g552315 ( .a(n_16326), .b(FE_OFN1266_n_16620), .c(n_16325), .o(n_17456) );
oa12f80 g552316 ( .a(n_16820), .b(n_17074), .c(n_16819), .o(n_18430) );
oa22f80 g552317 ( .a(n_16464), .b(FE_OFN201_n_29637), .c(n_51), .d(FE_OFN1146_n_4860), .o(n_17376) );
oa22f80 g552318 ( .a(FE_OFN596_n_16896), .b(FE_OFN410_n_28303), .c(n_191), .d(n_27709), .o(n_17847) );
oa22f80 g552319 ( .a(n_15951), .b(n_15949), .c(n_16847), .d(n_15948), .o(n_17788) );
oa22f80 g552320 ( .a(n_17533), .b(FE_OFN409_n_28303), .c(n_1335), .d(FE_OFN288_n_29266), .o(n_17082) );
oa22f80 g552321 ( .a(n_16665), .b(n_29683), .c(n_984), .d(n_29264), .o(n_17604) );
oa22f80 g552322 ( .a(n_16670), .b(FE_OFN264_n_4280), .c(n_97), .d(FE_OFN357_n_4860), .o(n_17603) );
oa22f80 g552323 ( .a(n_16669), .b(n_28303), .c(n_1549), .d(n_27449), .o(n_17602) );
oa22f80 g552324 ( .a(FE_OFN1015_n_16571), .b(FE_OFN235_n_4162), .c(n_1737), .d(n_29104), .o(n_16846) );
oa22f80 g552325 ( .a(n_16306), .b(FE_OFN405_n_28303), .c(n_519), .d(FE_OFN92_n_27449), .o(n_16610) );
oa22f80 g552326 ( .a(n_17080), .b(FE_OFN307_n_3069), .c(n_152), .d(FE_OFN99_n_27449), .o(n_17081) );
oa22f80 g552327 ( .a(n_17845), .b(n_28608), .c(n_865), .d(FE_OFN102_n_27449), .o(n_17846) );
oa22f80 g552328 ( .a(n_17374), .b(FE_OFN416_n_28303), .c(n_1759), .d(FE_OFN108_n_27449), .o(n_17375) );
oa22f80 g552329 ( .a(n_16454), .b(FE_OFN181_n_27681), .c(n_939), .d(FE_OFN1121_rst), .o(n_17373) );
oa22f80 g552330 ( .a(n_16239), .b(n_27681), .c(n_797), .d(FE_OFN98_n_27449), .o(n_17079) );
oa22f80 g552331 ( .a(n_16892), .b(FE_OFN240_n_4162), .c(n_254), .d(FE_OFN78_n_27012), .o(n_17844) );
oa22f80 g552332 ( .a(n_16452), .b(FE_OFN413_n_28303), .c(n_1220), .d(FE_OFN1121_rst), .o(n_17372) );
oa22f80 g552333 ( .a(n_16450), .b(FE_OFN307_n_3069), .c(n_85), .d(FE_OFN355_n_4860), .o(n_17371) );
oa22f80 g552334 ( .a(n_16575), .b(FE_OFN258_n_4280), .c(n_554), .d(FE_OFN1121_rst), .o(n_16609) );
oa22f80 g552335 ( .a(n_16447), .b(FE_OFN251_n_4162), .c(n_338), .d(rst), .o(n_17370) );
oa22f80 g552336 ( .a(n_16607), .b(FE_OFN251_n_4162), .c(n_642), .d(FE_OFN330_n_4860), .o(n_16608) );
ao22s80 g552337 ( .a(n_16446), .b(n_16233), .c(n_17369), .d(n_16232), .o(n_18299) );
oa22f80 g552338 ( .a(n_16463), .b(n_4162), .c(n_196), .d(FE_OFN116_n_27449), .o(n_17368) );
oa22f80 g552339 ( .a(n_16236), .b(FE_OFN258_n_4280), .c(n_1514), .d(FE_OFN352_n_4860), .o(n_17078) );
oa22f80 g552340 ( .a(n_16231), .b(FE_OFN249_n_4162), .c(n_943), .d(FE_OFN1110_rst), .o(n_17077) );
oa22f80 g552341 ( .a(n_17366), .b(FE_OFN256_n_4280), .c(n_1035), .d(FE_OFN336_n_4860), .o(n_17367) );
oa22f80 g552342 ( .a(n_16442), .b(n_4280), .c(n_969), .d(FE_OFN1112_rst), .o(n_17365) );
oa22f80 g552343 ( .a(n_16456), .b(FE_OFN296_n_3069), .c(n_1027), .d(n_28928), .o(n_17364) );
oa22f80 g552344 ( .a(n_16660), .b(FE_OFN251_n_4162), .c(n_1031), .d(FE_OFN1111_rst), .o(n_17601) );
oa22f80 g552345 ( .a(n_17075), .b(FE_OFN247_n_4162), .c(n_1305), .d(FE_OFN80_n_27012), .o(n_17076) );
oa22f80 g552346 ( .a(n_16659), .b(FE_OFN311_n_3069), .c(n_1016), .d(n_29068), .o(n_17600) );
ao22s80 g552347 ( .a(n_16905), .b(n_16451), .c(x_out_51_19), .d(FE_OFN274_n_16893), .o(n_17843) );
ao22s80 g552348 ( .a(n_16786), .b(n_16694), .c(x_out_38_19), .d(FE_OFN271_n_16028), .o(n_17363) );
ao22s80 g552349 ( .a(n_16695), .b(n_16580), .c(x_out_43_19), .d(FE_OFN280_n_16656), .o(n_17362) );
oa22f80 g552350 ( .a(n_16235), .b(n_15945), .c(n_17074), .d(n_15944), .o(n_18027) );
na02f80 g552384 ( .a(n_16844), .b(x_in_1_14), .o(n_16845) );
na02f80 g552385 ( .a(n_17526), .b(x_in_60_2), .o(n_17910) );
in01f80 g552386 ( .a(n_17360), .o(n_17361) );
no02f80 g552387 ( .a(n_17526), .b(x_in_60_2), .o(n_17360) );
in01f80 g552388 ( .a(n_16842), .o(n_16843) );
no02f80 g552389 ( .a(n_16606), .b(x_in_8_5), .o(n_16842) );
na02f80 g552390 ( .a(n_17325), .b(x_in_46_2), .o(n_18130) );
in01f80 g552391 ( .a(n_17072), .o(n_17073) );
no02f80 g552392 ( .a(n_16830), .b(x_in_56_4), .o(n_17072) );
na02f80 g552393 ( .a(n_16628), .b(n_16339), .o(n_16340) );
in01f80 g552394 ( .a(n_17598), .o(n_17599) );
no02f80 g552395 ( .a(n_17319), .b(x_in_2_2), .o(n_17598) );
no02f80 g552396 ( .a(n_17358), .b(n_17357), .o(n_17359) );
in01f80 g552397 ( .a(n_17596), .o(n_17597) );
no02f80 g552398 ( .a(n_17356), .b(x_in_34_2), .o(n_17596) );
na02f80 g552399 ( .a(n_17356), .b(x_in_34_2), .o(n_18142) );
na02f80 g552400 ( .a(n_16606), .b(x_in_8_5), .o(n_17412) );
no02f80 g552401 ( .a(n_16229), .b(n_16822), .o(n_17739) );
na02f80 g552402 ( .a(n_17595), .b(x_in_18_2), .o(n_18398) );
in01f80 g552403 ( .a(n_17840), .o(n_17841) );
no02f80 g552404 ( .a(n_17595), .b(x_in_18_2), .o(n_17840) );
no02f80 g552405 ( .a(n_17374), .b(n_17070), .o(n_17071) );
in01f80 g552406 ( .a(n_17354), .o(n_17355) );
no02f80 g552407 ( .a(n_17066), .b(x_in_26_2), .o(n_17354) );
na02f80 g552408 ( .a(n_17594), .b(x_in_50_2), .o(n_18407) );
in01f80 g552409 ( .a(n_17838), .o(n_17839) );
no02f80 g552410 ( .a(n_17594), .b(x_in_50_2), .o(n_17838) );
na02f80 g552411 ( .a(n_17051), .b(x_in_56_3), .o(n_17911) );
na02f80 g552412 ( .a(n_16847), .b(n_16604), .o(n_16605) );
na02f80 g552413 ( .a(n_17264), .b(x_in_6_2), .o(n_17699) );
in01f80 g552414 ( .a(n_17068), .o(n_17069) );
no02f80 g552415 ( .a(n_17264), .b(x_in_6_2), .o(n_17068) );
na02f80 g552416 ( .a(n_17353), .b(x_in_10_2), .o(n_18141) );
in01f80 g552417 ( .a(n_17592), .o(n_17593) );
no02f80 g552418 ( .a(n_17353), .b(x_in_10_2), .o(n_17592) );
na02f80 g552419 ( .a(n_17352), .b(x_in_42_2), .o(n_18138) );
in01f80 g552420 ( .a(n_17590), .o(n_17591) );
no02f80 g552421 ( .a(n_17352), .b(x_in_42_2), .o(n_17590) );
na02f80 g552422 ( .a(n_16859), .b(n_16602), .o(n_16603) );
na02f80 g552423 ( .a(n_16461), .b(n_16798), .o(n_17067) );
na02f80 g552424 ( .a(n_17341), .b(x_in_58_2), .o(n_18137) );
na02f80 g552425 ( .a(n_17066), .b(x_in_26_2), .o(n_17895) );
na02f80 g552426 ( .a(n_16841), .b(x_in_52_2), .o(n_17697) );
in01f80 g552427 ( .a(n_17064), .o(n_17065) );
no02f80 g552428 ( .a(n_16841), .b(x_in_52_2), .o(n_17064) );
na02f80 g552429 ( .a(n_17063), .b(x_in_38_3), .o(n_17897) );
in01f80 g552430 ( .a(n_17350), .o(n_17351) );
no02f80 g552431 ( .a(n_17063), .b(x_in_38_3), .o(n_17350) );
no02f80 g552432 ( .a(n_17588), .b(n_17587), .o(n_17589) );
in01f80 g552433 ( .a(n_17585), .o(n_17586) );
na02f80 g552434 ( .a(n_17349), .b(n_16747), .o(n_17585) );
na02f80 g552435 ( .a(n_17348), .b(x_in_22_2), .o(n_18122) );
in01f80 g552436 ( .a(n_17583), .o(n_17584) );
no02f80 g552437 ( .a(n_17348), .b(x_in_22_2), .o(n_17583) );
in01f80 g552438 ( .a(n_17836), .o(n_17837) );
no02f80 g552439 ( .a(n_17555), .b(x_in_54_3), .o(n_17836) );
na02f80 g552440 ( .a(n_17347), .b(x_in_54_2), .o(n_18123) );
in01f80 g552441 ( .a(n_17581), .o(n_17582) );
no02f80 g552442 ( .a(n_17347), .b(x_in_54_2), .o(n_17581) );
na02f80 g552443 ( .a(n_17062), .b(x_in_2_3), .o(n_17896) );
in01f80 g552444 ( .a(n_17345), .o(n_17346) );
no02f80 g552445 ( .a(n_17062), .b(x_in_2_3), .o(n_17345) );
na02f80 g552446 ( .a(n_17580), .b(x_in_22_3), .o(n_18406) );
na02f80 g552447 ( .a(n_16839), .b(n_16838), .o(n_16840) );
in01f80 g552448 ( .a(n_17834), .o(n_17835) );
no02f80 g552449 ( .a(n_17580), .b(x_in_22_3), .o(n_17834) );
na02f80 g552450 ( .a(n_16837), .b(x_in_40_2), .o(n_17693) );
na02f80 g552451 ( .a(n_17344), .b(x_in_14_2), .o(n_18132) );
in01f80 g552452 ( .a(n_17578), .o(n_17579) );
no02f80 g552453 ( .a(n_17344), .b(x_in_14_2), .o(n_17578) );
na02f80 g552454 ( .a(n_17343), .b(x_in_30_2), .o(n_18133) );
in01f80 g552455 ( .a(n_17576), .o(n_17577) );
no02f80 g552456 ( .a(n_17343), .b(x_in_30_2), .o(n_17576) );
na02f80 g552457 ( .a(n_17342), .b(x_in_62_2), .o(n_18119) );
in01f80 g552458 ( .a(n_17574), .o(n_17575) );
no02f80 g552459 ( .a(n_17342), .b(x_in_62_2), .o(n_17574) );
in01f80 g552460 ( .a(n_17572), .o(n_17573) );
no02f80 g552461 ( .a(n_17341), .b(x_in_58_2), .o(n_17572) );
in01f80 g552462 ( .a(n_17339), .o(n_17340) );
no02f80 g552463 ( .a(n_17061), .b(x_in_26_3), .o(n_17339) );
in01f80 g552464 ( .a(n_17570), .o(n_17571) );
no02f80 g552465 ( .a(n_17819), .b(x_in_36_2), .o(n_17570) );
na02f80 g552466 ( .a(n_16627), .b(n_16337), .o(n_16338) );
na02f80 g552467 ( .a(n_17569), .b(x_in_14_3), .o(n_18404) );
in01f80 g552468 ( .a(n_17832), .o(n_17833) );
no02f80 g552469 ( .a(n_17569), .b(x_in_14_3), .o(n_17832) );
na02f80 g552470 ( .a(n_17060), .b(x_in_34_3), .o(n_17907) );
in01f80 g552471 ( .a(n_17337), .o(n_17338) );
no02f80 g552472 ( .a(n_17060), .b(x_in_34_3), .o(n_17337) );
na02f80 g552473 ( .a(n_16626), .b(n_16335), .o(n_16336) );
na02f80 g552474 ( .a(n_17568), .b(x_in_46_3), .o(n_18403) );
in01f80 g552475 ( .a(n_17830), .o(n_17831) );
no02f80 g552476 ( .a(n_17568), .b(x_in_46_3), .o(n_17830) );
no02f80 g552477 ( .a(n_16625), .b(n_16333), .o(n_16334) );
na02f80 g552478 ( .a(n_17059), .b(x_in_16_3), .o(n_17906) );
in01f80 g552479 ( .a(n_17335), .o(n_17336) );
no02f80 g552480 ( .a(n_17059), .b(x_in_16_3), .o(n_17335) );
na02f80 g552481 ( .a(n_16624), .b(n_16331), .o(n_16332) );
na02f80 g552482 ( .a(n_17567), .b(x_in_30_3), .o(n_18402) );
in01f80 g552483 ( .a(n_17828), .o(n_17829) );
no02f80 g552484 ( .a(n_17567), .b(x_in_30_3), .o(n_17828) );
na02f80 g552485 ( .a(n_17250), .b(x_in_18_3), .o(n_17694) );
in01f80 g552486 ( .a(n_17057), .o(n_17058) );
no02f80 g552487 ( .a(n_17250), .b(x_in_18_3), .o(n_17057) );
na02f80 g552488 ( .a(n_16856), .b(n_16600), .o(n_16601) );
na02f80 g552489 ( .a(n_16623), .b(n_16329), .o(n_16330) );
na02f80 g552490 ( .a(n_17566), .b(x_in_62_3), .o(n_18401) );
na02f80 g552491 ( .a(n_17565), .b(x_in_12_3), .o(n_18400) );
in01f80 g552492 ( .a(n_17826), .o(n_17827) );
no02f80 g552493 ( .a(n_17566), .b(x_in_62_3), .o(n_17826) );
in01f80 g552494 ( .a(n_17824), .o(n_17825) );
no02f80 g552495 ( .a(n_17565), .b(x_in_12_3), .o(n_17824) );
no02f80 g552496 ( .a(n_16853), .b(n_16598), .o(n_16599) );
in01f80 g552497 ( .a(n_17563), .o(n_17564) );
na02f80 g552498 ( .a(n_17334), .b(n_16738), .o(n_17563) );
na02f80 g552499 ( .a(n_16836), .b(x_in_0_12), .o(n_17696) );
in01f80 g552500 ( .a(n_17055), .o(n_17056) );
no02f80 g552501 ( .a(n_16836), .b(x_in_0_12), .o(n_17055) );
no02f80 g552502 ( .a(n_16457), .b(n_17070), .o(n_18006) );
na02f80 g552503 ( .a(n_17054), .b(x_in_16_2), .o(n_17901) );
in01f80 g552504 ( .a(n_17332), .o(n_17333) );
no02f80 g552505 ( .a(n_17054), .b(x_in_16_2), .o(n_17332) );
no02f80 g552506 ( .a(n_17561), .b(n_17560), .o(n_17562) );
na02f80 g552507 ( .a(n_17561), .b(n_16753), .o(n_18128) );
na02f80 g552508 ( .a(n_17239), .b(x_in_50_3), .o(n_17417) );
in01f80 g552509 ( .a(n_16834), .o(n_16835) );
no02f80 g552510 ( .a(n_17239), .b(x_in_50_3), .o(n_16834) );
no02f80 g552511 ( .a(n_16230), .b(n_16824), .o(n_17742) );
no02f80 g552512 ( .a(n_16857), .b(n_16596), .o(n_16597) );
na02f80 g552513 ( .a(n_17559), .b(x_in_8_4), .o(n_18399) );
in01f80 g552514 ( .a(n_17822), .o(n_17823) );
no02f80 g552515 ( .a(n_17559), .b(x_in_8_4), .o(n_17822) );
na02f80 g552516 ( .a(n_17558), .b(n_16915), .o(n_18125) );
na02f80 g552517 ( .a(n_16595), .b(x_in_44_3), .o(n_17413) );
in01f80 g552518 ( .a(n_16832), .o(n_16833) );
no02f80 g552519 ( .a(n_16595), .b(x_in_44_3), .o(n_16832) );
na02f80 g552520 ( .a(n_16831), .b(x_in_32_2), .o(n_17689) );
in01f80 g552521 ( .a(n_17052), .o(n_17053) );
no02f80 g552522 ( .a(n_16831), .b(x_in_32_2), .o(n_17052) );
no02f80 g552523 ( .a(n_16622), .b(n_16327), .o(n_16328) );
na02f80 g552524 ( .a(n_16342), .b(n_15986), .o(n_15987) );
na02f80 g552525 ( .a(n_16858), .b(n_16593), .o(n_16594) );
na02f80 g552526 ( .a(n_17061), .b(x_in_26_3), .o(n_17894) );
in01f80 g552527 ( .a(n_17556), .o(n_17557) );
na02f80 g552528 ( .a(n_17331), .b(n_16745), .o(n_17556) );
in01f80 g552529 ( .a(n_17329), .o(n_17330) );
no02f80 g552530 ( .a(n_17051), .b(x_in_56_3), .o(n_17329) );
na02f80 g552531 ( .a(n_16976), .b(x_in_10_3), .o(n_17684) );
in01f80 g552532 ( .a(n_17049), .o(n_17050) );
no02f80 g552533 ( .a(n_16976), .b(x_in_10_3), .o(n_17049) );
na02f80 g552534 ( .a(n_17328), .b(n_16733), .o(n_17866) );
in01f80 g552535 ( .a(n_17047), .o(n_17048) );
no02f80 g552536 ( .a(n_16837), .b(x_in_40_2), .o(n_17047) );
na02f80 g552537 ( .a(n_16830), .b(x_in_56_4), .o(n_17698) );
na02f80 g552538 ( .a(n_17369), .b(n_16828), .o(n_16829) );
na02f80 g552539 ( .a(n_17816), .b(x_in_20_2), .o(n_18408) );
in01f80 g552540 ( .a(n_17820), .o(n_17821) );
no02f80 g552541 ( .a(n_17816), .b(x_in_20_2), .o(n_17820) );
in01f80 g552542 ( .a(n_16826), .o(n_16827) );
na02f80 g552543 ( .a(n_16592), .b(n_15976), .o(n_16826) );
na02f80 g552544 ( .a(n_16998), .b(x_in_42_3), .o(n_17683) );
in01f80 g552545 ( .a(n_17045), .o(n_17046) );
no02f80 g552546 ( .a(n_16998), .b(x_in_42_3), .o(n_17045) );
na02f80 g552547 ( .a(n_17555), .b(x_in_54_3), .o(n_18405) );
na02f80 g552548 ( .a(n_17399), .b(n_17326), .o(n_17327) );
no02f80 g552549 ( .a(n_17080), .b(n_16824), .o(n_16825) );
in01f80 g552550 ( .a(n_17553), .o(n_17554) );
no02f80 g552551 ( .a(n_17325), .b(x_in_46_2), .o(n_17553) );
in01f80 g552552 ( .a(n_17323), .o(n_17324) );
na02f80 g552553 ( .a(n_17044), .b(n_16543), .o(n_17323) );
na02f80 g552554 ( .a(n_17819), .b(x_in_36_2), .o(n_18143) );
no02f80 g552555 ( .a(n_17075), .b(n_16822), .o(n_16823) );
na02f80 g552556 ( .a(n_17322), .b(x_in_12_2), .o(n_18131) );
in01f80 g552557 ( .a(n_17551), .o(n_17552) );
no02f80 g552558 ( .a(n_17322), .b(x_in_12_2), .o(n_17551) );
na02f80 g552559 ( .a(n_17043), .b(x_in_44_2), .o(n_17912) );
in01f80 g552560 ( .a(n_17320), .o(n_17321) );
no02f80 g552561 ( .a(n_17043), .b(x_in_44_2), .o(n_17320) );
na02f80 g552562 ( .a(n_17319), .b(x_in_2_2), .o(n_18134) );
na02f80 g552563 ( .a(n_17042), .b(x_in_28_3), .o(n_17892) );
in01f80 g552564 ( .a(n_17317), .o(n_17318) );
no02f80 g552565 ( .a(n_17042), .b(x_in_28_3), .o(n_17317) );
na02f80 g552566 ( .a(FE_OFN1266_n_16620), .b(n_16325), .o(n_16326) );
na02f80 g552567 ( .a(n_16994), .b(x_in_58_3), .o(n_17700) );
no02f80 g552568 ( .a(n_16621), .b(n_16323), .o(n_16324) );
in01f80 g552569 ( .a(n_17040), .o(n_17041) );
no02f80 g552570 ( .a(n_16994), .b(x_in_58_3), .o(n_17040) );
oa12f80 g552571 ( .a(n_16459), .b(n_16405), .c(FE_OFN253_n_4280), .o(n_17316) );
oa12f80 g552572 ( .a(n_16458), .b(n_16403), .c(FE_OFN303_n_3069), .o(n_17315) );
oa12f80 g552573 ( .a(n_15947), .b(n_15888), .c(FE_OFN416_n_28303), .o(n_16821) );
oa12f80 g552574 ( .a(n_16449), .b(n_16404), .c(FE_OFN258_n_4280), .o(n_17314) );
na02f80 g552575 ( .a(n_16619), .b(n_16321), .o(n_16322) );
na02f80 g552576 ( .a(n_16844), .b(n_892), .o(n_17407) );
na02f80 g552577 ( .a(n_17074), .b(n_16819), .o(n_16820) );
no02f80 g552578 ( .a(n_16855), .b(n_16590), .o(n_16591) );
no02f80 g552579 ( .a(n_17038), .b(n_17037), .o(n_17039) );
na02f80 g552580 ( .a(n_17038), .b(n_16929), .o(n_17890) );
ao12f80 g552581 ( .a(n_3876), .b(n_15257), .c(n_4610), .o(n_15990) );
na02f80 g552582 ( .a(n_16618), .b(n_16319), .o(n_16320) );
na02f80 g552583 ( .a(n_16854), .b(n_16588), .o(n_16589) );
no02f80 g552584 ( .a(n_17394), .b(n_17035), .o(n_17036) );
no02f80 g552585 ( .a(n_16617), .b(n_16317), .o(n_16318) );
no02f80 g552586 ( .a(n_16852), .b(n_16586), .o(n_16587) );
na02f80 g552587 ( .a(n_16341), .b(n_15984), .o(n_15985) );
no02f80 g552588 ( .a(n_17033), .b(n_17032), .o(n_17034) );
no02f80 g552589 ( .a(n_17566), .b(n_17550), .o(n_18228) );
no02f80 g552590 ( .a(n_17569), .b(n_17549), .o(n_18231) );
no02f80 g552591 ( .a(n_17580), .b(n_17548), .o(n_18227) );
na02f80 g552592 ( .a(n_17312), .b(n_17546), .o(n_17313) );
no02f80 g552593 ( .a(n_17555), .b(n_17547), .o(n_18222) );
no02f80 g552594 ( .a(n_17568), .b(n_17546), .o(n_18218) );
no02f80 g552595 ( .a(n_17567), .b(n_17545), .o(n_18221) );
na02f80 g552596 ( .a(n_17310), .b(n_17545), .o(n_17311) );
na02f80 g552597 ( .a(n_17308), .b(n_17550), .o(n_17309) );
no02f80 g552598 ( .a(n_17033), .b(n_16049), .o(n_17681) );
no02f80 g552599 ( .a(n_17031), .b(n_16606), .o(n_17733) );
na02f80 g552600 ( .a(n_17031), .b(n_17029), .o(n_17030) );
na02f80 g552601 ( .a(n_17306), .b(n_17548), .o(n_17307) );
na02f80 g552602 ( .a(n_17304), .b(n_17549), .o(n_17305) );
na02f80 g552603 ( .a(n_17302), .b(n_17547), .o(n_17303) );
no02f80 g552604 ( .a(n_17565), .b(n_17544), .o(n_18215) );
na02f80 g552605 ( .a(n_17300), .b(n_17544), .o(n_17301) );
na02f80 g552606 ( .a(n_17299), .b(n_16911), .o(n_22092) );
na02f80 g552607 ( .a(n_16616), .b(n_16315), .o(n_16316) );
na02f80 g552608 ( .a(FE_OFN1236_n_16615), .b(n_16313), .o(n_16314) );
no02f80 g552609 ( .a(n_17845), .b(n_17542), .o(n_17543) );
no02f80 g552610 ( .a(n_16895), .b(n_17542), .o(n_18461) );
na02f80 g552611 ( .a(n_16584), .b(n_16607), .o(n_16585) );
no02f80 g552612 ( .a(n_16584), .b(n_16595), .o(n_17889) );
no02f80 g552613 ( .a(n_16817), .b(n_18203), .o(n_16818) );
no02f80 g552614 ( .a(n_17027), .b(n_18458), .o(n_17028) );
no02f80 g552615 ( .a(n_16815), .b(n_18209), .o(n_16816) );
no02f80 g552616 ( .a(n_16813), .b(n_18206), .o(n_16814) );
na02f80 g552617 ( .a(n_17025), .b(n_17024), .o(n_17026) );
no02f80 g552618 ( .a(n_16614), .b(n_16311), .o(n_16312) );
na02f80 g552619 ( .a(n_16613), .b(n_16309), .o(n_16310) );
na02f80 g552620 ( .a(n_17298), .b(n_15728), .o(n_17873) );
na02f80 g552621 ( .a(n_17298), .b(n_17296), .o(n_17297) );
na02f80 g552622 ( .a(n_16890), .b(FE_OFN46_n_17233), .o(n_17541) );
na02f80 g552623 ( .a(n_16888), .b(n_17258), .o(n_17540) );
no02f80 g552624 ( .a(n_16443), .b(n_17295), .o(n_17960) );
no02f80 g552625 ( .a(n_17366), .b(n_17295), .o(n_17294) );
na02f80 g552626 ( .a(n_16612), .b(n_16307), .o(n_16308) );
na02f80 g552627 ( .a(n_16889), .b(n_17261), .o(n_17539) );
no02f80 g552628 ( .a(n_16582), .b(n_16581), .o(n_16583) );
na02f80 g552629 ( .a(n_16306), .b(n_16581), .o(n_17444) );
oa12f80 g552630 ( .a(n_16460), .b(n_15884), .c(FE_OFN303_n_3069), .o(n_17023) );
no02f80 g552631 ( .a(n_16611), .b(n_16304), .o(n_16305) );
no02f80 g552632 ( .a(n_17293), .b(n_16553), .o(n_17870) );
na02f80 g552633 ( .a(n_17293), .b(n_17291), .o(n_17292) );
no02f80 g552634 ( .a(n_17021), .b(n_17020), .o(n_17022) );
no02f80 g552635 ( .a(n_17018), .b(n_17017), .o(n_17019) );
no02f80 g552636 ( .a(n_17289), .b(n_17288), .o(n_17290) );
no02f80 g552637 ( .a(n_17286), .b(n_17285), .o(n_17287) );
no02f80 g552638 ( .a(n_17283), .b(n_17282), .o(n_17284) );
no02f80 g552639 ( .a(n_17537), .b(n_17536), .o(n_17538) );
no02f80 g552640 ( .a(n_17015), .b(n_17014), .o(n_17016) );
no02f80 g552641 ( .a(n_17280), .b(n_17279), .o(n_17281) );
no02f80 g552642 ( .a(n_17277), .b(n_17276), .o(n_17278) );
no02f80 g552643 ( .a(n_16811), .b(n_16810), .o(n_16812) );
no02f80 g552644 ( .a(n_17012), .b(n_17011), .o(n_17013) );
no02f80 g552645 ( .a(n_17009), .b(n_17008), .o(n_17010) );
no02f80 g552646 ( .a(n_16808), .b(n_16807), .o(n_16809) );
no02f80 g552647 ( .a(n_16805), .b(n_16804), .o(n_16806) );
no02f80 g552648 ( .a(n_17006), .b(n_17005), .o(n_17007) );
no02f80 g552649 ( .a(n_17274), .b(n_17273), .o(n_17275) );
no02f80 g552650 ( .a(n_17271), .b(n_17270), .o(n_17272) );
no02f80 g552651 ( .a(n_17268), .b(n_17267), .o(n_17269) );
na02f80 g552652 ( .a(n_16238), .b(FE_OFN1120_rst), .o(n_17397) );
na02f80 g552653 ( .a(n_16801), .b(FE_OFN1114_rst), .o(n_17395) );
na02f80 g552654 ( .a(n_16448), .b(rst), .o(n_17621) );
no02f80 g552655 ( .a(n_17534), .b(n_17533), .o(n_17535) );
na02f80 g552656 ( .a(n_17062), .b(n_17247), .o(n_17004) );
na02f80 g552657 ( .a(n_17060), .b(n_17242), .o(n_17003) );
in01f80 g552658 ( .a(n_17002), .o(n_17931) );
oa12f80 g552659 ( .a(n_16424), .b(n_16803), .c(n_15683), .o(n_17002) );
oa12f80 g552660 ( .a(n_16991), .b(n_1527), .c(FE_OFN69_n_27012), .o(n_17001) );
oa12f80 g552661 ( .a(n_16779), .b(n_1441), .c(FE_OFN1120_rst), .o(n_16802) );
no02f80 g552662 ( .a(n_17250), .b(n_16649), .o(n_17730) );
in01f80 g552663 ( .a(n_17000), .o(n_17720) );
no02f80 g552664 ( .a(n_16801), .b(n_16800), .o(n_17000) );
no02f80 g552665 ( .a(n_16976), .b(n_16378), .o(n_17723) );
no02f80 g552666 ( .a(n_16998), .b(n_16377), .o(n_17724) );
na02f80 g552667 ( .a(n_16998), .b(n_16997), .o(n_16999) );
na02f80 g552668 ( .a(n_17266), .b(n_16662), .o(n_17954) );
na02f80 g552669 ( .a(n_17266), .b(n_17061), .o(n_16996) );
oa12f80 g552670 ( .a(n_16798), .b(n_327), .c(FE_OFN1119_rst), .o(n_16799) );
oa12f80 g552671 ( .a(n_16798), .b(n_796), .c(FE_OFN350_n_4860), .o(n_16797) );
na02f80 g552672 ( .a(n_16994), .b(n_16993), .o(n_16995) );
in01f80 g552673 ( .a(n_17532), .o(n_18188) );
na02f80 g552674 ( .a(n_16903), .b(n_17533), .o(n_17532) );
na02f80 g552675 ( .a(n_16841), .b(n_16795), .o(n_16796) );
oa12f80 g552676 ( .a(FE_OFN389_n_16991), .b(n_200), .c(n_28607), .o(n_16992) );
na02f80 g552677 ( .a(n_17264), .b(n_17263), .o(n_17265) );
na02f80 g552678 ( .a(n_16555), .b(n_4270), .o(n_17637) );
in01f80 g552679 ( .a(n_18491), .o(n_17531) );
oa12f80 g552680 ( .a(n_16551), .b(n_15920), .c(n_16365), .o(n_18491) );
in01f80 g552681 ( .a(n_19101), .o(n_16990) );
oa12f80 g552682 ( .a(n_16552), .b(n_15918), .c(n_15750), .o(n_19101) );
oa12f80 g552683 ( .a(n_16978), .b(n_710), .c(FE_OFN65_n_27012), .o(n_16989) );
na02f80 g552684 ( .a(n_16580), .b(n_16501), .o(n_17711) );
oa12f80 g552685 ( .a(n_17261), .b(n_799), .c(FE_OFN94_n_27449), .o(n_17262) );
oa12f80 g552686 ( .a(n_17261), .b(n_938), .c(FE_OFN72_n_27012), .o(n_17260) );
in01f80 g552687 ( .a(n_19098), .o(n_16988) );
oa12f80 g552688 ( .a(n_16546), .b(n_15913), .c(n_15748), .o(n_19098) );
oa12f80 g552689 ( .a(n_17258), .b(n_82), .c(FE_OFN99_n_27449), .o(n_17259) );
oa12f80 g552690 ( .a(n_17258), .b(n_1065), .c(FE_OFN1112_rst), .o(n_17257) );
no02f80 g552691 ( .a(n_16841), .b(n_15771), .o(n_18177) );
in01f80 g552692 ( .a(n_18237), .o(n_17530) );
oa12f80 g552693 ( .a(n_16730), .b(n_16173), .c(n_16366), .o(n_18237) );
oa12f80 g552694 ( .a(n_16971), .b(n_1900), .c(FE_OFN357_n_4860), .o(n_16987) );
in01f80 g552695 ( .a(n_19095), .o(n_16986) );
oa12f80 g552696 ( .a(n_16550), .b(n_15911), .c(n_15751), .o(n_19095) );
in01f80 g552697 ( .a(n_18487), .o(n_18101) );
oa12f80 g552698 ( .a(n_16742), .b(n_16887), .c(n_16205), .o(n_18487) );
in01f80 g552699 ( .a(n_19092), .o(n_16985) );
oa12f80 g552700 ( .a(n_16743), .b(n_16200), .c(n_15749), .o(n_19092) );
in01f80 g552701 ( .a(n_18484), .o(n_17256) );
oa12f80 g552702 ( .a(n_16741), .b(n_16064), .c(n_16198), .o(n_18484) );
oa12f80 g552703 ( .a(n_17254), .b(n_1144), .c(FE_OFN1124_rst), .o(n_17255) );
ao12f80 g552704 ( .a(n_10858), .b(n_16579), .c(n_12067), .o(n_17440) );
in01f80 g552705 ( .a(n_19089), .o(n_17253) );
oa12f80 g552706 ( .a(n_16919), .b(n_16420), .c(n_15745), .o(n_19089) );
in01f80 g552707 ( .a(n_18254), .o(n_17252) );
oa12f80 g552708 ( .a(n_16736), .b(n_16192), .c(n_16063), .o(n_18254) );
na02f80 g552709 ( .a(n_16485), .b(n_16984), .o(n_24548) );
in01f80 g552710 ( .a(n_19086), .o(n_16983) );
oa12f80 g552711 ( .a(n_16549), .b(n_15905), .c(n_15742), .o(n_19086) );
in01f80 g552712 ( .a(n_19083), .o(n_16982) );
oa12f80 g552713 ( .a(n_16288), .b(n_15612), .c(n_15741), .o(n_19083) );
na02f80 g552714 ( .a(n_17250), .b(n_17249), .o(n_17251) );
oa12f80 g552715 ( .a(n_16789), .b(n_472), .c(FE_OFN142_n_27449), .o(n_16794) );
no02f80 g552716 ( .a(n_16831), .b(n_15821), .o(n_18433) );
na02f80 g552717 ( .a(n_16831), .b(n_16792), .o(n_16793) );
no02f80 g552718 ( .a(n_16577), .b(n_16576), .o(n_16578) );
in01f80 g552719 ( .a(n_16791), .o(n_17437) );
na02f80 g552720 ( .a(n_16575), .b(n_16576), .o(n_16791) );
in01f80 g552721 ( .a(n_17946), .o(n_17529) );
na02f80 g552722 ( .a(n_16667), .b(n_17248), .o(n_17946) );
na02f80 g552723 ( .a(n_17059), .b(n_17248), .o(n_16981) );
no02f80 g552724 ( .a(n_16994), .b(n_16376), .o(n_17722) );
oa12f80 g552725 ( .a(n_16973), .b(n_72), .c(FE_OFN358_n_4860), .o(n_16980) );
in01f80 g552726 ( .a(n_17983), .o(n_17528) );
oa12f80 g552727 ( .a(n_16545), .b(n_16364), .c(n_15901), .o(n_17983) );
ao12f80 g552728 ( .a(n_16297), .b(n_16303), .c(n_13259), .o(n_16869) );
na02f80 g552729 ( .a(n_16671), .b(n_17247), .o(n_17957) );
na02f80 g552730 ( .a(n_17526), .b(n_17525), .o(n_17527) );
no02f80 g552731 ( .a(n_17245), .b(n_17244), .o(n_17246) );
no02f80 g552732 ( .a(n_17245), .b(n_16685), .o(n_17717) );
oa12f80 g552733 ( .a(FE_OFN387_n_17236), .b(n_107), .c(FE_OFN1123_rst), .o(n_17243) );
oa12f80 g552734 ( .a(n_16789), .b(n_988), .c(FE_OFN142_n_27449), .o(n_16790) );
na02f80 g552735 ( .a(n_16668), .b(n_17242), .o(n_17956) );
oa12f80 g552736 ( .a(n_16978), .b(n_1253), .c(FE_OFN124_n_27449), .o(n_16979) );
na02f80 g552737 ( .a(n_16976), .b(n_16975), .o(n_16977) );
no02f80 g552738 ( .a(n_16837), .b(n_16107), .o(n_17944) );
in01f80 g552739 ( .a(n_17979), .o(n_17241) );
oa12f80 g552740 ( .a(n_16287), .b(n_16060), .c(n_15601), .o(n_17979) );
na02f80 g552741 ( .a(n_16837), .b(n_16787), .o(n_16788) );
in01f80 g552742 ( .a(n_16574), .o(n_17430) );
oa12f80 g552743 ( .a(n_16286), .b(n_15616), .c(n_15081), .o(n_16574) );
na02f80 g552744 ( .a(n_16786), .b(n_16500), .o(n_18540) );
oa22f80 g552745 ( .a(n_15593), .b(n_12168), .c(n_14991), .d(n_12167), .o(n_17429) );
na02f80 g552746 ( .a(n_16785), .b(n_16096), .o(n_17713) );
na02f80 g552747 ( .a(n_16785), .b(n_16572), .o(n_16573) );
no02f80 g552748 ( .a(n_16783), .b(n_16782), .o(n_16784) );
in01f80 g552749 ( .a(n_18242), .o(n_17524) );
oa12f80 g552750 ( .a(n_16731), .b(n_16180), .c(n_16363), .o(n_18242) );
in01f80 g552751 ( .a(n_16781), .o(n_17432) );
na02f80 g552752 ( .a(FE_OFN1015_n_16571), .b(n_16782), .o(n_16781) );
oa12f80 g552753 ( .a(n_16973), .b(n_194), .c(FE_OFN141_n_27449), .o(n_16974) );
no02f80 g552754 ( .a(n_17239), .b(n_16648), .o(n_17727) );
oa12f80 g552755 ( .a(n_16971), .b(n_1558), .c(FE_OFN357_n_4860), .o(n_16972) );
no02f80 g552756 ( .a(n_17819), .b(n_17174), .o(n_18710) );
na02f80 g552757 ( .a(n_17819), .b(n_17522), .o(n_17523) );
na02f80 g552758 ( .a(n_17239), .b(n_17238), .o(n_17240) );
oa12f80 g552759 ( .a(n_15929), .b(n_14588), .c(n_14630), .o(n_16570) );
oa12f80 g552760 ( .a(FE_OFN387_n_17236), .b(n_1905), .c(FE_OFN1123_rst), .o(n_17237) );
in01f80 g552761 ( .a(n_18100), .o(n_18707) );
na02f80 g552762 ( .a(n_17818), .b(n_17169), .o(n_18100) );
oa12f80 g552763 ( .a(n_17518), .b(n_1520), .c(FE_OFN93_n_27449), .o(n_17521) );
na02f80 g552764 ( .a(n_17818), .b(n_17816), .o(n_17817) );
oa12f80 g552765 ( .a(n_15928), .b(n_14589), .c(n_14624), .o(n_16569) );
in01f80 g552766 ( .a(n_18465), .o(n_17520) );
oa12f80 g552767 ( .a(n_16726), .b(n_16183), .c(n_16362), .o(n_18465) );
oa12f80 g552768 ( .a(n_16779), .b(n_1155), .c(FE_OFN1120_rst), .o(n_16780) );
oa12f80 g552769 ( .a(FE_OFN46_n_17233), .b(n_631), .c(FE_OFN288_n_29266), .o(n_17234) );
oa12f80 g552770 ( .a(FE_OFN46_n_17233), .b(n_1575), .c(n_29104), .o(n_17232) );
oa12f80 g552771 ( .a(n_16798), .b(n_321), .c(FE_OFN350_n_4860), .o(n_16778) );
in01f80 g552772 ( .a(n_18268), .o(n_17231) );
oa12f80 g552773 ( .a(n_16735), .b(n_16055), .c(n_16213), .o(n_18268) );
oa12f80 g552774 ( .a(n_17518), .b(n_174), .c(FE_OFN93_n_27449), .o(n_17519) );
in01f80 g552775 ( .a(n_17517), .o(n_18178) );
na02f80 g552776 ( .a(n_16462), .b(n_17263), .o(n_17517) );
in01f80 g552777 ( .a(n_17815), .o(n_18429) );
na02f80 g552778 ( .a(n_16672), .b(n_17525), .o(n_17815) );
oa12f80 g552779 ( .a(n_16240), .b(n_14613), .c(FE_OFN25_n_11489), .o(n_16777) );
oa12f80 g552780 ( .a(n_16897), .b(n_16001), .c(n_13853), .o(n_17516) );
in01f80 g552781 ( .a(n_16568), .o(n_17426) );
oa12f80 g552782 ( .a(n_2810), .b(n_16299), .c(n_2169), .o(n_16568) );
oa12f80 g552783 ( .a(n_12466), .b(n_16302), .c(n_13656), .o(n_17119) );
in01f80 g552784 ( .a(n_16776), .o(n_17706) );
oa12f80 g552785 ( .a(n_13312), .b(n_16559), .c(n_12123), .o(n_16776) );
oa12f80 g552786 ( .a(n_16894), .b(n_16003), .c(n_11415), .o(n_17515) );
in01f80 g552787 ( .a(n_16567), .o(n_17424) );
ao12f80 g552788 ( .a(n_2156), .b(n_16295), .c(n_3160), .o(n_16567) );
oa12f80 g552789 ( .a(n_16237), .b(n_14612), .c(n_10719), .o(n_16775) );
in01f80 g552790 ( .a(n_17230), .o(n_18164) );
oa12f80 g552791 ( .a(n_16921), .b(n_16422), .c(n_13660), .o(n_17230) );
in01f80 g552792 ( .a(n_16970), .o(n_17938) );
oa12f80 g552793 ( .a(n_16729), .b(n_16178), .c(n_11114), .o(n_16970) );
in01f80 g552794 ( .a(n_16774), .o(n_17703) );
ao12f80 g552795 ( .a(n_12115), .b(n_16562), .c(n_13343), .o(n_16774) );
oa12f80 g552796 ( .a(n_15946), .b(n_14587), .c(n_14628), .o(n_16566) );
oa12f80 g552797 ( .a(n_16440), .b(n_15015), .c(n_11493), .o(n_16969) );
oa12f80 g552798 ( .a(n_17222), .b(n_1623), .c(FE_OFN116_n_27449), .o(n_17229) );
oa12f80 g552799 ( .a(n_17227), .b(n_1930), .c(FE_OFN119_n_27449), .o(n_17228) );
oa12f80 g552800 ( .a(n_17217), .b(n_331), .c(FE_OFN1120_rst), .o(n_17226) );
oa12f80 g552801 ( .a(n_17220), .b(n_390), .c(FE_OFN72_n_27012), .o(n_17225) );
oa12f80 g552802 ( .a(n_16658), .b(n_15436), .c(n_14208), .o(n_17224) );
oa12f80 g552803 ( .a(n_17222), .b(n_364), .c(FE_OFN1143_n_27012), .o(n_17223) );
oa12f80 g552804 ( .a(n_16430), .b(n_15242), .c(n_11075), .o(n_16968) );
oa12f80 g552805 ( .a(n_17220), .b(n_1920), .c(FE_OFN355_n_4860), .o(n_17221) );
oa12f80 g552806 ( .a(n_16657), .b(n_15435), .c(n_14632), .o(n_17219) );
oa12f80 g552807 ( .a(n_17217), .b(n_921), .c(FE_OFN135_n_27449), .o(n_17218) );
ao12f80 g552808 ( .a(n_4354), .b(n_14990), .c(n_5729), .o(n_15993) );
oa12f80 g552809 ( .a(n_10695), .b(n_15640), .c(n_11804), .o(n_16636) );
ao12f80 g552810 ( .a(n_9427), .b(n_16773), .c(n_9426), .o(n_17715) );
oa12f80 g552811 ( .a(n_11481), .b(n_15983), .c(n_12479), .o(n_16877) );
oa12f80 g552812 ( .a(n_11530), .b(n_16565), .c(n_12496), .o(n_17441) );
oa12f80 g552813 ( .a(n_8332), .b(n_16772), .c(n_9534), .o(n_17404) );
na03f80 g552814 ( .a(n_5355), .b(n_16719), .c(FE_OFN63_n_27012), .o(n_17631) );
na03f80 g552815 ( .a(n_5371), .b(n_16723), .c(FE_OFN74_n_27012), .o(n_17628) );
na03f80 g552816 ( .a(n_5376), .b(n_16721), .c(FE_OFN78_n_27012), .o(n_17634) );
oa12f80 g552817 ( .a(n_11809), .b(n_16301), .c(n_13110), .o(n_17118) );
in01f80 g552818 ( .a(n_18455), .o(n_17514) );
oa12f80 g552819 ( .a(n_17216), .b(n_17215), .c(n_17196), .o(n_18455) );
in01f80 g552820 ( .a(n_18754), .o(n_17513) );
oa12f80 g552821 ( .a(n_16067), .b(n_17214), .c(n_16065), .o(n_18754) );
in01f80 g552822 ( .a(n_18751), .o(n_17512) );
oa12f80 g552823 ( .a(n_16644), .b(n_17213), .c(n_16643), .o(n_18751) );
in01f80 g552824 ( .a(n_19072), .o(n_17212) );
oa12f80 g552825 ( .a(n_15744), .b(n_16967), .c(n_15743), .o(n_19072) );
in01f80 g552826 ( .a(n_19069), .o(n_17211) );
oa12f80 g552827 ( .a(n_16062), .b(n_16966), .c(n_16061), .o(n_19069) );
in01f80 g552828 ( .a(n_18200), .o(n_17511) );
oa12f80 g552829 ( .a(n_17210), .b(n_17209), .c(n_16939), .o(n_18200) );
in01f80 g552830 ( .a(n_18748), .o(n_16965) );
oa12f80 g552831 ( .a(n_16059), .b(n_16771), .c(n_16058), .o(n_18748) );
in01f80 g552832 ( .a(n_18742), .o(n_16964) );
oa12f80 g552833 ( .a(n_16069), .b(n_16770), .c(n_16068), .o(n_18742) );
in01f80 g552834 ( .a(n_18452), .o(n_17208) );
oa12f80 g552835 ( .a(n_16057), .b(n_16963), .c(n_16056), .o(n_18452) );
in01f80 g552836 ( .a(n_18745), .o(n_16962) );
oa12f80 g552837 ( .a(n_15737), .b(n_16769), .c(n_15736), .o(n_18745) );
in01f80 g552838 ( .a(n_18739), .o(n_16961) );
oa12f80 g552839 ( .a(n_15473), .b(n_16768), .c(n_15472), .o(n_18739) );
in01f80 g552840 ( .a(n_18733), .o(n_16960) );
oa12f80 g552841 ( .a(n_15469), .b(n_16767), .c(n_15468), .o(n_18733) );
in01f80 g552842 ( .a(n_18730), .o(n_16959) );
oa12f80 g552843 ( .a(n_15471), .b(n_16766), .c(n_15470), .o(n_18730) );
in01f80 g552844 ( .a(n_18727), .o(n_16958) );
oa12f80 g552845 ( .a(n_15467), .b(n_16765), .c(n_15466), .o(n_18727) );
in01f80 g552846 ( .a(n_18724), .o(n_16957) );
oa12f80 g552847 ( .a(n_15465), .b(n_16764), .c(n_15464), .o(n_18724) );
in01f80 g552848 ( .a(n_18721), .o(n_17814) );
oa12f80 g552849 ( .a(n_17510), .b(n_17509), .c(n_17508), .o(n_18721) );
in01f80 g552850 ( .a(n_18449), .o(n_16956) );
oa12f80 g552851 ( .a(n_15747), .b(n_16763), .c(n_15746), .o(n_18449) );
in01f80 g552852 ( .a(n_18191), .o(n_17207) );
oa12f80 g552853 ( .a(n_16955), .b(n_16954), .c(n_16455), .o(n_18191) );
in01f80 g552854 ( .a(n_18197), .o(n_17507) );
oa12f80 g552855 ( .a(n_17206), .b(n_17205), .c(n_16663), .o(n_18197) );
in01f80 g552856 ( .a(n_18542), .o(n_17506) );
oa12f80 g552857 ( .a(n_17204), .b(n_17203), .c(n_16453), .o(n_18542) );
in01f80 g552858 ( .a(n_19075), .o(n_17813) );
oa12f80 g552859 ( .a(n_17505), .b(n_17504), .c(n_17499), .o(n_19075) );
in01f80 g552860 ( .a(n_18718), .o(n_16953) );
oa12f80 g552861 ( .a(n_15463), .b(n_16762), .c(n_15462), .o(n_18718) );
in01f80 g552862 ( .a(n_18736), .o(n_16952) );
oa12f80 g552863 ( .a(n_15475), .b(n_16761), .c(n_15474), .o(n_18736) );
in01f80 g552864 ( .a(n_18194), .o(n_17202) );
oa12f80 g552865 ( .a(n_16951), .b(n_16950), .c(n_16441), .o(n_18194) );
in01f80 g552866 ( .a(n_18446), .o(n_16949) );
oa12f80 g552867 ( .a(n_15740), .b(n_16760), .c(n_15739), .o(n_18446) );
na03f80 g552868 ( .a(n_2624), .b(n_16281), .c(FE_OFN77_n_27012), .o(n_17099) );
ao12f80 g552869 ( .a(n_16528), .b(n_16527), .c(n_17666), .o(n_16948) );
ao22s80 g552870 ( .a(n_17214), .b(n_16026), .c(n_16642), .d(x_in_2_1), .o(n_18117) );
ao12f80 g552871 ( .a(n_16533), .b(n_16534), .c(n_16532), .o(n_16947) );
ao22s80 g552872 ( .a(FE_OFN748_n_16529), .b(n_16033), .c(x_out_49_19), .d(FE_OFN277_n_16893), .o(n_16759) );
ao22s80 g552873 ( .a(n_17213), .b(n_16351), .c(n_16641), .d(x_in_34_1), .o(n_18114) );
ao22s80 g552874 ( .a(n_16963), .b(n_16007), .c(n_16359), .d(x_in_26_1), .o(n_17878) );
ao12f80 g552875 ( .a(n_17183), .b(n_17182), .c(n_17181), .o(n_17812) );
ao22s80 g552876 ( .a(n_16967), .b(n_16354), .c(n_16357), .d(x_in_18_1), .o(n_17883) );
ao22s80 g552877 ( .a(n_16966), .b(n_16031), .c(n_16355), .d(x_in_50_1), .o(n_17875) );
ao22s80 g552878 ( .a(n_16771), .b(n_15988), .c(n_16046), .d(x_in_10_1), .o(n_17675) );
ao22s80 g552879 ( .a(n_16652), .b(n_16803), .c(n_16651), .d(n_16073), .o(n_17503) );
ao22s80 g552880 ( .a(n_16769), .b(n_15723), .c(n_16052), .d(x_in_58_1), .o(n_17667) );
ao12f80 g552881 ( .a(n_15962), .b(n_16293), .c(n_15961), .o(n_16564) );
in01f80 g552882 ( .a(n_17868), .o(n_16758) );
oa12f80 g552883 ( .a(n_15974), .b(n_16302), .c(n_15973), .o(n_17868) );
oa12f80 g552884 ( .a(n_16700), .b(n_16701), .c(n_16699), .o(n_17898) );
ao22s80 g552885 ( .a(n_16768), .b(n_15720), .c(n_16045), .d(x_in_22_1), .o(n_17664) );
ao22s80 g552886 ( .a(n_16562), .b(n_13755), .c(n_15479), .d(n_13754), .o(n_16563) );
oa12f80 g552887 ( .a(n_16276), .b(n_16275), .c(n_16277), .o(n_17414) );
ao12f80 g552888 ( .a(n_16526), .b(n_16525), .c(n_17663), .o(n_16946) );
ao22s80 g552889 ( .a(n_16761), .b(n_15724), .c(n_16047), .d(x_in_14_1), .o(n_17658) );
ao22s80 g552890 ( .a(n_16766), .b(n_15810), .c(n_16050), .d(x_in_46_1), .o(n_17655) );
ao22s80 g552891 ( .a(n_16765), .b(n_16013), .c(n_16040), .d(x_in_30_1), .o(n_17652) );
ao22s80 g552892 ( .a(n_16764), .b(n_16012), .c(n_16041), .d(x_in_62_1), .o(n_17649) );
ao12f80 g552893 ( .a(n_16715), .b(n_16714), .c(n_18116), .o(n_17201) );
in01f80 g552894 ( .a(FE_OFN450_n_17680), .o(n_17678) );
ao12f80 g552895 ( .a(n_16285), .b(n_16565), .c(n_16284), .o(n_17680) );
ao12f80 g552896 ( .a(n_16503), .b(n_16502), .c(n_17660), .o(n_16945) );
ao12f80 g552897 ( .a(n_16698), .b(n_16697), .c(n_16696), .o(n_17200) );
ao22s80 g552898 ( .a(n_16299), .b(n_3720), .c(n_15204), .d(n_3719), .o(n_16300) );
ao12f80 g552899 ( .a(n_16524), .b(n_16523), .c(n_17657), .o(n_16944) );
ao12f80 g552900 ( .a(n_16522), .b(n_16521), .c(n_17654), .o(n_16943) );
ao22s80 g552901 ( .a(n_16770), .b(n_15877), .c(n_16054), .d(x_in_42_1), .o(n_17672) );
ao12f80 g552902 ( .a(n_16713), .b(n_16712), .c(n_18113), .o(n_17199) );
ao12f80 g552903 ( .a(n_16274), .b(n_16273), .c(n_17645), .o(n_16757) );
in01f80 g552904 ( .a(n_16942), .o(n_18127) );
oa12f80 g552905 ( .a(n_16280), .b(n_16579), .c(n_16279), .o(n_16942) );
ao12f80 g552906 ( .a(n_16520), .b(n_16519), .c(n_17651), .o(n_16941) );
in01f80 g552907 ( .a(n_16862), .o(n_16561) );
oa12f80 g552908 ( .a(n_15635), .b(n_15983), .c(n_15634), .o(n_16862) );
ao12f80 g552909 ( .a(n_16518), .b(n_16517), .c(n_17648), .o(n_16940) );
ao12f80 g552910 ( .a(n_16711), .b(n_16710), .c(n_17882), .o(n_17198) );
oa12f80 g552911 ( .a(n_16531), .b(n_16530), .c(x_in_1_13), .o(n_17695) );
ao22s80 g552912 ( .a(n_16559), .b(n_13743), .c(n_15480), .d(n_13742), .o(n_16560) );
in01f80 g552913 ( .a(n_17934), .o(n_17197) );
ao12f80 g552914 ( .a(n_16484), .b(n_16939), .c(n_16675), .o(n_17934) );
ao22s80 g552915 ( .a(n_16763), .b(n_15444), .c(n_16044), .d(x_in_16_1), .o(n_17646) );
ao12f80 g552916 ( .a(n_16516), .b(n_16515), .c(n_17642), .o(n_16938) );
ao12f80 g552917 ( .a(n_16918), .b(n_16917), .c(n_16916), .o(n_17502) );
in01f80 g552918 ( .a(n_18171), .o(n_17501) );
ao12f80 g552919 ( .a(n_16692), .b(n_17196), .c(n_16899), .o(n_18171) );
in01f80 g552920 ( .a(n_15991), .o(n_16347) );
ao12f80 g552921 ( .a(n_14583), .b(n_14990), .c(n_14582), .o(n_15991) );
oa12f80 g552922 ( .a(n_14495), .b(n_16303), .c(n_16297), .o(n_16298) );
in01f80 g552923 ( .a(n_17109), .o(n_16756) );
oa12f80 g552924 ( .a(n_15972), .b(n_16303), .c(n_15971), .o(n_17109) );
ao22s80 g552925 ( .a(n_16767), .b(n_15717), .c(n_16051), .d(x_in_54_1), .o(n_17661) );
ao12f80 g552926 ( .a(n_16482), .b(n_16481), .c(n_16480), .o(n_16937) );
ao22s80 g552927 ( .a(n_16295), .b(n_3722), .c(n_15202), .d(n_3721), .o(n_16296) );
ao12f80 g552928 ( .a(n_16709), .b(n_16708), .c(n_17874), .o(n_17195) );
ao12f80 g552929 ( .a(n_16537), .b(n_16536), .c(n_16535), .o(n_16936) );
in01f80 g552930 ( .a(n_17194), .o(n_18151) );
oa12f80 g552931 ( .a(n_16539), .b(n_16773), .c(n_16538), .o(n_17194) );
ao12f80 g552932 ( .a(n_16908), .b(n_16907), .c(n_16906), .o(n_17500) );
in01f80 g552933 ( .a(n_17692), .o(n_17888) );
oa12f80 g552934 ( .a(n_16477), .b(n_16772), .c(n_16476), .o(n_17692) );
ao12f80 g552935 ( .a(n_15250), .b(n_15249), .c(n_15248), .o(n_15982) );
in01f80 g552936 ( .a(n_16343), .o(n_16630) );
ao12f80 g552937 ( .a(n_14989), .b(n_15257), .c(n_14988), .o(n_16343) );
in01f80 g552938 ( .a(n_16866), .o(n_16873) );
ao12f80 g552939 ( .a(n_15253), .b(n_15640), .c(n_15252), .o(n_16866) );
ao12f80 g552940 ( .a(n_16514), .b(n_16513), .c(n_17639), .o(n_16935) );
ao12f80 g552941 ( .a(n_16512), .b(n_16511), .c(n_16510), .o(n_16934) );
in01f80 g552942 ( .a(n_17871), .o(n_17411) );
ao12f80 g552943 ( .a(n_15970), .b(n_16301), .c(n_15969), .o(n_17871) );
ao12f80 g552944 ( .a(n_16509), .b(n_16508), .c(n_17674), .o(n_16933) );
ao12f80 g552945 ( .a(n_16507), .b(n_16506), .c(n_17671), .o(n_16932) );
in01f80 g552946 ( .a(n_18694), .o(n_18099) );
ao12f80 g552947 ( .a(n_17173), .b(n_17508), .c(n_17172), .o(n_18694) );
in01f80 g552948 ( .a(n_18421), .o(n_17811) );
ao12f80 g552949 ( .a(n_16901), .b(n_17499), .c(n_17170), .o(n_18421) );
ao12f80 g552950 ( .a(n_16505), .b(n_16504), .c(n_17877), .o(n_16931) );
ao22s80 g552951 ( .a(n_16762), .b(n_15678), .c(n_16039), .d(x_in_12_1), .o(n_17643) );
ao12f80 g552952 ( .a(n_15255), .b(n_15636), .c(n_15254), .o(n_15981) );
ao22s80 g552953 ( .a(n_16760), .b(n_15992), .c(FE_OFN834_n_16760), .d(x_in_44_1), .o(n_17640) );
oa12f80 g552954 ( .a(n_16707), .b(n_16706), .c(n_16705), .o(n_17893) );
ao12f80 g552955 ( .a(n_16703), .b(n_16704), .c(n_16702), .o(n_17193) );
oa22f80 g552956 ( .a(n_16293), .b(FE_OFN312_n_3069), .c(n_1972), .d(FE_OFN60_n_27012), .o(n_16294) );
oa22f80 g552957 ( .a(n_16929), .b(FE_OFN406_n_28303), .c(n_760), .d(FE_OFN127_n_27449), .o(n_16930) );
oa22f80 g552958 ( .a(n_16360), .b(FE_OFN236_n_4162), .c(n_140), .d(FE_OFN127_n_27449), .o(n_17192) );
ao22s80 g552959 ( .a(n_17196), .b(n_17191), .c(n_16900), .d(x_in_60_1), .o(n_17880) );
ao22s80 g552960 ( .a(n_16939), .b(n_16928), .c(n_16676), .d(x_in_6_1), .o(n_17669) );
ao22s80 g552961 ( .a(n_17499), .b(n_17498), .c(n_17171), .d(x_in_20_1), .o(n_18109) );
oa22f80 g552962 ( .a(n_15460), .b(n_29698), .c(n_653), .d(FE_OFN89_n_27449), .o(n_16558) );
oa22f80 g552963 ( .a(n_15639), .b(FE_OFN416_n_28303), .c(n_318), .d(FE_OFN108_n_27449), .o(n_16557) );
oa22f80 g552964 ( .a(n_15734), .b(FE_OFN400_n_28303), .c(n_1059), .d(n_27449), .o(n_16755) );
oa22f80 g552965 ( .a(n_16358), .b(FE_OFN292_n_3069), .c(n_821), .d(FE_OFN1115_rst), .o(n_17190) );
oa22f80 g552966 ( .a(n_16349), .b(FE_OFN294_n_3069), .c(n_592), .d(FE_OFN100_n_27449), .o(n_16927) );
oa22f80 g552967 ( .a(n_14973), .b(FE_OFN312_n_3069), .c(n_271), .d(FE_OFN18_n_29617), .o(n_15980) );
oa22f80 g552968 ( .a(n_16352), .b(FE_OFN303_n_3069), .c(n_1813), .d(FE_OFN69_n_27012), .o(n_16926) );
oa22f80 g552969 ( .a(n_17032), .b(n_29698), .c(n_706), .d(FE_OFN347_n_4860), .o(n_16925) );
oa22f80 g552970 ( .a(n_14977), .b(n_29698), .c(n_116), .d(FE_OFN56_n_27012), .o(n_15979) );
ao22s80 g552971 ( .a(n_17508), .b(n_17497), .c(n_16902), .d(x_in_36_1), .o(n_18111) );
oa22f80 g552972 ( .a(n_15456), .b(FE_OFN269_n_4280), .c(n_1162), .d(FE_OFN1113_rst), .o(n_16556) );
oa22f80 g552973 ( .a(n_16753), .b(FE_OFN240_n_4162), .c(n_1961), .d(FE_OFN352_n_4860), .o(n_16754) );
oa22f80 g552974 ( .a(n_15195), .b(FE_OFN410_n_28303), .c(n_923), .d(FE_OFN127_n_27449), .o(n_16292) );
oa22f80 g552975 ( .a(n_15636), .b(n_29496), .c(n_658), .d(FE_OFN129_n_27449), .o(n_15637) );
oa22f80 g552976 ( .a(n_14975), .b(FE_OFN295_n_3069), .c(n_1428), .d(FE_OFN127_n_27449), .o(n_15978) );
oa22f80 g552977 ( .a(n_15729), .b(FE_OFN406_n_28303), .c(n_1214), .d(FE_OFN355_n_4860), .o(n_16752) );
oa22f80 g552978 ( .a(n_15193), .b(FE_OFN264_n_4280), .c(n_1615), .d(FE_OFN329_n_4860), .o(n_16291) );
oa22f80 g552979 ( .a(n_15197), .b(FE_OFN257_n_4280), .c(n_964), .d(FE_OFN1118_rst), .o(n_16290) );
oa22f80 g552980 ( .a(FE_OFN981_n_16353), .b(FE_OFN292_n_3069), .c(n_302), .d(n_25680), .o(n_16924) );
oa22f80 g552981 ( .a(n_14972), .b(FE_OFN265_n_4280), .c(n_1804), .d(FE_OFN129_n_27449), .o(n_15977) );
oa22f80 g552982 ( .a(FE_OFN835_n_16760), .b(n_23291), .c(n_972), .d(FE_OFN89_n_27449), .o(n_16751) );
ao22s80 g552983 ( .a(n_16356), .b(n_15441), .c(x_out_47_19), .d(FE_OFN273_n_16893), .o(n_17189) );
ao12f80 g552984 ( .a(n_16282), .b(x_out_56_31), .c(FE_OFN37_n_17184), .o(n_16750) );
ao22s80 g552985 ( .a(n_16554), .b(n_2892), .c(x_out_57_31), .d(n_17184), .o(n_16749) );
ao12f80 g552986 ( .a(n_16724), .b(x_out_58_31), .c(FE_OFN37_n_17184), .o(n_17188) );
ao12f80 g552987 ( .a(n_16722), .b(x_out_59_31), .c(FE_OFN37_n_17184), .o(n_17187) );
ao12f80 g552988 ( .a(n_16720), .b(x_out_62_31), .c(n_17184), .o(n_17185) );
no02f80 g553052 ( .a(n_16554), .b(x_in_39_15), .o(n_16555) );
in01f80 g553053 ( .a(n_15975), .o(n_15976) );
no02f80 g553054 ( .a(n_16275), .b(x_in_24_4), .o(n_15975) );
na03f80 g553055 ( .a(n_15677), .b(n_18822), .c(FE_OFN422_n_16909), .o(n_16991) );
no02f80 g553056 ( .a(n_17182), .b(n_17181), .o(n_17183) );
in01f80 g553057 ( .a(n_16922), .o(n_16923) );
na02f80 g553058 ( .a(n_16748), .b(n_16211), .o(n_16922) );
na02f80 g553059 ( .a(n_16275), .b(x_in_24_4), .o(n_16592) );
na03f80 g553060 ( .a(n_15292), .b(n_18209), .c(FE_OFN384_n_16289), .o(n_16779) );
na02f80 g553061 ( .a(n_16553), .b(x_in_38_5), .o(n_17349) );
in01f80 g553062 ( .a(n_16746), .o(n_16747) );
no02f80 g553063 ( .a(n_16553), .b(x_in_38_5), .o(n_16746) );
na02f80 g553064 ( .a(n_16302), .b(n_15973), .o(n_15974) );
na02f80 g553065 ( .a(n_16921), .b(n_16423), .o(n_17588) );
in01f80 g553066 ( .a(n_17179), .o(n_17180) );
na02f80 g553067 ( .a(n_16920), .b(n_16407), .o(n_17179) );
in01f80 g553068 ( .a(n_16744), .o(n_16745) );
no02f80 g553069 ( .a(n_16544), .b(x_in_24_3), .o(n_16744) );
na02f80 g553070 ( .a(n_16552), .b(n_15919), .o(n_17021) );
na02f80 g553071 ( .a(n_16551), .b(n_15921), .o(n_17006) );
na02f80 g553072 ( .a(n_16550), .b(n_15912), .o(n_17018) );
na02f80 g553073 ( .a(n_16743), .b(n_16201), .o(n_17289) );
na02f80 g553074 ( .a(n_16742), .b(n_16206), .o(n_17286) );
na02f80 g553075 ( .a(n_16741), .b(n_16199), .o(n_17283) );
na02f80 g553076 ( .a(n_16919), .b(n_16421), .o(n_17537) );
na02f80 g553077 ( .a(n_16549), .b(n_15906), .o(n_17015) );
in01f80 g553078 ( .a(n_16739), .o(n_16740) );
na02f80 g553079 ( .a(n_16548), .b(n_15904), .o(n_16739) );
na02f80 g553080 ( .a(n_16547), .b(x_in_0_11), .o(n_17334) );
in01f80 g553081 ( .a(n_16737), .o(n_16738) );
no02f80 g553082 ( .a(n_16547), .b(x_in_0_11), .o(n_16737) );
na02f80 g553083 ( .a(n_16736), .b(n_16193), .o(n_17280) );
na02f80 g553084 ( .a(n_16735), .b(n_16214), .o(n_17277) );
no02f80 g553085 ( .a(n_16917), .b(n_16916), .o(n_16918) );
no02f80 g553086 ( .a(n_16917), .b(n_15325), .o(n_17561) );
na03f80 g553087 ( .a(n_16022), .b(n_18203), .c(n_16289), .o(n_16973) );
na02f80 g553088 ( .a(n_16288), .b(n_15613), .o(n_16811) );
na02f80 g553089 ( .a(n_16546), .b(n_15914), .o(n_17012) );
na02f80 g553090 ( .a(n_16734), .b(x_in_8_3), .o(n_17558) );
in01f80 g553091 ( .a(n_16914), .o(n_16915) );
no02f80 g553092 ( .a(n_16734), .b(x_in_8_3), .o(n_16914) );
na02f80 g553093 ( .a(n_16545), .b(n_15902), .o(n_17009) );
na03f80 g553094 ( .a(n_16034), .b(n_19414), .c(FE_OFN422_n_16909), .o(n_17236) );
na03f80 g553095 ( .a(n_15346), .b(n_18206), .c(n_16289), .o(n_16789) );
na03f80 g553096 ( .a(n_15714), .b(n_18458), .c(FE_OFN419_n_16909), .o(n_16978) );
no02f80 g553097 ( .a(n_14580), .b(n_15254), .o(n_16346) );
na02f80 g553098 ( .a(n_16544), .b(x_in_24_3), .o(n_17331) );
in01f80 g553099 ( .a(n_16542), .o(n_16543) );
no02f80 g553100 ( .a(n_17296), .b(x_in_28_5), .o(n_16542) );
na02f80 g553101 ( .a(n_16287), .b(n_15602), .o(n_16808) );
na02f80 g553102 ( .a(n_16286), .b(n_15617), .o(n_16805) );
na02f80 g553103 ( .a(n_16541), .b(x_in_56_2), .o(n_17328) );
in01f80 g553104 ( .a(n_16732), .o(n_16733) );
no02f80 g553105 ( .a(n_16541), .b(x_in_56_2), .o(n_16732) );
na02f80 g553106 ( .a(n_17296), .b(x_in_28_5), .o(n_17044) );
na02f80 g553107 ( .a(n_16731), .b(n_16181), .o(n_17274) );
in01f80 g553108 ( .a(n_17177), .o(n_17178) );
na02f80 g553109 ( .a(n_16913), .b(n_16411), .o(n_17177) );
in01f80 g553110 ( .a(n_16911), .o(n_16912) );
na02f80 g553111 ( .a(n_16072), .b(x_in_4_11), .o(n_16911) );
na02f80 g553112 ( .a(n_16071), .b(n_1168), .o(n_17299) );
na03f80 g553113 ( .a(n_16015), .b(n_19737), .c(FE_OFN419_n_16909), .o(n_16971) );
na02f80 g553114 ( .a(n_16730), .b(n_16174), .o(n_17271) );
na02f80 g553115 ( .a(n_16729), .b(n_16179), .o(n_17358) );
in01f80 g553116 ( .a(n_17175), .o(n_17176) );
na02f80 g553117 ( .a(n_16910), .b(n_16413), .o(n_17175) );
na03f80 g553118 ( .a(n_16021), .b(n_19129), .c(FE_OFN419_n_16909), .o(n_17518) );
in01f80 g553119 ( .a(n_16727), .o(n_16728) );
na02f80 g553120 ( .a(n_16540), .b(n_15895), .o(n_16727) );
na02f80 g553121 ( .a(n_16726), .b(n_16184), .o(n_17268) );
no02f80 g553122 ( .a(n_15636), .b(n_15254), .o(n_15255) );
no02f80 g553123 ( .a(n_14990), .b(n_14582), .o(n_14583) );
no02f80 g553124 ( .a(n_15893), .b(x_in_1_13), .o(n_16844) );
no02f80 g553125 ( .a(n_15640), .b(n_15252), .o(n_15253) );
na02f80 g553126 ( .a(n_16075), .b(x_in_4_14), .o(n_16725) );
na02f80 g553127 ( .a(n_16773), .b(n_16538), .o(n_16539) );
na02f80 g553128 ( .a(n_15983), .b(n_15634), .o(n_15635) );
no02f80 g553129 ( .a(n_16565), .b(n_16284), .o(n_16285) );
no02f80 g553130 ( .a(n_16536), .b(n_16535), .o(n_16537) );
no02f80 g553131 ( .a(n_16536), .b(n_15063), .o(n_17038) );
na02f80 g553132 ( .a(n_15281), .b(n_15967), .o(n_16283) );
no02f80 g553133 ( .a(n_16281), .b(n_7261), .o(n_16282) );
no02f80 g553134 ( .a(n_16723), .b(n_8204), .o(n_16724) );
no02f80 g553135 ( .a(n_16721), .b(n_7361), .o(n_16722) );
na02f80 g553136 ( .a(n_16579), .b(n_16279), .o(n_16280) );
no02f80 g553137 ( .a(n_16719), .b(n_7575), .o(n_16720) );
oa12f80 g553138 ( .a(n_15289), .b(n_14998), .c(n_4280), .o(n_16278) );
no02f80 g553139 ( .a(n_15257), .b(n_14988), .o(n_14989) );
na02f80 g553140 ( .a(n_16534), .b(n_15940), .o(n_17033) );
no02f80 g553141 ( .a(n_16534), .b(n_16532), .o(n_16533) );
na02f80 g553142 ( .a(n_16530), .b(x_in_1_13), .o(n_16531) );
na02f80 g553143 ( .a(n_15192), .b(n_16277), .o(n_16865) );
na02f80 g553144 ( .a(n_16275), .b(n_16277), .o(n_16276) );
na02f80 g553145 ( .a(n_16070), .b(FE_OFN1124_rst), .o(n_17254) );
na02f80 g553146 ( .a(FE_OFN748_n_16529), .b(n_15707), .o(n_17542) );
oa12f80 g553147 ( .a(n_16029), .b(n_15650), .c(FE_OFN186_n_29496), .o(n_16718) );
oa12f80 g553148 ( .a(n_16030), .b(n_15646), .c(FE_OFN293_n_3069), .o(n_16717) );
oa12f80 g553149 ( .a(n_16027), .b(n_15644), .c(FE_OFN406_n_28303), .o(n_16716) );
no02f80 g553150 ( .a(n_16527), .b(n_17666), .o(n_16528) );
no02f80 g553151 ( .a(n_16525), .b(n_17663), .o(n_16526) );
no02f80 g553152 ( .a(n_16714), .b(n_18116), .o(n_16715) );
no02f80 g553153 ( .a(n_16523), .b(n_17657), .o(n_16524) );
no02f80 g553154 ( .a(n_16521), .b(n_17654), .o(n_16522) );
no02f80 g553155 ( .a(n_16712), .b(n_18113), .o(n_16713) );
no02f80 g553156 ( .a(n_16273), .b(n_17645), .o(n_16274) );
no02f80 g553157 ( .a(n_16519), .b(n_17651), .o(n_16520) );
no02f80 g553158 ( .a(n_16517), .b(n_17648), .o(n_16518) );
no02f80 g553159 ( .a(n_16710), .b(n_17882), .o(n_16711) );
no02f80 g553160 ( .a(n_16515), .b(n_17642), .o(n_16516) );
no02f80 g553161 ( .a(n_16708), .b(n_17874), .o(n_16709) );
no02f80 g553162 ( .a(n_16513), .b(n_17639), .o(n_16514) );
no02f80 g553163 ( .a(n_16511), .b(n_16510), .o(n_16512) );
no02f80 g553164 ( .a(n_16508), .b(n_17674), .o(n_16509) );
no02f80 g553165 ( .a(n_16506), .b(n_17671), .o(n_16507) );
no02f80 g553166 ( .a(n_16504), .b(n_17877), .o(n_16505) );
no02f80 g553167 ( .a(n_16502), .b(n_17660), .o(n_16503) );
na02f80 g553168 ( .a(n_16271), .b(n_16270), .o(n_16272) );
na02f80 g553169 ( .a(n_16706), .b(n_16705), .o(n_16707) );
no02f80 g553170 ( .a(n_16706), .b(n_16182), .o(n_17298) );
na02f80 g553171 ( .a(n_16704), .b(n_16219), .o(n_17295) );
no02f80 g553172 ( .a(n_16704), .b(n_16702), .o(n_16703) );
na02f80 g553173 ( .a(n_16303), .b(n_15971), .o(n_15972) );
no02f80 g553174 ( .a(n_16301), .b(n_15969), .o(n_15970) );
na02f80 g553175 ( .a(n_16701), .b(n_15686), .o(n_17293) );
na02f80 g553176 ( .a(n_16701), .b(n_16699), .o(n_16700) );
no02f80 g553177 ( .a(n_16697), .b(n_16696), .o(n_16698) );
no02f80 g553178 ( .a(n_16907), .b(n_16906), .o(n_16908) );
in01f80 g553179 ( .a(n_16695), .o(n_17217) );
no02f80 g553180 ( .a(n_16501), .b(n_2022), .o(n_16695) );
na02f80 g553181 ( .a(n_16687), .b(rst), .o(n_17227) );
in01f80 g553182 ( .a(n_17222), .o(n_16905) );
na02f80 g553183 ( .a(n_16800), .b(FE_OFN1114_rst), .o(n_17222) );
in01f80 g553184 ( .a(n_16694), .o(n_17220) );
no02f80 g553185 ( .a(n_16500), .b(n_2022), .o(n_16694) );
na02f80 g553186 ( .a(n_15574), .b(n_16269), .o(n_16839) );
na02f80 g553187 ( .a(n_15812), .b(n_16498), .o(n_24559) );
no02f80 g553188 ( .a(n_16129), .b(n_16693), .o(n_24455) );
no02f80 g553189 ( .a(n_17196), .b(n_16899), .o(n_16692) );
na02f80 g553190 ( .a(n_16092), .b(n_16691), .o(n_17326) );
no02f80 g553191 ( .a(n_16497), .b(n_16496), .o(n_26103) );
no02f80 g553192 ( .a(n_16268), .b(n_15561), .o(n_20470) );
no02f80 g553193 ( .a(n_16385), .b(n_16904), .o(n_22247) );
no02f80 g553194 ( .a(n_16267), .b(n_15565), .o(n_22584) );
na02f80 g553195 ( .a(n_15856), .b(n_16495), .o(n_21167) );
no02f80 g553196 ( .a(n_15842), .b(n_16494), .o(n_18366) );
no02f80 g553197 ( .a(n_16125), .b(n_16690), .o(n_20082) );
no02f80 g553198 ( .a(n_16109), .b(n_16689), .o(n_24176) );
no02f80 g553199 ( .a(n_16086), .b(n_16688), .o(n_20412) );
no02f80 g553200 ( .a(n_15833), .b(n_16493), .o(n_25905) );
oa12f80 g553201 ( .a(n_15967), .b(n_397), .c(FE_OFN326_n_4860), .o(n_15968) );
oa12f80 g553202 ( .a(n_15967), .b(n_339), .c(FE_OFN91_n_27449), .o(n_15966) );
oa12f80 g553203 ( .a(n_15967), .b(n_1965), .c(FE_OFN91_n_27449), .o(n_15965) );
na02f80 g553204 ( .a(n_15858), .b(n_16492), .o(n_21500) );
na02f80 g553205 ( .a(n_15562), .b(n_16266), .o(n_21569) );
no02f80 g553206 ( .a(n_15760), .b(n_16491), .o(n_18616) );
no02f80 g553207 ( .a(n_15550), .b(n_16265), .o(n_16884) );
na02f80 g553208 ( .a(n_15566), .b(n_16264), .o(n_17467) );
na02f80 g553209 ( .a(n_15558), .b(n_16263), .o(n_19394) );
no02f80 g553210 ( .a(n_15764), .b(n_16490), .o(n_24544) );
in01f80 g553211 ( .a(n_16489), .o(n_17400) );
oa12f80 g553212 ( .a(n_16215), .b(n_15656), .c(n_14619), .o(n_16489) );
na02f80 g553213 ( .a(n_15568), .b(n_16262), .o(n_19364) );
na02f80 g553214 ( .a(n_15781), .b(n_16488), .o(n_24754) );
in01f80 g553215 ( .a(n_16903), .o(n_17534) );
no02f80 g553216 ( .a(n_16687), .b(n_16686), .o(n_16903) );
no02f80 g553217 ( .a(n_15830), .b(n_16487), .o(n_24879) );
no02f80 g553218 ( .a(n_15556), .b(n_16261), .o(n_18681) );
in01f80 g553219 ( .a(n_16485), .o(n_16486) );
na02f80 g553220 ( .a(n_15731), .b(n_13831), .o(n_16485) );
na02f80 g553221 ( .a(n_15732), .b(n_13832), .o(n_16984) );
no02f80 g553222 ( .a(n_16939), .b(n_16675), .o(n_16484) );
no02f80 g553223 ( .a(n_15805), .b(n_16483), .o(n_24534) );
na02f80 g553224 ( .a(n_15482), .b(n_16260), .o(n_23577) );
no02f80 g553225 ( .a(n_16481), .b(n_16480), .o(n_16482) );
in01f80 g553226 ( .a(n_16685), .o(n_17244) );
na02f80 g553227 ( .a(n_16481), .b(FE_OFN897_n_15930), .o(n_16685) );
in01f80 g553228 ( .a(n_18124), .o(n_16684) );
oa12f80 g553229 ( .a(n_16414), .b(n_15680), .c(n_14199), .o(n_18124) );
in01f80 g553230 ( .a(n_17522), .o(n_17174) );
no02f80 g553231 ( .a(n_16902), .b(n_17172), .o(n_17522) );
na02f80 g553232 ( .a(n_16479), .b(n_15802), .o(n_22897) );
oa12f80 g553233 ( .a(n_15967), .b(n_421), .c(FE_OFN91_n_27449), .o(n_15964) );
no02f80 g553234 ( .a(n_16478), .b(n_15795), .o(n_23758) );
na02f80 g553235 ( .a(n_16772), .b(n_16476), .o(n_16477) );
no02f80 g553236 ( .a(n_17499), .b(n_17170), .o(n_16901) );
no02f80 g553237 ( .a(n_15525), .b(n_16259), .o(n_21946) );
na02f80 g553238 ( .a(n_15799), .b(n_16475), .o(n_20842) );
na02f80 g553239 ( .a(n_15521), .b(n_16258), .o(n_19029) );
no02f80 g553240 ( .a(n_15519), .b(n_16257), .o(n_18057) );
na02f80 g553241 ( .a(n_15517), .b(n_16256), .o(n_17128) );
no02f80 g553242 ( .a(n_15797), .b(n_16474), .o(n_17024) );
no02f80 g553243 ( .a(n_15523), .b(n_16255), .o(n_19688) );
no02f80 g553244 ( .a(n_15511), .b(n_16254), .o(n_23853) );
no02f80 g553245 ( .a(n_15249), .b(n_15248), .o(n_15250) );
no02f80 g553246 ( .a(n_15249), .b(n_14572), .o(n_16629) );
no02f80 g553247 ( .a(n_16683), .b(n_16094), .o(n_17973) );
in01f80 g553248 ( .a(n_15963), .o(n_16849) );
ao12f80 g553249 ( .a(n_10966), .b(n_15633), .c(n_12094), .o(n_15963) );
no02f80 g553250 ( .a(n_16293), .b(n_15961), .o(n_15962) );
na02f80 g553251 ( .a(n_15783), .b(n_16473), .o(n_24542) );
na02f80 g553252 ( .a(n_15792), .b(n_16472), .o(n_22791) );
no02f80 g553253 ( .a(n_16103), .b(n_16682), .o(n_21856) );
na02f80 g553254 ( .a(n_16101), .b(n_16681), .o(n_20742) );
no02f80 g553255 ( .a(n_16099), .b(n_16680), .o(n_19946) );
na02f80 g553256 ( .a(n_16097), .b(n_16679), .o(n_18927) );
na02f80 g553257 ( .a(n_16678), .b(n_16127), .o(n_23216) );
no02f80 g553258 ( .a(n_16253), .b(n_15510), .o(n_17975) );
na02f80 g553259 ( .a(n_15779), .b(n_16471), .o(n_22786) );
na02f80 g553260 ( .a(n_15776), .b(n_16470), .o(n_24540) );
no02f80 g553261 ( .a(n_15504), .b(n_16252), .o(n_21852) );
na02f80 g553262 ( .a(n_15502), .b(n_16251), .o(n_20738) );
no02f80 g553263 ( .a(n_15532), .b(n_16250), .o(n_19942) );
no02f80 g553264 ( .a(n_17508), .b(n_17172), .o(n_17173) );
no02f80 g553265 ( .a(n_16249), .b(n_15497), .o(n_23749) );
na02f80 g553266 ( .a(n_15494), .b(n_16248), .o(n_24750) );
no02f80 g553267 ( .a(n_17171), .b(n_17170), .o(n_17818) );
na02f80 g553268 ( .a(n_16677), .b(n_16091), .o(n_23501) );
no02f80 g553269 ( .a(n_16676), .b(n_16675), .o(n_17263) );
na02f80 g553270 ( .a(n_15767), .b(n_16469), .o(n_24536) );
na02f80 g553271 ( .a(n_15500), .b(n_16247), .o(n_18923) );
in01f80 g553272 ( .a(n_16246), .o(n_16860) );
na02f80 g553273 ( .a(n_16293), .b(n_14916), .o(n_16246) );
no02f80 g553274 ( .a(n_16088), .b(n_16674), .o(n_22521) );
na02f80 g553275 ( .a(n_16080), .b(n_16673), .o(n_19609) );
no02f80 g553276 ( .a(n_16900), .b(n_16899), .o(n_17525) );
na02f80 g553277 ( .a(n_16245), .b(n_15483), .o(n_17734) );
na02f80 g553278 ( .a(n_15552), .b(n_16244), .o(n_17807) );
in01f80 g553279 ( .a(n_16898), .o(n_17860) );
oa12f80 g553280 ( .a(n_16653), .b(n_16024), .c(n_15427), .o(n_16898) );
oa12f80 g553281 ( .a(n_15950), .b(n_15960), .c(n_13915), .o(n_16847) );
oa12f80 g553282 ( .a(n_14962), .b(n_15959), .c(n_14006), .o(n_16859) );
oa12f80 g553283 ( .a(n_13658), .b(n_15606), .c(n_14795), .o(n_16838) );
ao12f80 g553284 ( .a(n_15343), .b(n_16169), .c(n_14759), .o(n_16628) );
ao12f80 g553285 ( .a(n_15403), .b(n_16208), .c(n_14667), .o(n_16627) );
ao12f80 g553286 ( .a(n_15393), .b(n_16203), .c(n_14732), .o(n_16626) );
ao12f80 g553287 ( .a(n_14372), .b(n_15909), .c(n_15138), .o(n_16625) );
ao12f80 g553288 ( .a(n_15381), .b(n_16196), .c(n_14700), .o(n_16624) );
oa12f80 g553289 ( .a(n_15655), .b(n_15958), .c(n_14838), .o(n_16856) );
ao12f80 g553290 ( .a(n_15363), .b(n_16190), .c(n_14678), .o(n_16623) );
ao12f80 g553291 ( .a(n_11475), .b(n_15957), .c(n_12460), .o(n_16853) );
ao12f80 g553292 ( .a(n_13628), .b(n_15956), .c(n_14662), .o(n_16857) );
in01f80 g553293 ( .a(n_15955), .o(n_16851) );
ao12f80 g553294 ( .a(n_12296), .b(n_15628), .c(n_12955), .o(n_15955) );
ao12f80 g553295 ( .a(n_15413), .b(n_16186), .c(n_14774), .o(n_16858) );
oa12f80 g553296 ( .a(n_11454), .b(n_15246), .c(n_12446), .o(n_16342) );
ao12f80 g553297 ( .a(n_16243), .b(n_16445), .c(n_15021), .o(n_17369) );
oa12f80 g553298 ( .a(n_14644), .b(n_16468), .c(n_15374), .o(n_17399) );
ao12f80 g553299 ( .a(n_12257), .b(n_15632), .c(n_12934), .o(n_16622) );
oa22f80 g553300 ( .a(n_15674), .b(FE_OFN400_n_28303), .c(n_926), .d(FE_OFN347_n_4860), .o(n_16467) );
oa12f80 g553301 ( .a(n_16234), .b(n_16242), .c(n_13856), .o(n_17074) );
na03f80 g553302 ( .a(n_2536), .b(n_15293), .c(FE_OFN1119_rst), .o(n_16798) );
oa12f80 g553303 ( .a(n_8825), .b(n_15954), .c(n_10343), .o(n_16855) );
oa12f80 g553304 ( .a(n_11198), .b(n_15631), .c(n_12819), .o(n_16618) );
ao12f80 g553305 ( .a(n_12071), .b(n_15953), .c(n_13235), .o(n_16854) );
ao12f80 g553306 ( .a(n_13644), .b(n_16466), .c(n_14728), .o(n_17394) );
oa12f80 g553307 ( .a(n_14312), .b(n_15882), .c(n_15169), .o(n_16617) );
oa12f80 g553308 ( .a(n_14407), .b(n_15952), .c(n_15151), .o(n_16852) );
oa12f80 g553309 ( .a(n_10727), .b(n_15245), .c(n_11794), .o(n_16341) );
na03f80 g553310 ( .a(n_16270), .b(n_16271), .c(n_12894), .o(n_16465) );
ao12f80 g553311 ( .a(n_13655), .b(n_15582), .c(n_14653), .o(n_17025) );
ao12f80 g553312 ( .a(n_14229), .b(n_15866), .c(n_15117), .o(n_16614) );
ao12f80 g553313 ( .a(n_10675), .b(n_15630), .c(n_11802), .o(n_16612) );
oa12f80 g553314 ( .a(n_8833), .b(n_15629), .c(n_9535), .o(n_16611) );
na03f80 g553315 ( .a(n_5368), .b(n_16397), .c(FE_OFN64_n_27012), .o(n_17233) );
na03f80 g553316 ( .a(n_5042), .b(n_16399), .c(FE_OFN68_n_27012), .o(n_17258) );
na03f80 g553317 ( .a(n_5363), .b(n_16401), .c(FE_OFN64_n_27012), .o(n_17261) );
in01f80 g553318 ( .a(n_17526), .o(n_16672) );
oa12f80 g553319 ( .a(n_15892), .b(n_16242), .c(n_15891), .o(n_17526) );
oa12f80 g553320 ( .a(n_16085), .b(n_16084), .c(n_16387), .o(n_17319) );
ao22s80 g553321 ( .a(n_15439), .b(n_15184), .c(x_out_48_19), .d(n_16028), .o(n_16240) );
ao12f80 g553322 ( .a(n_15876), .b(n_15875), .c(n_16035), .o(n_16464) );
ao12f80 g553323 ( .a(n_15786), .b(n_15827), .c(n_15935), .o(n_16463) );
oa12f80 g553324 ( .a(n_16383), .b(n_16384), .c(n_16382), .o(n_17595) );
oa12f80 g553325 ( .a(n_16146), .b(n_16147), .c(n_16145), .o(n_17325) );
ao12f80 g553326 ( .a(n_16429), .b(x_out_50_19), .c(n_16028), .o(n_16897) );
ao12f80 g553327 ( .a(n_16427), .b(n_16426), .c(n_16425), .o(n_16896) );
oa12f80 g553328 ( .a(n_16380), .b(n_16379), .c(n_16381), .o(n_17594) );
ao12f80 g553329 ( .a(n_14965), .b(n_15960), .c(n_15950), .o(n_15951) );
ao12f80 g553330 ( .a(n_15220), .b(n_15949), .c(n_15948), .o(n_16604) );
in01f80 g553331 ( .a(n_17264), .o(n_16462) );
oa12f80 g553332 ( .a(n_15619), .b(n_15960), .c(n_15618), .o(n_17264) );
oa12f80 g553333 ( .a(n_16113), .b(n_16124), .c(n_16112), .o(n_17353) );
ao12f80 g553334 ( .a(n_15615), .b(n_15959), .c(n_15614), .o(n_17533) );
ao22s80 g553335 ( .a(n_15294), .b(n_2773), .c(x_out_54_30), .d(FE_OFN37_n_17184), .o(n_16461) );
ao22s80 g553336 ( .a(n_15591), .b(n_4308), .c(x_out_56_30), .d(FE_OFN280_n_16656), .o(n_15947) );
ao12f80 g553337 ( .a(n_15926), .b(x_out_57_30), .c(n_5003), .o(n_16460) );
oa12f80 g553338 ( .a(n_16153), .b(n_16152), .c(n_16151), .o(n_17348) );
ao22s80 g553339 ( .a(n_16159), .b(n_4320), .c(x_out_58_30), .d(FE_OFN276_n_16893), .o(n_16459) );
oa12f80 g553340 ( .a(n_16136), .b(n_16140), .c(n_16135), .o(n_17347) );
in01f80 g553341 ( .a(n_17062), .o(n_16671) );
oa12f80 g553342 ( .a(n_15883), .b(n_15882), .c(n_15881), .o(n_17062) );
oa12f80 g553343 ( .a(n_16144), .b(n_16393), .c(n_16194), .o(n_17343) );
ao12f80 g553344 ( .a(n_16163), .b(n_16162), .c(x_in_47_14), .o(n_16670) );
ao22s80 g553345 ( .a(n_16155), .b(n_4888), .c(x_out_62_30), .d(FE_OFN279_n_16656), .o(n_16458) );
oa12f80 g553346 ( .a(n_16142), .b(n_16143), .c(n_16141), .o(n_17342) );
ao12f80 g553347 ( .a(n_16165), .b(n_16164), .c(x_in_63_14), .o(n_16669) );
in01f80 g553348 ( .a(n_17306), .o(n_17580) );
ao12f80 g553349 ( .a(n_16187), .b(n_16186), .c(n_16185), .o(n_17306) );
ao12f80 g553350 ( .a(n_15576), .b(n_15575), .c(n_15754), .o(n_16239) );
in01f80 g553351 ( .a(n_16580), .o(n_16238) );
ao12f80 g553352 ( .a(n_15234), .b(n_15631), .c(n_15233), .o(n_16580) );
oa12f80 g553353 ( .a(n_16115), .b(n_16116), .c(n_16114), .o(n_17341) );
in01f80 g553354 ( .a(n_17304), .o(n_17569) );
ao12f80 g553355 ( .a(n_16209), .b(n_16208), .c(n_16207), .o(n_17304) );
in01f80 g553356 ( .a(n_17060), .o(n_16668) );
oa12f80 g553357 ( .a(n_15880), .b(n_15952), .c(n_15879), .o(n_17060) );
in01f80 g553358 ( .a(n_17312), .o(n_17568) );
ao12f80 g553359 ( .a(n_16204), .b(n_16203), .c(n_16202), .o(n_17312) );
in01f80 g553360 ( .a(n_17059), .o(n_16667) );
oa12f80 g553361 ( .a(n_15910), .b(n_15909), .c(n_15908), .o(n_17059) );
in01f80 g553362 ( .a(n_16895), .o(n_17845) );
oa12f80 g553363 ( .a(n_16161), .b(n_16466), .c(n_16160), .o(n_16895) );
in01f80 g553364 ( .a(n_17310), .o(n_17567) );
ao12f80 g553365 ( .a(n_16197), .b(n_16196), .c(n_16195), .o(n_17310) );
oa12f80 g553366 ( .a(n_15597), .b(n_15625), .c(n_15596), .o(n_17250) );
ao12f80 g553367 ( .a(n_15540), .b(n_15539), .c(n_15538), .o(n_25633) );
in01f80 g553368 ( .a(n_17029), .o(n_16606) );
ao22s80 g553369 ( .a(n_14573), .b(n_13509), .c(n_15628), .d(n_13508), .o(n_17029) );
in01f80 g553370 ( .a(n_17308), .o(n_17566) );
ao12f80 g553371 ( .a(n_16191), .b(n_16190), .c(n_16189), .o(n_17308) );
in01f80 g553372 ( .a(n_17300), .o(n_17565) );
ao22s80 g553373 ( .a(n_15995), .b(n_14901), .c(n_15994), .d(n_15958), .o(n_17300) );
in01f80 g553374 ( .a(n_16457), .o(n_17374) );
oa12f80 g553375 ( .a(n_15610), .b(n_15957), .c(n_15609), .o(n_16457) );
oa12f80 g553376 ( .a(n_15621), .b(n_15620), .c(x_in_1_12), .o(n_16836) );
ao12f80 g553377 ( .a(n_15917), .b(n_15916), .c(n_15915), .o(n_16456) );
in01f80 g553378 ( .a(n_17393), .o(n_16666) );
ao12f80 g553379 ( .a(n_15820), .b(n_16455), .c(n_15819), .o(n_17393) );
ao12f80 g553380 ( .a(n_15816), .b(n_15815), .c(n_16222), .o(n_16454) );
oa12f80 g553381 ( .a(n_15814), .b(n_15813), .c(n_15907), .o(n_17054) );
ao12f80 g553382 ( .a(n_16428), .b(x_out_34_19), .c(FE_OFN277_n_16893), .o(n_16894) );
ao12f80 g553383 ( .a(n_16417), .b(n_16416), .c(n_16415), .o(n_16892) );
oa12f80 g553384 ( .a(n_15227), .b(n_15622), .c(n_15226), .o(n_17239) );
ao12f80 g553385 ( .a(n_16167), .b(n_16166), .c(x_in_15_14), .o(n_16665) );
in01f80 g553386 ( .a(n_17392), .o(n_16664) );
ao12f80 g553387 ( .a(n_15808), .b(n_16453), .c(n_15807), .o(n_17392) );
ao22s80 g553388 ( .a(n_15437), .b(n_15007), .c(x_out_35_19), .d(FE_OFN280_n_16656), .o(n_16237) );
ao12f80 g553389 ( .a(n_15925), .b(n_15924), .c(FE_OFN895_n_15923), .o(n_16452) );
in01f80 g553390 ( .a(n_17245), .o(n_16236) );
oa12f80 g553391 ( .a(n_15232), .b(n_15629), .c(n_15231), .o(n_17245) );
oa12f80 g553392 ( .a(n_16123), .b(n_16374), .c(n_16122), .o(n_17356) );
in01f80 g553393 ( .a(n_16801), .o(n_16451) );
oa12f80 g553394 ( .a(n_15604), .b(n_15956), .c(n_15603), .o(n_16801) );
oa12f80 g553395 ( .a(n_16396), .b(n_16395), .c(n_16394), .o(n_17559) );
ao12f80 g553396 ( .a(n_14920), .b(n_16242), .c(n_16234), .o(n_16235) );
ao12f80 g553397 ( .a(n_15887), .b(n_15886), .c(n_15885), .o(n_16450) );
in01f80 g553398 ( .a(n_16607), .o(n_16595) );
ao12f80 g553399 ( .a(n_14983), .b(n_14982), .c(n_14981), .o(n_16607) );
oa12f80 g553400 ( .a(n_15578), .b(n_15953), .c(n_15577), .o(n_16837) );
in01f80 g553401 ( .a(n_17618), .o(n_16891) );
ao12f80 g553402 ( .a(n_16106), .b(n_16663), .c(n_16105), .o(n_17618) );
oa12f80 g553403 ( .a(n_15583), .b(n_15582), .c(n_15581), .o(n_16831) );
oa12f80 g553404 ( .a(n_16119), .b(n_16120), .c(n_16118), .o(n_17352) );
oa12f80 g553405 ( .a(n_15863), .b(n_15862), .c(n_16131), .o(n_17063) );
ao22s80 g553406 ( .a(n_16157), .b(n_2987), .c(x_out_59_30), .d(n_16893), .o(n_16449) );
in01f80 g553407 ( .a(n_16575), .o(n_16577) );
ao12f80 g553408 ( .a(n_14987), .b(n_15246), .c(n_14986), .o(n_16575) );
oa12f80 g553409 ( .a(n_15846), .b(n_15845), .c(n_16117), .o(n_17066) );
in01f80 g553410 ( .a(n_16786), .o(n_16448) );
ao12f80 g553411 ( .a(n_15589), .b(n_15592), .c(n_15588), .o(n_16786) );
ao12f80 g553412 ( .a(n_15870), .b(n_15869), .c(n_15868), .o(n_16447) );
in01f80 g553413 ( .a(n_16785), .o(n_16830) );
ao12f80 g553414 ( .a(n_15240), .b(n_15633), .c(n_15239), .o(n_16785) );
oa12f80 g553415 ( .a(n_15788), .b(n_15789), .c(n_15787), .o(n_17051) );
in01f80 g553416 ( .a(FE_OFN1015_n_16571), .o(n_16783) );
ao12f80 g553417 ( .a(n_15225), .b(n_15630), .c(n_15224), .o(n_16571) );
oa12f80 g553418 ( .a(n_15587), .b(n_15624), .c(n_15586), .o(n_16976) );
oa12f80 g553419 ( .a(n_15692), .b(n_16445), .c(n_16243), .o(n_16446) );
oa12f80 g553420 ( .a(n_15506), .b(n_16233), .c(n_16232), .o(n_16828) );
in01f80 g553421 ( .a(n_17816), .o(n_17169) );
oa12f80 g553422 ( .a(n_16409), .b(n_16445), .c(n_16408), .o(n_17816) );
oa22f80 g553423 ( .a(n_23062), .b(n_2608), .c(n_16444), .d(x_in_4_15), .o(n_25711) );
ao22s80 g553424 ( .a(n_14995), .b(n_14081), .c(x_out_40_19), .d(FE_OFN271_n_16028), .o(n_15946) );
ao12f80 g553425 ( .a(n_15580), .b(n_15937), .c(n_15579), .o(n_16231) );
in01f80 g553426 ( .a(n_16306), .o(n_16582) );
ao12f80 g553427 ( .a(n_14985), .b(n_15245), .c(n_14984), .o(n_16306) );
oa12f80 g553428 ( .a(n_15585), .b(n_15623), .c(n_15584), .o(n_16998) );
in01f80 g553429 ( .a(n_16443), .o(n_17366) );
oa12f80 g553430 ( .a(n_15595), .b(n_15954), .c(n_15594), .o(n_16443) );
oa12f80 g553431 ( .a(n_16172), .b(n_16468), .c(n_16171), .o(n_17819) );
ao12f80 g553432 ( .a(n_15492), .b(n_15491), .c(n_15490), .o(n_25459) );
ao12f80 g553433 ( .a(n_15898), .b(n_15897), .c(n_15896), .o(n_16442) );
in01f80 g553434 ( .a(n_16230), .o(n_17080) );
oa12f80 g553435 ( .a(n_15238), .b(n_15632), .c(n_15237), .o(n_16230) );
in01f80 g553436 ( .a(n_17302), .o(n_17555) );
ao12f80 g553437 ( .a(n_16170), .b(n_16169), .c(n_16168), .o(n_17302) );
in01f80 g553438 ( .a(n_17061), .o(n_16662) );
oa12f80 g553439 ( .a(n_15867), .b(n_15866), .c(n_15865), .o(n_17061) );
in01f80 g553440 ( .a(n_17391), .o(n_16661) );
ao12f80 g553441 ( .a(n_15770), .b(n_16441), .c(n_15769), .o(n_17391) );
oa12f80 g553442 ( .a(n_16139), .b(n_16138), .c(n_16137), .o(n_17322) );
oa12f80 g553443 ( .a(n_15608), .b(n_15607), .c(n_15606), .o(n_16841) );
in01f80 g553444 ( .a(n_17043), .o(n_16660) );
oa12f80 g553445 ( .a(n_15872), .b(n_15874), .c(n_15871), .o(n_17043) );
oa12f80 g553446 ( .a(n_15864), .b(n_15900), .c(n_16132), .o(n_17042) );
in01f80 g553447 ( .a(n_16229), .o(n_17075) );
oa12f80 g553448 ( .a(n_15236), .b(n_15627), .c(n_15235), .o(n_16229) );
ao22s80 g553449 ( .a(n_15701), .b(n_15638), .c(x_out_46_19), .d(n_16028), .o(n_16440) );
ao12f80 g553450 ( .a(n_16218), .b(n_16217), .c(FE_OFN690_n_16216), .o(n_16659) );
oa12f80 g553451 ( .a(n_15599), .b(n_15626), .c(n_15598), .o(n_16994) );
oa12f80 g553452 ( .a(n_16149), .b(n_16150), .c(n_16148), .o(n_17344) );
ao12f80 g553453 ( .a(n_15208), .b(n_15945), .c(n_15944), .o(n_16819) );
oa22f80 g553454 ( .a(n_16535), .b(FE_OFN234_n_4162), .c(n_236), .d(FE_OFN360_n_4860), .o(n_16228) );
oa22f80 g553455 ( .a(n_14885), .b(FE_OFN404_n_28303), .c(n_1450), .d(FE_OFN133_n_27449), .o(n_15943) );
oa22f80 g553456 ( .a(n_14887), .b(n_28608), .c(n_1601), .d(FE_OFN336_n_4860), .o(n_15942) );
oa22f80 g553457 ( .a(n_15331), .b(FE_OFN299_n_3069), .c(n_1355), .d(FE_OFN363_n_4860), .o(n_16439) );
ao22s80 g553458 ( .a(n_16663), .b(n_16438), .c(n_15798), .d(x_in_40_1), .o(n_17027) );
oa22f80 g553459 ( .a(n_15323), .b(FE_OFN307_n_3069), .c(n_1187), .d(FE_OFN76_n_27012), .o(n_16437) );
oa22f80 g553460 ( .a(n_15330), .b(FE_OFN306_n_3069), .c(n_1565), .d(rst), .o(n_16436) );
oa22f80 g553461 ( .a(n_15305), .b(FE_OFN303_n_3069), .c(n_173), .d(FE_OFN122_n_27449), .o(n_16435) );
oa22f80 g553462 ( .a(n_15940), .b(FE_OFN309_n_3069), .c(n_64), .d(FE_OFN122_n_27449), .o(n_15941) );
oa22f80 g553463 ( .a(n_15328), .b(FE_OFN293_n_3069), .c(n_1384), .d(FE_OFN17_n_29617), .o(n_16434) );
oa22f80 g553464 ( .a(n_14886), .b(n_23813), .c(n_829), .d(FE_OFN89_n_27449), .o(n_15939) );
oa22f80 g553465 ( .a(n_15937), .b(FE_OFN405_n_28303), .c(n_992), .d(FE_OFN1110_rst), .o(n_15938) );
ao22s80 g553466 ( .a(n_16441), .b(n_16227), .c(n_15489), .d(x_in_52_1), .o(n_16815) );
oa22f80 g553467 ( .a(n_15935), .b(FE_OFN221_n_23315), .c(n_550), .d(FE_OFN116_n_27449), .o(n_15936) );
oa22f80 g553468 ( .a(n_15600), .b(FE_OFN307_n_3069), .c(n_587), .d(FE_OFN357_n_4860), .o(n_15934) );
oa22f80 g553469 ( .a(n_16916), .b(FE_OFN413_n_28303), .c(n_1639), .d(FE_OFN1121_rst), .o(n_16433) );
oa22f80 g553470 ( .a(n_16225), .b(FE_OFN201_n_29637), .c(n_1619), .d(FE_OFN80_n_27012), .o(n_16226) );
oa22f80 g553471 ( .a(n_15326), .b(FE_OFN311_n_3069), .c(n_1167), .d(FE_OFN134_n_27449), .o(n_16432) );
oa22f80 g553472 ( .a(FE_OFN628_n_15605), .b(FE_OFN256_n_4280), .c(n_727), .d(n_27709), .o(n_15933) );
ao22s80 g553473 ( .a(n_16455), .b(n_16224), .c(n_15536), .d(x_in_32_1), .o(n_16813) );
oa22f80 g553474 ( .a(n_16222), .b(FE_OFN297_n_3069), .c(n_1146), .d(FE_OFN1121_rst), .o(n_16223) );
oa22f80 g553475 ( .a(n_15873), .b(n_23813), .c(n_299), .d(FE_OFN288_n_29266), .o(n_15932) );
ao22s80 g553476 ( .a(n_16453), .b(n_16221), .c(n_15529), .d(x_in_48_1), .o(n_16817) );
oa22f80 g553477 ( .a(FE_OFN897_n_15930), .b(FE_OFN292_n_3069), .c(n_386), .d(n_29261), .o(n_15931) );
oa22f80 g553478 ( .a(n_16219), .b(FE_OFN410_n_28303), .c(n_1149), .d(n_27709), .o(n_16220) );
ao22s80 g553479 ( .a(n_15000), .b(n_13497), .c(x_out_41_19), .d(FE_OFN271_n_16028), .o(n_15929) );
ao22s80 g553480 ( .a(n_15002), .b(n_13492), .c(x_out_42_19), .d(n_16893), .o(n_15928) );
oa22f80 g553481 ( .a(n_15322), .b(n_23315), .c(n_1505), .d(FE_OFN352_n_4860), .o(n_16431) );
ao22s80 g553482 ( .a(n_14525), .b(n_12314), .c(n_15627), .d(FE_OFN642_n_12432), .o(n_16621) );
oa22f80 g553483 ( .a(FE_OFN831_n_14863), .b(n_23813), .c(n_510), .d(FE_OFN56_n_27012), .o(n_15927) );
ao22s80 g553484 ( .a(n_14532), .b(n_14882), .c(n_15626), .d(n_14881), .o(n_16620) );
ao12f80 g553485 ( .a(n_16398), .b(x_out_60_31), .c(FE_OFN38_n_17184), .o(n_16890) );
ao12f80 g553486 ( .a(n_16402), .b(x_out_61_31), .c(FE_OFN38_n_17184), .o(n_16889) );
ao12f80 g553487 ( .a(n_16400), .b(x_out_63_31), .c(FE_OFN38_n_17184), .o(n_16888) );
ao22s80 g553488 ( .a(n_15706), .b(n_15124), .c(x_out_33_19), .d(FE_OFN277_n_16893), .o(n_16658) );
ao22s80 g553489 ( .a(n_15443), .b(n_8965), .c(x_out_36_19), .d(FE_OFN271_n_16028), .o(n_16430) );
ao22s80 g553490 ( .a(n_15704), .b(n_15100), .c(x_out_39_19), .d(FE_OFN279_n_16656), .o(n_16657) );
ao22s80 g553491 ( .a(n_14539), .b(n_14880), .c(n_15625), .d(n_14879), .o(n_16619) );
ao22s80 g553492 ( .a(n_16444), .b(x_in_4_13), .c(n_23062), .d(n_96), .o(n_24669) );
ao22s80 g553493 ( .a(n_16444), .b(x_in_4_14), .c(n_23062), .d(n_2403), .o(n_24673) );
in01f80 g553494 ( .a(n_16654), .o(n_16655) );
oa22f80 g553495 ( .a(n_23062), .b(n_2112), .c(n_16444), .d(x_in_4_12), .o(n_16654) );
ao22s80 g553496 ( .a(n_14530), .b(n_14877), .c(n_15624), .d(n_14876), .o(n_16616) );
ao22s80 g553497 ( .a(n_14527), .b(n_14856), .c(n_15623), .d(n_14855), .o(n_16615) );
oa22f80 g553498 ( .a(n_14536), .b(n_14534), .c(n_15622), .d(n_14533), .o(n_16613) );
no02f80 g553510 ( .a(n_16368), .b(FE_OFN600_n_16000), .o(n_16429) );
no02f80 g553511 ( .a(n_15922), .b(n_7424), .o(n_15926) );
na02f80 g553512 ( .a(n_15620), .b(x_in_1_12), .o(n_15621) );
no02f80 g553513 ( .a(n_16370), .b(n_16002), .o(n_16428) );
no02f80 g553514 ( .a(n_15924), .b(FE_OFN895_n_15923), .o(n_15925) );
no02f80 g553515 ( .a(n_15922), .b(x_in_39_14), .o(n_16554) );
no02f80 g553516 ( .a(n_16217), .b(FE_OFN690_n_16216), .o(n_16218) );
na02f80 g553517 ( .a(n_16653), .b(n_16025), .o(n_17182) );
no02f80 g553518 ( .a(n_16426), .b(n_16425), .o(n_16427) );
na02f80 g553519 ( .a(n_15960), .b(n_15618), .o(n_15619) );
in01f80 g553520 ( .a(n_15616), .o(n_15617) );
no02f80 g553521 ( .a(n_15241), .b(x_in_24_2), .o(n_15616) );
in01f80 g553522 ( .a(n_16651), .o(n_16652) );
na02f80 g553523 ( .a(n_16424), .b(n_15684), .o(n_16651) );
no02f80 g553524 ( .a(n_15959), .b(n_15614), .o(n_15615) );
na02f80 g553525 ( .a(n_16215), .b(n_15657), .o(n_16697) );
in01f80 g553526 ( .a(n_16213), .o(n_16214) );
no02f80 g553527 ( .a(n_16114), .b(x_in_58_2), .o(n_16213) );
na02f80 g553528 ( .a(n_16699), .b(x_in_38_4), .o(n_16920) );
na02f80 g553529 ( .a(n_16212), .b(x_in_38_3), .o(n_16921) );
in01f80 g553530 ( .a(n_16422), .o(n_16423) );
no02f80 g553531 ( .a(n_16212), .b(x_in_38_3), .o(n_16422) );
na02f80 g553532 ( .a(n_16387), .b(x_in_2_2), .o(n_16551) );
in01f80 g553533 ( .a(n_15920), .o(n_15921) );
no02f80 g553534 ( .a(n_16387), .b(x_in_2_2), .o(n_15920) );
na02f80 g553535 ( .a(n_16151), .b(x_in_22_2), .o(n_16552) );
in01f80 g553536 ( .a(n_15918), .o(n_15919) );
no02f80 g553537 ( .a(n_16151), .b(x_in_22_2), .o(n_15918) );
na02f80 g553538 ( .a(n_16118), .b(x_in_42_2), .o(n_16730) );
in01f80 g553539 ( .a(n_16210), .o(n_16211) );
no02f80 g553540 ( .a(n_16394), .b(x_in_8_4), .o(n_16210) );
no02f80 g553541 ( .a(n_16217), .b(n_14206), .o(n_16704) );
no02f80 g553542 ( .a(n_15916), .b(n_15915), .o(n_15917) );
na02f80 g553543 ( .a(n_16394), .b(x_in_8_4), .o(n_16748) );
in01f80 g553544 ( .a(n_15913), .o(n_15914) );
no02f80 g553545 ( .a(n_16135), .b(x_in_54_2), .o(n_15913) );
no02f80 g553546 ( .a(n_16208), .b(n_16207), .o(n_16209) );
na02f80 g553547 ( .a(n_16148), .b(x_in_14_2), .o(n_16550) );
in01f80 g553548 ( .a(n_15911), .o(n_15912) );
no02f80 g553549 ( .a(n_16148), .b(x_in_14_2), .o(n_15911) );
na02f80 g553550 ( .a(n_16374), .b(x_in_34_2), .o(n_16742) );
in01f80 g553551 ( .a(n_16205), .o(n_16206) );
no02f80 g553552 ( .a(n_16374), .b(x_in_34_2), .o(n_16205) );
no02f80 g553553 ( .a(n_16203), .b(n_16202), .o(n_16204) );
na02f80 g553554 ( .a(n_16145), .b(x_in_46_2), .o(n_16743) );
in01f80 g553555 ( .a(n_16200), .o(n_16201) );
no02f80 g553556 ( .a(n_16145), .b(x_in_46_2), .o(n_16200) );
na02f80 g553557 ( .a(n_15909), .b(n_15908), .o(n_15910) );
na02f80 g553558 ( .a(n_15907), .b(x_in_16_2), .o(n_16741) );
in01f80 g553559 ( .a(n_16198), .o(n_16199) );
no02f80 g553560 ( .a(n_15907), .b(x_in_16_2), .o(n_16198) );
no02f80 g553561 ( .a(n_16196), .b(n_16195), .o(n_16197) );
na02f80 g553562 ( .a(n_16194), .b(x_in_30_2), .o(n_16919) );
in01f80 g553563 ( .a(n_16420), .o(n_16421) );
no02f80 g553564 ( .a(n_16194), .b(x_in_30_2), .o(n_16420) );
na02f80 g553565 ( .a(n_16382), .b(x_in_18_2), .o(n_16736) );
in01f80 g553566 ( .a(n_16192), .o(n_16193) );
no02f80 g553567 ( .a(n_16382), .b(x_in_18_2), .o(n_16192) );
no02f80 g553568 ( .a(n_16190), .b(n_16189), .o(n_16191) );
na02f80 g553569 ( .a(n_16141), .b(x_in_62_2), .o(n_16549) );
in01f80 g553570 ( .a(n_15905), .o(n_15906) );
no02f80 g553571 ( .a(n_16141), .b(x_in_62_2), .o(n_15905) );
na02f80 g553572 ( .a(n_16137), .b(x_in_12_2), .o(n_16288) );
in01f80 g553573 ( .a(n_15612), .o(n_15613) );
no02f80 g553574 ( .a(n_16137), .b(x_in_12_2), .o(n_15612) );
na02f80 g553575 ( .a(n_15611), .b(x_in_0_10), .o(n_16548) );
in01f80 g553576 ( .a(n_15903), .o(n_15904) );
no02f80 g553577 ( .a(n_15611), .b(x_in_0_10), .o(n_15903) );
na02f80 g553578 ( .a(n_15957), .b(n_15609), .o(n_15610) );
in01f80 g553579 ( .a(n_16418), .o(n_16419) );
na02f80 g553580 ( .a(n_16188), .b(n_15659), .o(n_16418) );
no02f80 g553581 ( .a(n_16186), .b(n_16185), .o(n_16187) );
no02f80 g553582 ( .a(n_16416), .b(n_16415), .o(n_16417) );
na02f80 g553583 ( .a(n_16416), .b(n_16008), .o(n_16917) );
na02f80 g553584 ( .a(n_16379), .b(x_in_50_2), .o(n_16545) );
in01f80 g553585 ( .a(n_15901), .o(n_15902) );
no02f80 g553586 ( .a(n_16379), .b(x_in_50_2), .o(n_15901) );
no02f80 g553587 ( .a(n_14555), .b(n_12941), .o(n_16303) );
na02f80 g553588 ( .a(n_15607), .b(n_15606), .o(n_15608) );
na02f80 g553589 ( .a(n_16426), .b(n_16225), .o(n_17070) );
no02f80 g553590 ( .a(n_15924), .b(n_13845), .o(n_16481) );
in01f80 g553591 ( .a(n_16183), .o(n_16184) );
no02f80 g553592 ( .a(n_16117), .b(x_in_26_2), .o(n_16183) );
na02f80 g553593 ( .a(FE_OFN628_n_15605), .b(n_15915), .o(n_16822) );
na02f80 g553594 ( .a(n_15956), .b(n_15603), .o(n_15604) );
na02f80 g553595 ( .a(n_16414), .b(n_15681), .o(n_16907) );
na02f80 g553596 ( .a(n_15871), .b(x_in_44_2), .o(n_16287) );
in01f80 g553597 ( .a(n_15601), .o(n_15602) );
no02f80 g553598 ( .a(n_15871), .b(x_in_44_2), .o(n_15601) );
no02f80 g553599 ( .a(n_15246), .b(n_14986), .o(n_14987) );
na02f80 g553600 ( .a(n_15241), .b(x_in_24_2), .o(n_16286) );
na02f80 g553601 ( .a(n_16182), .b(x_in_28_4), .o(n_16910) );
no02f80 g553602 ( .a(n_15633), .b(n_15239), .o(n_15240) );
na02f80 g553603 ( .a(n_16112), .b(x_in_10_2), .o(n_16731) );
in01f80 g553604 ( .a(n_16180), .o(n_16181) );
no02f80 g553605 ( .a(n_16112), .b(x_in_10_2), .o(n_16180) );
na02f80 g553606 ( .a(n_16135), .b(x_in_54_2), .o(n_16546) );
in01f80 g553607 ( .a(n_16412), .o(n_16413) );
no02f80 g553608 ( .a(n_16182), .b(x_in_28_4), .o(n_16412) );
na02f80 g553609 ( .a(n_15900), .b(x_in_28_3), .o(n_16729) );
in01f80 g553610 ( .a(n_16178), .o(n_16179) );
no02f80 g553611 ( .a(n_15900), .b(x_in_28_3), .o(n_16178) );
na02f80 g553612 ( .a(n_16177), .b(x_in_4_10), .o(n_16913) );
in01f80 g553613 ( .a(n_16410), .o(n_16411) );
no02f80 g553614 ( .a(n_16177), .b(x_in_4_10), .o(n_16410) );
na02f80 g553615 ( .a(n_16445), .b(n_16408), .o(n_16409) );
in01f80 g553616 ( .a(n_16175), .o(n_16176) );
na02f80 g553617 ( .a(n_15899), .b(n_15279), .o(n_16175) );
in01f80 g553618 ( .a(n_16173), .o(n_16174) );
no02f80 g553619 ( .a(n_16118), .b(x_in_42_2), .o(n_16173) );
na02f80 g553620 ( .a(n_16468), .b(n_16171), .o(n_16172) );
no02f80 g553621 ( .a(n_15897), .b(n_15896), .o(n_15898) );
na02f80 g553622 ( .a(n_15600), .b(n_15896), .o(n_16824) );
na02f80 g553623 ( .a(n_15632), .b(n_15237), .o(n_15238) );
in01f80 g553624 ( .a(n_16406), .o(n_16407) );
no02f80 g553625 ( .a(n_16699), .b(x_in_38_4), .o(n_16406) );
na02f80 g553626 ( .a(n_15787), .b(x_in_56_3), .o(n_16540) );
in01f80 g553627 ( .a(n_15894), .o(n_15895) );
no02f80 g553628 ( .a(n_15787), .b(x_in_56_3), .o(n_15894) );
na02f80 g553629 ( .a(n_16117), .b(x_in_26_2), .o(n_16726) );
no02f80 g553630 ( .a(n_16169), .b(n_16168), .o(n_16170) );
na02f80 g553631 ( .a(n_15627), .b(n_15235), .o(n_15236) );
na02f80 g553632 ( .a(n_15626), .b(n_15598), .o(n_15599) );
na02f80 g553633 ( .a(n_16114), .b(x_in_58_2), .o(n_16735) );
na02f80 g553634 ( .a(n_15625), .b(n_15596), .o(n_15597) );
no02f80 g553635 ( .a(n_16166), .b(x_in_15_14), .o(n_16167) );
no02f80 g553636 ( .a(n_16164), .b(x_in_63_14), .o(n_16165) );
no02f80 g553637 ( .a(n_16162), .b(x_in_47_14), .o(n_16163) );
in01f80 g553638 ( .a(n_15893), .o(n_16530) );
na02f80 g553639 ( .a(n_15620), .b(n_1808), .o(n_15893) );
na02f80 g553640 ( .a(n_16016), .b(n_16158), .o(n_16405) );
na02f80 g553641 ( .a(n_16014), .b(n_16156), .o(n_16404) );
na02f80 g553642 ( .a(n_16242), .b(n_15891), .o(n_15892) );
na02f80 g553643 ( .a(n_16020), .b(n_16154), .o(n_16403) );
na02f80 g553644 ( .a(n_15009), .b(n_15590), .o(n_15888) );
no02f80 g553645 ( .a(n_15886), .b(n_15885), .o(n_15887) );
na02f80 g553646 ( .a(n_15886), .b(n_15715), .o(n_16536) );
na02f80 g553647 ( .a(n_15954), .b(n_15594), .o(n_15595) );
no02f80 g553648 ( .a(n_16401), .b(n_7406), .o(n_16402) );
no02f80 g553649 ( .a(n_16399), .b(n_8198), .o(n_16400) );
no02f80 g553650 ( .a(n_16397), .b(n_8056), .o(n_16398) );
na02f80 g553651 ( .a(n_15922), .b(n_2343), .o(n_15884) );
no02f80 g553652 ( .a(n_15592), .b(n_12169), .o(n_15593) );
na02f80 g553653 ( .a(n_16466), .b(n_16160), .o(n_16161) );
na02f80 g553654 ( .a(n_15882), .b(n_15881), .o(n_15883) );
no02f80 g553655 ( .a(n_15631), .b(n_15233), .o(n_15234) );
na02f80 g553656 ( .a(n_15952), .b(n_15879), .o(n_15880) );
na02f80 g553657 ( .a(n_16159), .b(n_16158), .o(n_16723) );
na02f80 g553658 ( .a(n_16157), .b(n_16156), .o(n_16721) );
na02f80 g553659 ( .a(n_16155), .b(n_16154), .o(n_16719) );
na02f80 g553660 ( .a(n_15591), .b(n_15590), .o(n_16281) );
no02f80 g553661 ( .a(n_15592), .b(n_15588), .o(n_15589) );
no02f80 g553662 ( .a(n_15245), .b(n_14984), .o(n_14985) );
na02f80 g553663 ( .a(n_16152), .b(n_16151), .o(n_16153) );
na02f80 g553664 ( .a(n_16150), .b(n_15074), .o(n_17549) );
na02f80 g553665 ( .a(n_16150), .b(n_16148), .o(n_16149) );
na02f80 g553666 ( .a(n_16147), .b(n_15327), .o(n_17546) );
na02f80 g553667 ( .a(n_16147), .b(n_16145), .o(n_16146) );
na02f80 g553668 ( .a(n_16393), .b(n_16194), .o(n_16144) );
na02f80 g553669 ( .a(n_16143), .b(n_15068), .o(n_17550) );
na02f80 g553670 ( .a(n_16143), .b(n_16141), .o(n_16142) );
na02f80 g553671 ( .a(n_16140), .b(n_15077), .o(n_17547) );
no02f80 g553672 ( .a(n_15875), .b(n_16035), .o(n_15876) );
no02f80 g553673 ( .a(n_15875), .b(n_15018), .o(n_16534) );
na02f80 g553674 ( .a(n_16395), .b(n_16394), .o(n_16396) );
na02f80 g553675 ( .a(n_16138), .b(n_16137), .o(n_16139) );
na02f80 g553676 ( .a(n_16393), .b(n_15685), .o(n_17545) );
na02f80 g553677 ( .a(n_16395), .b(n_15321), .o(n_17031) );
na02f80 g553678 ( .a(n_16140), .b(n_16135), .o(n_16136) );
na02f80 g553679 ( .a(n_16152), .b(n_15071), .o(n_17548) );
na02f80 g553680 ( .a(n_16138), .b(n_14878), .o(n_17544) );
na02f80 g553681 ( .a(n_15624), .b(n_15586), .o(n_15587) );
na02f80 g553682 ( .a(n_15623), .b(n_15584), .o(n_15585) );
na02f80 g553683 ( .a(n_16389), .b(x_in_60_1), .o(n_17216) );
na02f80 g553684 ( .a(n_16392), .b(x_in_6_1), .o(n_17210) );
no02f80 g553685 ( .a(n_16392), .b(x_in_6_1), .o(n_17209) );
na02f80 g553686 ( .a(n_15874), .b(n_15873), .o(n_16584) );
na02f80 g553687 ( .a(n_16134), .b(x_in_52_1), .o(n_16951) );
no02f80 g553688 ( .a(n_16134), .b(x_in_52_1), .o(n_16950) );
na02f80 g553689 ( .a(n_16391), .b(x_in_48_1), .o(n_17204) );
no02f80 g553690 ( .a(n_16391), .b(x_in_48_1), .o(n_17203) );
na02f80 g553691 ( .a(n_16390), .b(x_in_40_1), .o(n_17206) );
no02f80 g553692 ( .a(n_16390), .b(x_in_40_1), .o(n_17205) );
na02f80 g553693 ( .a(n_16133), .b(x_in_32_1), .o(n_16955) );
no02f80 g553694 ( .a(n_16133), .b(x_in_32_1), .o(n_16954) );
no02f80 g553695 ( .a(n_16389), .b(x_in_60_1), .o(n_17215) );
na02f80 g553696 ( .a(n_16650), .b(x_in_20_1), .o(n_17505) );
no02f80 g553697 ( .a(n_16650), .b(x_in_20_1), .o(n_17504) );
no02f80 g553698 ( .a(n_16388), .b(x_in_36_1), .o(n_17509) );
na02f80 g553699 ( .a(n_16388), .b(x_in_36_1), .o(n_17510) );
na02f80 g553700 ( .a(n_15874), .b(n_15871), .o(n_15872) );
na02f80 g553701 ( .a(n_15629), .b(n_15231), .o(n_15232) );
no02f80 g553702 ( .a(n_15869), .b(n_15868), .o(n_15870) );
na02f80 g553703 ( .a(n_15582), .b(n_15581), .o(n_15583) );
na02f80 g553704 ( .a(n_15866), .b(n_15865), .o(n_15867) );
na02f80 g553705 ( .a(n_15622), .b(n_15226), .o(n_15227) );
na02f80 g553706 ( .a(n_15311), .b(n_16132), .o(n_16706) );
na02f80 g553707 ( .a(n_15900), .b(n_16132), .o(n_15864) );
no02f80 g553708 ( .a(n_15630), .b(n_15224), .o(n_15225) );
no02f80 g553709 ( .a(n_14857), .b(n_15579), .o(n_16581) );
no02f80 g553710 ( .a(n_15937), .b(n_15579), .o(n_15580) );
no02f80 g553711 ( .a(n_16212), .b(n_16131), .o(n_16701) );
na02f80 g553712 ( .a(n_15862), .b(n_16131), .o(n_15863) );
na02f80 g553713 ( .a(n_15953), .b(n_15577), .o(n_15578) );
no02f80 g553714 ( .a(n_15575), .b(n_15754), .o(n_15576) );
no02f80 g553715 ( .a(n_14982), .b(n_14981), .o(n_14983) );
in01f80 g553716 ( .a(n_15573), .o(n_15574) );
no02f80 g553717 ( .a(n_15223), .b(n_15222), .o(n_15573) );
na02f80 g553718 ( .a(n_15223), .b(n_15222), .o(n_16269) );
na02f80 g553719 ( .a(n_15531), .b(n_15530), .o(n_16498) );
in01f80 g553720 ( .a(n_16129), .o(n_16130) );
no02f80 g553721 ( .a(n_15336), .b(n_13025), .o(n_16129) );
no02f80 g553722 ( .a(n_15571), .b(n_9364), .o(n_15572) );
oa12f80 g553723 ( .a(FE_OFN391_n_15554), .b(n_654), .c(n_29264), .o(n_15570) );
no02f80 g553724 ( .a(n_15700), .b(n_16387), .o(n_17247) );
no02f80 g553725 ( .a(n_15337), .b(n_13026), .o(n_16693) );
na02f80 g553726 ( .a(n_15180), .b(n_15861), .o(n_25185) );
in01f80 g553727 ( .a(n_16127), .o(n_16128) );
na02f80 g553728 ( .a(n_15332), .b(n_15012), .o(n_16127) );
no02f80 g553729 ( .a(n_15079), .b(n_14186), .o(n_16496) );
oa12f80 g553730 ( .a(FE_OFN373_n_15853), .b(n_286), .c(FE_OFN1110_rst), .o(n_15860) );
in01f80 g553731 ( .a(n_16385), .o(n_16386) );
no02f80 g553732 ( .a(n_15687), .b(n_14162), .o(n_16385) );
in01f80 g553733 ( .a(n_15858), .o(n_15859) );
na02f80 g553734 ( .a(n_15043), .b(n_14134), .o(n_15858) );
no02f80 g553735 ( .a(n_15688), .b(n_14163), .o(n_16904) );
in01f80 g553736 ( .a(n_15856), .o(n_15857) );
na02f80 g553737 ( .a(n_15075), .b(n_14609), .o(n_15856) );
oa12f80 g553738 ( .a(n_15213), .b(n_190), .c(FE_OFN1124_rst), .o(n_15221) );
in01f80 g553739 ( .a(n_16649), .o(n_17249) );
na02f80 g553740 ( .a(n_16384), .b(n_15324), .o(n_16649) );
na02f80 g553741 ( .a(n_16384), .b(n_16382), .o(n_16383) );
na02f80 g553742 ( .a(n_15076), .b(n_14610), .o(n_16495) );
in01f80 g553743 ( .a(n_16125), .o(n_16126) );
no02f80 g553744 ( .a(n_15334), .b(n_13815), .o(n_16125) );
no02f80 g553745 ( .a(n_15335), .b(n_13816), .o(n_16690) );
in01f80 g553746 ( .a(n_15568), .o(n_15569) );
na02f80 g553747 ( .a(n_14874), .b(n_13813), .o(n_15568) );
no02f80 g553748 ( .a(n_15219), .b(n_15218), .o(n_16267) );
no02f80 g553749 ( .a(n_15548), .b(n_15547), .o(n_16494) );
in01f80 g553750 ( .a(n_15566), .o(n_15567) );
na02f80 g553751 ( .a(n_14894), .b(n_13811), .o(n_15566) );
oa12f80 g553752 ( .a(FE_OFN371_n_15817), .b(n_822), .c(FE_OFN116_n_27449), .o(n_15855) );
in01f80 g553753 ( .a(n_16648), .o(n_17238) );
na02f80 g553754 ( .a(n_15067), .b(n_16381), .o(n_16648) );
no02f80 g553755 ( .a(n_15212), .b(n_15211), .o(n_16253) );
na02f80 g553756 ( .a(n_16379), .b(n_16381), .o(n_16380) );
no02f80 g553757 ( .a(n_15080), .b(n_14187), .o(n_16497) );
oa12f80 g553758 ( .a(FE_OFN373_n_15853), .b(n_241), .c(FE_OFN91_n_27449), .o(n_15854) );
no02f80 g553759 ( .a(n_15949), .b(n_15948), .o(n_15220) );
in01f80 g553760 ( .a(n_15564), .o(n_15565) );
na02f80 g553761 ( .a(n_15219), .b(n_15218), .o(n_15564) );
oa12f80 g553762 ( .a(n_15790), .b(n_272), .c(FE_OFN136_n_27449), .o(n_15852) );
in01f80 g553763 ( .a(n_16378), .o(n_16975) );
na02f80 g553764 ( .a(n_16124), .b(n_15312), .o(n_16378) );
na02f80 g553765 ( .a(n_16374), .b(n_16122), .o(n_16123) );
no02f80 g553766 ( .a(n_15217), .b(n_15216), .o(n_16268) );
no02f80 g553767 ( .a(n_15804), .b(n_15803), .o(n_16689) );
in01f80 g553768 ( .a(n_15562), .o(n_15563) );
na02f80 g553769 ( .a(n_14892), .b(n_13771), .o(n_15562) );
na02f80 g553770 ( .a(n_15425), .b(n_16121), .o(n_24898) );
in01f80 g553771 ( .a(n_15560), .o(n_15561) );
na02f80 g553772 ( .a(n_15217), .b(n_15216), .o(n_15560) );
in01f80 g553773 ( .a(n_16377), .o(n_16997) );
na02f80 g553774 ( .a(n_16120), .b(n_15310), .o(n_16377) );
na02f80 g553775 ( .a(n_16120), .b(n_16118), .o(n_16119) );
no02f80 g553776 ( .a(n_15167), .b(n_15851), .o(n_23212) );
na02f80 g553777 ( .a(n_15850), .b(n_15849), .o(n_26585) );
oa12f80 g553778 ( .a(n_15773), .b(n_387), .c(FE_OFN105_n_27449), .o(n_15848) );
na02f80 g553779 ( .a(n_14893), .b(n_13772), .o(n_16266) );
no02f80 g553780 ( .a(n_15417), .b(n_16117), .o(n_17266) );
in01f80 g553781 ( .a(n_15558), .o(n_15559) );
na02f80 g553782 ( .a(n_14890), .b(n_13817), .o(n_15558) );
in01f80 g553783 ( .a(n_15556), .o(n_15557) );
no02f80 g553784 ( .a(n_14843), .b(n_13819), .o(n_15556) );
in01f80 g553785 ( .a(n_16376), .o(n_16993) );
na02f80 g553786 ( .a(n_16116), .b(n_15298), .o(n_16376) );
oa12f80 g553787 ( .a(n_15554), .b(n_714), .c(FE_OFN69_n_27012), .o(n_15555) );
no02f80 g553788 ( .a(n_15507), .b(n_15847), .o(n_25621) );
na02f80 g553789 ( .a(n_15845), .b(n_16117), .o(n_15846) );
in01f80 g553790 ( .a(n_15552), .o(n_15553) );
na02f80 g553791 ( .a(n_14888), .b(n_13821), .o(n_15552) );
in01f80 g553792 ( .a(n_15550), .o(n_15551) );
no02f80 g553793 ( .a(n_14861), .b(n_13828), .o(n_15550) );
na02f80 g553794 ( .a(n_14889), .b(n_13822), .o(n_16244) );
no02f80 g553795 ( .a(n_14862), .b(n_13829), .o(n_16265) );
na02f80 g553796 ( .a(n_15207), .b(n_15206), .o(n_16260) );
no02f80 g553797 ( .a(n_15516), .b(n_15515), .o(n_16474) );
na02f80 g553798 ( .a(n_14959), .b(n_15549), .o(n_24171) );
na02f80 g553799 ( .a(n_15165), .b(n_15844), .o(n_23859) );
no02f80 g553800 ( .a(n_15419), .b(n_15843), .o(n_24894) );
no02f80 g553801 ( .a(n_15488), .b(n_15487), .o(n_16490) );
na02f80 g553802 ( .a(n_16116), .b(n_16114), .o(n_16115) );
no02f80 g553803 ( .a(n_14844), .b(n_13820), .o(n_16261) );
in01f80 g553804 ( .a(n_15841), .o(n_15842) );
na02f80 g553805 ( .a(n_15548), .b(n_15547), .o(n_15841) );
no02f80 g553806 ( .a(n_14938), .b(n_15546), .o(n_24201) );
na02f80 g553807 ( .a(n_25728), .b(n_15840), .o(n_25356) );
no02f80 g553808 ( .a(n_15162), .b(n_15839), .o(n_22924) );
na02f80 g553809 ( .a(n_14956), .b(n_15545), .o(n_23880) );
no02f80 g553810 ( .a(n_15356), .b(n_15838), .o(n_24697) );
no02f80 g553811 ( .a(n_15571), .b(n_15837), .o(n_25686) );
oa12f80 g553812 ( .a(n_14994), .b(n_581), .c(n_29068), .o(n_15215) );
oa12f80 g553813 ( .a(n_16372), .b(n_622), .c(FE_OFN361_n_4860), .o(n_16375) );
na02f80 g553814 ( .a(n_14875), .b(n_13814), .o(n_16262) );
no02f80 g553815 ( .a(n_15158), .b(n_15836), .o(n_22922) );
na02f80 g553816 ( .a(n_14954), .b(n_15544), .o(n_23878) );
no02f80 g553817 ( .a(n_15401), .b(n_15835), .o(n_24648) );
in01f80 g553818 ( .a(n_15833), .o(n_15834) );
no02f80 g553819 ( .a(n_15069), .b(n_14148), .o(n_15833) );
na02f80 g553820 ( .a(n_15148), .b(n_15832), .o(n_24161) );
na02f80 g553821 ( .a(n_16124), .b(n_16112), .o(n_16113) );
in01f80 g553822 ( .a(n_15830), .o(n_15831) );
no02f80 g553823 ( .a(n_15072), .b(n_13846), .o(n_15830) );
no02f80 g553824 ( .a(n_15073), .b(n_13847), .o(n_16487) );
no02f80 g553825 ( .a(n_15146), .b(n_15829), .o(n_22920) );
na02f80 g553826 ( .a(n_14949), .b(n_15543), .o(n_23876) );
no02f80 g553827 ( .a(n_15391), .b(n_15828), .o(n_24563) );
oa12f80 g553828 ( .a(n_15534), .b(n_674), .c(FE_OFN136_n_27449), .o(n_15542) );
no02f80 g553829 ( .a(n_15827), .b(n_14858), .o(n_16782) );
oa12f80 g553830 ( .a(n_15213), .b(n_1617), .c(n_28928), .o(n_15214) );
no02f80 g553831 ( .a(n_15134), .b(n_15826), .o(n_22916) );
na02f80 g553832 ( .a(n_14947), .b(n_15541), .o(n_23872) );
no02f80 g553833 ( .a(n_15379), .b(n_15825), .o(n_24554) );
no02f80 g553834 ( .a(n_15127), .b(n_15824), .o(n_23863) );
no02f80 g553835 ( .a(n_15539), .b(n_15538), .o(n_15540) );
no02f80 g553836 ( .a(n_15125), .b(n_15823), .o(n_22914) );
na02f80 g553837 ( .a(n_14939), .b(n_15537), .o(n_23870) );
no02f80 g553838 ( .a(n_15361), .b(n_15822), .o(n_24552) );
in01f80 g553839 ( .a(n_16792), .o(n_15821) );
no02f80 g553840 ( .a(n_15536), .b(n_15819), .o(n_16792) );
no02f80 g553841 ( .a(n_16455), .b(n_15819), .o(n_15820) );
oa12f80 g553842 ( .a(FE_OFN371_n_15817), .b(n_604), .c(FE_OFN353_n_4860), .o(n_15818) );
no02f80 g553843 ( .a(n_15815), .b(n_16222), .o(n_15816) );
no02f80 g553844 ( .a(n_15815), .b(n_15056), .o(n_16576) );
oa12f80 g553845 ( .a(n_15534), .b(n_221), .c(FE_OFN136_n_27449), .o(n_15535) );
no02f80 g553846 ( .a(n_15123), .b(n_15907), .o(n_17248) );
in01f80 g553847 ( .a(n_15532), .o(n_15533) );
no02f80 g553848 ( .a(n_14849), .b(n_13776), .o(n_15532) );
na02f80 g553849 ( .a(n_15813), .b(n_15907), .o(n_15814) );
in01f80 g553850 ( .a(n_15811), .o(n_15812) );
no02f80 g553851 ( .a(n_15531), .b(n_15530), .o(n_15811) );
na02f80 g553852 ( .a(n_15118), .b(n_15809), .o(n_23849) );
no02f80 g553853 ( .a(n_15529), .b(n_15807), .o(n_17401) );
no02f80 g553854 ( .a(n_16453), .b(n_15807), .o(n_15808) );
in01f80 g553855 ( .a(n_15805), .o(n_15806) );
no02f80 g553856 ( .a(n_15065), .b(n_13823), .o(n_15805) );
no02f80 g553857 ( .a(n_15070), .b(n_14149), .o(n_16493) );
no02f80 g553858 ( .a(n_15066), .b(n_13824), .o(n_16483) );
na02f80 g553859 ( .a(n_14895), .b(n_13812), .o(n_16264) );
na02f80 g553860 ( .a(n_15064), .b(n_12259), .o(n_16772) );
oa12f80 g553861 ( .a(n_16082), .b(n_1281), .c(FE_OFN193_n_28928), .o(n_16110) );
no02f80 g553862 ( .a(n_16374), .b(n_15693), .o(n_17242) );
na02f80 g553863 ( .a(n_15528), .b(n_15527), .o(n_16479) );
no02f80 g553864 ( .a(n_15514), .b(n_15513), .o(n_16478) );
in01f80 g553865 ( .a(n_16108), .o(n_16109) );
na02f80 g553866 ( .a(n_15804), .b(n_15803), .o(n_16108) );
in01f80 g553867 ( .a(n_15801), .o(n_15802) );
no02f80 g553868 ( .a(n_15528), .b(n_15527), .o(n_15801) );
in01f80 g553869 ( .a(n_15525), .o(n_15526) );
no02f80 g553870 ( .a(n_14872), .b(n_13841), .o(n_15525) );
no02f80 g553871 ( .a(n_14873), .b(n_13842), .o(n_16259) );
in01f80 g553872 ( .a(n_15799), .o(n_15800) );
na02f80 g553873 ( .a(n_15061), .b(n_13794), .o(n_15799) );
na02f80 g553874 ( .a(n_15062), .b(n_13795), .o(n_16475) );
in01f80 g553875 ( .a(n_15523), .o(n_15524) );
no02f80 g553876 ( .a(n_14870), .b(n_13792), .o(n_15523) );
no02f80 g553877 ( .a(n_14871), .b(n_13793), .o(n_16255) );
in01f80 g553878 ( .a(n_15521), .o(n_15522) );
na02f80 g553879 ( .a(n_14868), .b(n_13790), .o(n_15521) );
na02f80 g553880 ( .a(n_14869), .b(n_13791), .o(n_16258) );
in01f80 g553881 ( .a(n_15519), .o(n_15520) );
no02f80 g553882 ( .a(n_14866), .b(n_13788), .o(n_15519) );
no02f80 g553883 ( .a(n_14867), .b(n_13789), .o(n_16257) );
in01f80 g553884 ( .a(n_15517), .o(n_15518) );
na02f80 g553885 ( .a(n_14859), .b(n_13839), .o(n_15517) );
in01f80 g553886 ( .a(n_16787), .o(n_16107) );
no02f80 g553887 ( .a(n_15798), .b(n_16105), .o(n_16787) );
na02f80 g553888 ( .a(n_14860), .b(n_13840), .o(n_16256) );
in01f80 g553889 ( .a(n_15796), .o(n_15797) );
na02f80 g553890 ( .a(n_15516), .b(n_15515), .o(n_15796) );
in01f80 g553891 ( .a(n_15794), .o(n_15795) );
na02f80 g553892 ( .a(n_15514), .b(n_15513), .o(n_15794) );
in01f80 g553893 ( .a(n_15792), .o(n_15793) );
na02f80 g553894 ( .a(n_15057), .b(n_13014), .o(n_15792) );
no02f80 g553895 ( .a(n_16663), .b(n_16105), .o(n_16106) );
in01f80 g553896 ( .a(n_15511), .o(n_15512) );
no02f80 g553897 ( .a(n_14864), .b(n_13843), .o(n_15511) );
no02f80 g553898 ( .a(n_14865), .b(n_13844), .o(n_16254) );
in01f80 g553899 ( .a(n_16103), .o(n_16104) );
no02f80 g553900 ( .a(n_15319), .b(n_13009), .o(n_16103) );
no02f80 g553901 ( .a(n_15320), .b(n_13008), .o(n_16682) );
na02f80 g553902 ( .a(n_15058), .b(n_13013), .o(n_16472) );
in01f80 g553903 ( .a(n_16101), .o(n_16102) );
na02f80 g553904 ( .a(n_15317), .b(n_14606), .o(n_16101) );
na02f80 g553905 ( .a(n_15318), .b(n_14607), .o(n_16681) );
in01f80 g553906 ( .a(n_16099), .o(n_16100) );
no02f80 g553907 ( .a(n_15315), .b(n_14604), .o(n_16099) );
no02f80 g553908 ( .a(n_15316), .b(n_14605), .o(n_16680) );
in01f80 g553909 ( .a(n_16097), .o(n_16098) );
na02f80 g553910 ( .a(n_15313), .b(n_13362), .o(n_16097) );
oa12f80 g553911 ( .a(n_15790), .b(n_147), .c(FE_OFN136_n_27449), .o(n_15791) );
na02f80 g553912 ( .a(n_15314), .b(n_13363), .o(n_16679) );
in01f80 g553913 ( .a(n_15509), .o(n_15510) );
na02f80 g553914 ( .a(n_15212), .b(n_15211), .o(n_15509) );
in01f80 g553915 ( .a(n_16572), .o(n_16096) );
na02f80 g553916 ( .a(n_15789), .b(n_15055), .o(n_16572) );
na02f80 g553917 ( .a(n_15789), .b(n_15787), .o(n_15788) );
no02f80 g553918 ( .a(n_15827), .b(n_15935), .o(n_15786) );
no02f80 g553919 ( .a(n_15096), .b(n_15785), .o(n_23857) );
in01f80 g553920 ( .a(n_15783), .o(n_15784) );
na02f80 g553921 ( .a(n_15053), .b(n_13837), .o(n_15783) );
na02f80 g553922 ( .a(n_15054), .b(n_13838), .o(n_16473) );
no02f80 g553923 ( .a(n_15507), .b(n_10131), .o(n_15508) );
na02f80 g553924 ( .a(n_16233), .b(n_16232), .o(n_15506) );
in01f80 g553925 ( .a(n_15781), .o(n_15782) );
na02f80 g553926 ( .a(n_15051), .b(n_13782), .o(n_15781) );
na02f80 g553927 ( .a(n_15052), .b(n_13783), .o(n_16488) );
in01f80 g553928 ( .a(n_15779), .o(n_15780) );
na02f80 g553929 ( .a(n_15049), .b(n_13780), .o(n_15779) );
no02f80 g553930 ( .a(n_15090), .b(n_15778), .o(n_23855) );
na02f80 g553931 ( .a(n_15050), .b(n_13781), .o(n_16471) );
in01f80 g553932 ( .a(n_15504), .o(n_15505) );
no02f80 g553933 ( .a(n_14853), .b(n_13778), .o(n_15504) );
no02f80 g553934 ( .a(n_14854), .b(n_13779), .o(n_16252) );
in01f80 g553935 ( .a(n_15502), .o(n_15503) );
na02f80 g553936 ( .a(n_14851), .b(n_13360), .o(n_15502) );
na02f80 g553937 ( .a(n_14852), .b(n_13361), .o(n_16251) );
in01f80 g553938 ( .a(n_15776), .o(n_15777) );
na02f80 g553939 ( .a(n_15047), .b(n_13835), .o(n_15776) );
no02f80 g553940 ( .a(n_14850), .b(n_13777), .o(n_16250) );
in01f80 g553941 ( .a(n_15500), .o(n_15501) );
na02f80 g553942 ( .a(n_14847), .b(n_14600), .o(n_15500) );
na02f80 g553943 ( .a(n_15048), .b(n_13836), .o(n_16470) );
na02f80 g553944 ( .a(n_14848), .b(n_14601), .o(n_16247) );
in01f80 g553945 ( .a(n_16094), .o(n_16095) );
no02f80 g553946 ( .a(n_15308), .b(n_14614), .o(n_16094) );
no02f80 g553947 ( .a(n_15498), .b(n_15775), .o(n_25619) );
no02f80 g553948 ( .a(n_15309), .b(n_14615), .o(n_16683) );
in01f80 g553949 ( .a(n_16092), .o(n_16093) );
na02f80 g553950 ( .a(n_15306), .b(n_12975), .o(n_16092) );
na02f80 g553951 ( .a(n_15307), .b(n_12976), .o(n_16691) );
no02f80 g553952 ( .a(n_15498), .b(n_10129), .o(n_15499) );
no02f80 g553953 ( .a(n_15210), .b(n_15209), .o(n_16249) );
in01f80 g553954 ( .a(n_15496), .o(n_15497) );
na02f80 g553955 ( .a(n_15210), .b(n_15209), .o(n_15496) );
in01f80 g553956 ( .a(n_15494), .o(n_15495) );
na02f80 g553957 ( .a(n_14845), .b(n_13364), .o(n_15494) );
na02f80 g553958 ( .a(n_15493), .b(n_14922), .o(n_24538) );
na02f80 g553959 ( .a(n_14846), .b(n_13365), .o(n_16248) );
oa12f80 g553960 ( .a(n_15773), .b(n_1329), .c(n_29204), .o(n_15774) );
oa12f80 g553961 ( .a(n_16372), .b(n_527), .c(FE_OFN139_n_27449), .o(n_16373) );
no02f80 g553962 ( .a(n_15491), .b(n_15490), .o(n_15492) );
na02f80 g553963 ( .a(n_15766), .b(n_15765), .o(n_16677) );
na02f80 g553964 ( .a(n_14891), .b(n_13818), .o(n_16263) );
no02f80 g553965 ( .a(n_15087), .b(n_15772), .o(n_23851) );
in01f80 g553966 ( .a(n_16795), .o(n_15771) );
no02f80 g553967 ( .a(n_15489), .b(n_15769), .o(n_16795) );
no02f80 g553968 ( .a(n_16441), .b(n_15769), .o(n_15770) );
in01f80 g553969 ( .a(n_15767), .o(n_15768) );
na02f80 g553970 ( .a(n_15045), .b(n_13833), .o(n_15767) );
in01f80 g553971 ( .a(n_16090), .o(n_16091) );
no02f80 g553972 ( .a(n_15766), .b(n_15765), .o(n_16090) );
in01f80 g553973 ( .a(n_15763), .o(n_15764) );
na02f80 g553974 ( .a(n_15488), .b(n_15487), .o(n_15763) );
in01f80 g553975 ( .a(n_16088), .o(n_16089) );
no02f80 g553976 ( .a(n_15303), .b(n_14136), .o(n_16088) );
na02f80 g553977 ( .a(n_15046), .b(n_13834), .o(n_16469) );
no02f80 g553978 ( .a(n_15485), .b(n_15762), .o(n_25607) );
no02f80 g553979 ( .a(n_15304), .b(n_14137), .o(n_16674) );
no02f80 g553980 ( .a(n_15485), .b(n_10127), .o(n_15486) );
na02f80 g553981 ( .a(n_15044), .b(n_14135), .o(n_16492) );
in01f80 g553982 ( .a(n_16086), .o(n_16087) );
no02f80 g553983 ( .a(n_15301), .b(n_14598), .o(n_16086) );
na02f80 g553984 ( .a(n_16084), .b(n_16387), .o(n_16085) );
no02f80 g553985 ( .a(n_15302), .b(n_14599), .o(n_16688) );
oa12f80 g553986 ( .a(n_16082), .b(n_1622), .c(FE_OFN1110_rst), .o(n_16083) );
in01f80 g553987 ( .a(n_16080), .o(n_16081) );
na02f80 g553988 ( .a(n_15299), .b(n_14132), .o(n_16080) );
na02f80 g553989 ( .a(n_15333), .b(n_15013), .o(n_16678) );
na02f80 g553990 ( .a(n_15300), .b(n_14133), .o(n_16673) );
in01f80 g553991 ( .a(n_15760), .o(n_15761) );
no02f80 g553992 ( .a(n_15041), .b(n_13809), .o(n_15760) );
no02f80 g553993 ( .a(n_15042), .b(n_13810), .o(n_16491) );
in01f80 g553994 ( .a(n_15483), .o(n_15484) );
na02f80 g553995 ( .a(n_14841), .b(n_13773), .o(n_15483) );
na02f80 g553996 ( .a(n_14842), .b(n_13774), .o(n_16245) );
no02f80 g553997 ( .a(n_15083), .b(n_15759), .o(n_23865) );
no02f80 g553998 ( .a(n_15945), .b(n_15944), .o(n_15208) );
in01f80 g553999 ( .a(n_15481), .o(n_15482) );
no02f80 g554000 ( .a(n_15207), .b(n_15206), .o(n_15481) );
ao12f80 g554001 ( .a(n_12477), .b(n_15205), .c(n_13673), .o(n_16302) );
in01f80 g554002 ( .a(n_15204), .o(n_16299) );
oa12f80 g554003 ( .a(n_3224), .b(n_14976), .c(n_2160), .o(n_15204) );
oa12f80 g554004 ( .a(n_14999), .b(n_378), .c(FE_OFN1112_rst), .o(n_15203) );
in01f80 g554005 ( .a(n_15480), .o(n_16559) );
oa12f80 g554006 ( .a(n_12548), .b(n_15194), .c(n_11617), .o(n_15480) );
in01f80 g554007 ( .a(n_15202), .o(n_16295) );
oa12f80 g554008 ( .a(n_3153), .b(n_14974), .c(n_2173), .o(n_15202) );
in01f80 g554009 ( .a(n_15479), .o(n_16562) );
oa12f80 g554010 ( .a(n_12131), .b(n_15196), .c(n_10977), .o(n_15479) );
oa12f80 g554011 ( .a(n_15001), .b(n_759), .c(FE_OFN80_n_27012), .o(n_15201) );
oa12f80 g554012 ( .a(n_15755), .b(n_1539), .c(rst), .o(n_15758) );
oa12f80 g554013 ( .a(n_16645), .b(n_1410), .c(FE_OFN139_n_27449), .o(n_16647) );
oa12f80 g554014 ( .a(n_15442), .b(n_1331), .c(FE_OFN355_n_4860), .o(n_15757) );
oa12f80 g554015 ( .a(n_15755), .b(n_872), .c(FE_OFN93_n_27449), .o(n_15756) );
oa12f80 g554016 ( .a(n_14840), .b(n_13099), .c(n_12814), .o(n_15478) );
oa12f80 g554017 ( .a(n_15440), .b(n_1761), .c(n_25680), .o(n_16079) );
oa12f80 g554018 ( .a(n_15703), .b(n_1770), .c(FE_OFN353_n_4860), .o(n_16078) );
oa12f80 g554019 ( .a(n_16645), .b(n_259), .c(FE_OFN139_n_27449), .o(n_16646) );
oa12f80 g554020 ( .a(n_16370), .b(n_1895), .c(FE_OFN141_n_27449), .o(n_16371) );
oa12f80 g554021 ( .a(n_16368), .b(n_1077), .c(FE_OFN1124_rst), .o(n_16369) );
oa12f80 g554022 ( .a(n_15705), .b(n_1969), .c(FE_OFN142_n_27449), .o(n_16077) );
oa12f80 g554023 ( .a(n_15438), .b(n_13), .c(FE_OFN352_n_4860), .o(n_16076) );
oa12f80 g554024 ( .a(n_15702), .b(n_707), .c(FE_OFN190_n_28362), .o(n_16367) );
ao12f80 g554025 ( .a(n_11700), .b(n_13489), .c(n_5264), .o(n_14990) );
ao12f80 g554026 ( .a(n_10803), .b(n_14581), .c(n_12049), .o(n_15640) );
oa12f80 g554027 ( .a(n_3117), .b(n_14079), .c(n_6461), .o(n_15257) );
in01f80 g554028 ( .a(n_16074), .o(n_16075) );
ao12f80 g554029 ( .a(n_16444), .b(x_in_4_13), .c(x_in_4_12), .o(n_16074) );
in01f80 g554030 ( .a(n_16803), .o(n_16073) );
ao12f80 g554031 ( .a(n_14057), .b(n_14992), .c(n_15754), .o(n_16803) );
ao12f80 g554032 ( .a(n_8378), .b(n_15753), .c(n_9553), .o(n_16773) );
ao12f80 g554033 ( .a(n_11516), .b(n_14978), .c(n_12494), .o(n_15983) );
ao12f80 g554034 ( .a(n_11577), .b(n_15477), .c(n_12512), .o(n_16565) );
oa12f80 g554035 ( .a(n_10809), .b(n_15476), .c(n_12051), .o(n_16579) );
in01f80 g554036 ( .a(n_16071), .o(n_16072) );
ao12f80 g554037 ( .a(n_16444), .b(n_15329), .c(n_15752), .o(n_16071) );
oa12f80 g554038 ( .a(n_14924), .b(n_14309), .c(n_14308), .o(n_16271) );
na03f80 g554039 ( .a(n_2394), .b(n_15005), .c(FE_OFN35_n_15183), .o(n_15967) );
in01f80 g554040 ( .a(FE_OFN748_n_16529), .o(n_16070) );
ao22s80 g554041 ( .a(n_15654), .b(n_12065), .c(n_14621), .d(n_15653), .o(n_16529) );
ao12f80 g554042 ( .a(n_11806), .b(n_15200), .c(n_13209), .o(n_16301) );
in01f80 g554043 ( .a(n_17270), .o(n_16366) );
oa12f80 g554044 ( .a(n_16069), .b(n_15878), .c(n_16068), .o(n_17270) );
in01f80 g554045 ( .a(n_17005), .o(n_16365) );
oa12f80 g554046 ( .a(n_16067), .b(n_16066), .c(n_16065), .o(n_17005) );
in01f80 g554047 ( .a(n_17017), .o(n_15751) );
oa12f80 g554048 ( .a(n_15475), .b(n_15725), .c(n_15474), .o(n_17017) );
in01f80 g554049 ( .a(n_17020), .o(n_15750) );
oa12f80 g554050 ( .a(n_15473), .b(n_15721), .c(n_15472), .o(n_17020) );
in01f80 g554051 ( .a(n_17285), .o(n_16887) );
oa12f80 g554052 ( .a(n_16644), .b(n_16643), .c(n_16361), .o(n_17285) );
in01f80 g554053 ( .a(n_17288), .o(n_15749) );
oa12f80 g554054 ( .a(n_15471), .b(n_15733), .c(n_15470), .o(n_17288) );
in01f80 g554055 ( .a(n_17011), .o(n_15748) );
oa12f80 g554056 ( .a(n_15469), .b(n_15718), .c(n_15468), .o(n_17011) );
in01f80 g554057 ( .a(n_17282), .o(n_16064) );
oa12f80 g554058 ( .a(n_15747), .b(n_15746), .c(n_15730), .o(n_17282) );
in01f80 g554059 ( .a(n_17536), .o(n_15745) );
oa12f80 g554060 ( .a(n_15467), .b(n_15726), .c(n_15466), .o(n_17536) );
in01f80 g554061 ( .a(n_17279), .o(n_16063) );
oa12f80 g554062 ( .a(n_15744), .b(n_16048), .c(n_15743), .o(n_17279) );
in01f80 g554063 ( .a(n_17014), .o(n_15742) );
oa12f80 g554064 ( .a(n_15465), .b(n_15727), .c(n_15464), .o(n_17014) );
in01f80 g554065 ( .a(n_16810), .o(n_15741) );
oa12f80 g554066 ( .a(n_15463), .b(n_15679), .c(n_15462), .o(n_16810) );
in01f80 g554067 ( .a(n_17008), .o(n_16364) );
oa12f80 g554068 ( .a(n_16062), .b(n_16061), .c(n_16042), .o(n_17008) );
in01f80 g554069 ( .a(n_16807), .o(n_16060) );
oa12f80 g554070 ( .a(n_15740), .b(n_15890), .c(n_15739), .o(n_16807) );
in01f80 g554071 ( .a(n_17865), .o(n_15738) );
oa12f80 g554072 ( .a(n_14201), .b(n_15461), .c(n_14200), .o(n_17865) );
in01f80 g554073 ( .a(n_17273), .o(n_16363) );
oa12f80 g554074 ( .a(n_16059), .b(n_15989), .c(n_16058), .o(n_17273) );
in01f80 g554075 ( .a(n_17267), .o(n_16362) );
oa12f80 g554076 ( .a(n_16057), .b(n_16053), .c(n_16056), .o(n_17267) );
in01f80 g554077 ( .a(n_17276), .o(n_16055) );
oa12f80 g554078 ( .a(n_15737), .b(n_15736), .c(n_15735), .o(n_17276) );
in01f80 g554079 ( .a(n_17196), .o(n_16900) );
ao12f80 g554080 ( .a(n_15447), .b(n_15446), .c(n_15445), .o(n_17196) );
ao22s80 g554081 ( .a(n_15461), .b(n_13769), .c(n_14603), .d(x_in_56_1), .o(n_16511) );
in01f80 g554082 ( .a(n_17214), .o(n_16642) );
ao12f80 g554083 ( .a(n_15690), .b(n_16066), .c(n_15689), .o(n_17214) );
ao12f80 g554084 ( .a(n_14585), .b(n_14978), .c(n_14584), .o(n_16293) );
in01f80 g554085 ( .a(n_17213), .o(n_16641) );
ao12f80 g554086 ( .a(n_15699), .b(n_16361), .c(n_15698), .o(n_17213) );
ao12f80 g554087 ( .a(n_15713), .b(n_15712), .c(n_15711), .o(n_16360) );
oa12f80 g554088 ( .a(n_15103), .b(n_15264), .c(n_15102), .o(n_16541) );
in01f80 g554089 ( .a(n_16939), .o(n_16676) );
ao12f80 g554090 ( .a(n_15272), .b(n_15271), .c(n_15270), .o(n_16939) );
in01f80 g554091 ( .a(n_16770), .o(n_16054) );
ao12f80 g554092 ( .a(n_15175), .b(n_15878), .c(n_15377), .o(n_16770) );
in01f80 g554093 ( .a(n_16963), .o(n_16359) );
ao12f80 g554094 ( .a(n_15422), .b(n_16053), .c(n_15421), .o(n_16963) );
in01f80 g554095 ( .a(n_16769), .o(n_16052) );
ao12f80 g554096 ( .a(n_15173), .b(n_15735), .c(n_15358), .o(n_16769) );
ao12f80 g554097 ( .a(n_14968), .b(n_14967), .c(n_14966), .o(n_15460) );
in01f80 g554098 ( .a(n_17291), .o(n_16553) );
ao12f80 g554099 ( .a(n_14980), .b(n_15205), .c(n_14979), .o(n_17291) );
ao12f80 g554100 ( .a(n_15269), .b(n_15268), .c(x_in_39_13), .o(n_15734) );
ao12f80 g554101 ( .a(n_15710), .b(n_15709), .c(n_15708), .o(n_16358) );
in01f80 g554102 ( .a(n_16767), .o(n_16051) );
ao12f80 g554103 ( .a(n_15251), .b(n_15718), .c(n_15647), .o(n_16767) );
oa12f80 g554104 ( .a(n_14576), .b(n_14575), .c(n_14574), .o(n_25628) );
in01f80 g554105 ( .a(n_16766), .o(n_16050) );
ao12f80 g554106 ( .a(n_15244), .b(n_15733), .c(n_15672), .o(n_16766) );
in01f80 g554107 ( .a(n_16049), .o(n_17032) );
oa12f80 g554108 ( .a(n_15199), .b(n_15477), .c(n_15198), .o(n_16049) );
in01f80 g554109 ( .a(n_16967), .o(n_16357) );
ao12f80 g554110 ( .a(n_15411), .b(n_16048), .c(n_15694), .o(n_16967) );
ao22s80 g554111 ( .a(n_15196), .b(n_12554), .c(n_13850), .d(n_12553), .o(n_15197) );
ao22s80 g554112 ( .a(n_14976), .b(n_4044), .c(n_13388), .d(n_4043), .o(n_14977) );
oa12f80 g554113 ( .a(n_14953), .b(n_14952), .c(n_14951), .o(n_25870) );
in01f80 g554114 ( .a(n_16761), .o(n_16047) );
ao12f80 g554115 ( .a(n_15243), .b(n_15725), .c(n_15285), .o(n_16761) );
in01f80 g554116 ( .a(n_16771), .o(n_16046) );
ao12f80 g554117 ( .a(n_15178), .b(n_15989), .c(n_15428), .o(n_16771) );
in01f80 g554118 ( .a(n_16753), .o(n_17560) );
ao12f80 g554119 ( .a(n_15259), .b(n_15476), .c(n_15258), .o(n_16753) );
in01f80 g554120 ( .a(n_15731), .o(n_15732) );
oa12f80 g554121 ( .a(n_14944), .b(n_14943), .c(n_14942), .o(n_15731) );
oa12f80 g554122 ( .a(n_15266), .b(n_15265), .c(x_in_1_11), .o(n_16547) );
in01f80 g554123 ( .a(n_16768), .o(n_16045) );
ao12f80 g554124 ( .a(n_15026), .b(n_15721), .c(n_15340), .o(n_16768) );
ao22s80 g554125 ( .a(n_15194), .b(n_12958), .c(n_13851), .d(n_12957), .o(n_15195) );
ao12f80 g554126 ( .a(n_14970), .b(n_14969), .c(n_16510), .o(n_15456) );
in01f80 g554127 ( .a(n_16763), .o(n_16044) );
ao12f80 g554128 ( .a(n_15122), .b(n_15730), .c(n_15121), .o(n_16763) );
in01f80 g554129 ( .a(n_14580), .o(n_15636) );
oa12f80 g554130 ( .a(n_12861), .b(n_13489), .c(n_12860), .o(n_14580) );
oa12f80 g554131 ( .a(n_14928), .b(n_14927), .c(n_14926), .o(n_25604) );
ao22s80 g554132 ( .a(n_14974), .b(n_4075), .c(n_13387), .d(n_4074), .o(n_14975) );
oa12f80 g554133 ( .a(n_15459), .b(n_15458), .c(n_15457), .o(n_16800) );
oa12f80 g554134 ( .a(n_15668), .b(n_15667), .c(n_15997), .o(n_16734) );
ao12f80 g554135 ( .a(n_15230), .b(n_15229), .c(n_15228), .o(n_15729) );
in01f80 g554136 ( .a(n_16929), .o(n_17037) );
ao12f80 g554137 ( .a(n_15666), .b(n_15753), .c(n_15665), .o(n_16929) );
in01f80 g554138 ( .a(n_16687), .o(n_16356) );
oa12f80 g554139 ( .a(n_15297), .b(n_15296), .c(n_15295), .o(n_16687) );
ao12f80 g554140 ( .a(n_14567), .b(n_14566), .c(n_14565), .o(n_15193) );
in01f80 g554141 ( .a(n_15249), .o(n_14973) );
oa12f80 g554142 ( .a(n_13491), .b(n_14079), .c(n_13490), .o(n_15249) );
in01f80 g554143 ( .a(n_16275), .o(n_15192) );
oa12f80 g554144 ( .a(n_14078), .b(n_14581), .c(n_14077), .o(n_16275) );
oa12f80 g554145 ( .a(n_15274), .b(n_15661), .c(n_15273), .o(n_16544) );
in01f80 g554146 ( .a(n_16500), .o(n_16043) );
ao12f80 g554147 ( .a(n_15188), .b(n_15187), .c(n_15186), .o(n_16500) );
in01f80 g554148 ( .a(n_16966), .o(n_16355) );
ao12f80 g554149 ( .a(n_15349), .b(n_16042), .c(n_15696), .o(n_16966) );
in01f80 g554150 ( .a(n_17296), .o(n_15728) );
oa12f80 g554151 ( .a(n_15004), .b(n_15200), .c(n_15003), .o(n_17296) );
in01f80 g554152 ( .a(n_17499), .o(n_17171) );
ao12f80 g554153 ( .a(n_16006), .b(n_16005), .c(n_16004), .o(n_17499) );
in01f80 g554154 ( .a(n_16764), .o(n_16041) );
ao12f80 g554155 ( .a(n_15256), .b(n_15727), .c(n_15287), .o(n_16764) );
oa12f80 g554156 ( .a(n_14564), .b(n_14563), .c(n_14562), .o(n_25462) );
in01f80 g554157 ( .a(n_16765), .o(n_16040) );
ao12f80 g554158 ( .a(n_15277), .b(n_15726), .c(n_15641), .o(n_16765) );
in01f80 g554159 ( .a(n_16902), .o(n_17508) );
oa12f80 g554160 ( .a(n_16019), .b(n_16018), .c(n_16017), .o(n_16902) );
in01f80 g554161 ( .a(n_16762), .o(n_16039) );
ao12f80 g554162 ( .a(n_15022), .b(n_15679), .c(n_15662), .o(n_16762) );
ao12f80 g554163 ( .a(n_13787), .b(n_13786), .c(n_14080), .o(n_14972) );
in01f80 g554164 ( .a(n_16501), .o(n_16038) );
ao12f80 g554165 ( .a(n_15263), .b(n_15262), .c(n_15261), .o(n_16501) );
ao22s80 g554166 ( .a(n_15735), .b(n_15723), .c(n_15359), .d(x_in_58_1), .o(n_16527) );
oa22f80 g554167 ( .a(FE_OFN1029_n_14570), .b(FE_OFN412_n_28303), .c(n_641), .d(FE_OFN1111_rst), .o(n_14971) );
oa22f80 g554168 ( .a(n_13766), .b(FE_OFN204_n_28771), .c(n_1475), .d(FE_OFN1110_rst), .o(n_15191) );
oa22f80 g554169 ( .a(n_14188), .b(FE_OFN154_n_22615), .c(n_1766), .d(FE_OFN355_n_4860), .o(n_15455) );
oa22f80 g554170 ( .a(n_13764), .b(FE_OFN294_n_3069), .c(n_1346), .d(FE_OFN78_n_27012), .o(n_15190) );
oa22f80 g554171 ( .a(n_13765), .b(FE_OFN230_n_4162), .c(n_1849), .d(FE_OFN108_n_27449), .o(n_15189) );
oa22f80 g554172 ( .a(n_15014), .b(n_28303), .c(n_1116), .d(FE_OFN95_n_27449), .o(n_16037) );
oa22f80 g554173 ( .a(n_14185), .b(n_26454), .c(n_209), .d(FE_OFN68_n_27012), .o(n_15454) );
oa22f80 g554174 ( .a(n_14597), .b(FE_OFN235_n_4162), .c(n_303), .d(n_27449), .o(n_15722) );
oa22f80 g554175 ( .a(n_14127), .b(FE_OFN169_n_22948), .c(n_214), .d(FE_OFN100_n_27449), .o(n_15453) );
oa22f80 g554176 ( .a(n_14076), .b(FE_OFN249_n_4162), .c(n_798), .d(FE_OFN98_n_27449), .o(n_14579) );
ao22s80 g554177 ( .a(n_15721), .b(n_15720), .c(n_15341), .d(x_in_22_1), .o(n_16525) );
oa22f80 g554178 ( .a(n_14126), .b(FE_OFN171_n_22948), .c(n_1143), .d(FE_OFN1112_rst), .o(n_15452) );
oa22f80 g554179 ( .a(FE_OFN859_n_14125), .b(n_21076), .c(n_676), .d(FE_OFN324_n_4860), .o(n_15451) );
oa22f80 g554180 ( .a(n_14124), .b(FE_OFN234_n_4162), .c(n_930), .d(FE_OFN1182_rst), .o(n_15450) );
ao22s80 g554181 ( .a(n_16066), .b(n_16026), .c(n_15430), .d(x_in_2_1), .o(n_16714) );
oa22f80 g554182 ( .a(n_16035), .b(FE_OFN265_n_4280), .c(n_374), .d(FE_OFN1146_n_4860), .o(n_16036) );
oa22f80 g554183 ( .a(n_14123), .b(n_4280), .c(n_1013), .d(n_27449), .o(n_15449) );
ao22s80 g554184 ( .a(n_15718), .b(n_15717), .c(n_15648), .d(x_in_54_1), .o(n_16502) );
oa22f80 g554185 ( .a(n_14131), .b(FE_OFN256_n_4280), .c(n_834), .d(FE_OFN1123_rst), .o(n_15448) );
oa22f80 g554186 ( .a(n_12859), .b(FE_OFN267_n_4280), .c(n_1656), .d(FE_OFN92_n_27449), .o(n_14577) );
ao22s80 g554187 ( .a(n_15725), .b(n_15724), .c(n_15286), .d(x_in_14_1), .o(n_16523) );
ao22s80 g554188 ( .a(n_15733), .b(n_15810), .c(n_15673), .d(x_in_46_1), .o(n_16521) );
ao22s80 g554189 ( .a(n_16361), .b(n_16351), .c(n_15352), .d(x_in_34_1), .o(n_16712) );
ao22s80 g554190 ( .a(n_15730), .b(n_15444), .c(n_14935), .d(x_in_16_1), .o(n_16273) );
oa22f80 g554191 ( .a(n_16008), .b(FE_OFN253_n_4280), .c(n_1633), .d(FE_OFN141_n_27449), .o(n_16009) );
oa22f80 g554192 ( .a(n_15715), .b(FE_OFN223_n_21642), .c(n_1593), .d(FE_OFN1112_rst), .o(n_15716) );
ao22s80 g554193 ( .a(n_15726), .b(n_16013), .c(n_15642), .d(x_in_30_1), .o(n_16519) );
ao22s80 g554194 ( .a(n_15727), .b(n_16012), .c(n_15288), .d(x_in_62_1), .o(n_16517) );
ao22s80 g554195 ( .a(n_16048), .b(n_16354), .c(n_15695), .d(x_in_18_1), .o(n_16710) );
oa22f80 g554196 ( .a(n_13367), .b(FE_OFN234_n_4162), .c(n_150), .d(FE_OFN76_n_27012), .o(n_14591) );
ao22s80 g554197 ( .a(n_15679), .b(n_15678), .c(n_15663), .d(x_in_12_1), .o(n_16515) );
oa22f80 g554198 ( .a(n_13761), .b(FE_OFN310_n_3069), .c(n_117), .d(FE_OFN129_n_27449), .o(n_13762) );
oa22f80 g554199 ( .a(n_12857), .b(FE_OFN234_n_4162), .c(n_810), .d(FE_OFN360_n_4860), .o(n_14426) );
ao22s80 g554200 ( .a(n_16042), .b(n_16031), .c(n_15697), .d(x_in_50_1), .o(n_16708) );
oa22f80 g554201 ( .a(n_14176), .b(n_21988), .c(n_703), .d(FE_OFN324_n_4860), .o(n_15664) );
oa22f80 g554202 ( .a(n_15890), .b(FE_OFN1176_n_28597), .c(n_253), .d(FE_OFN1111_rst), .o(n_15719) );
ao22s80 g554203 ( .a(n_15878), .b(n_15877), .c(n_15378), .d(x_in_42_1), .o(n_16506) );
ao22s80 g554204 ( .a(n_15989), .b(n_15988), .c(n_15429), .d(x_in_10_1), .o(n_16508) );
oa22f80 g554205 ( .a(FE_OFN460_n_13371), .b(FE_OFN257_n_4280), .c(n_950), .d(FE_OFN190_n_28362), .o(n_14993) );
ao22s80 g554206 ( .a(n_16053), .b(n_16007), .c(n_15171), .d(x_in_26_1), .o(n_16504) );
oa22f80 g554207 ( .a(FE_OFN534_n_13775), .b(FE_OFN266_n_4280), .c(n_1909), .d(n_25680), .o(n_15276) );
oa22f80 g554208 ( .a(n_14122), .b(FE_OFN230_n_4162), .c(n_1807), .d(FE_OFN21_n_27452), .o(n_15669) );
oa22f80 g554209 ( .a(FE_OFN895_n_15923), .b(FE_OFN240_n_4162), .c(n_1062), .d(FE_OFN1121_rst), .o(n_14665) );
ao12f80 g554210 ( .a(n_15006), .b(x_out_53_29), .c(n_17184), .o(n_15281) );
ao22s80 g554211 ( .a(n_15059), .b(n_4882), .c(x_out_54_29), .d(FE_OFN271_n_16028), .o(n_15289) );
ao22s80 g554212 ( .a(n_15996), .b(n_4193), .c(x_out_60_29), .d(FE_OFN273_n_16893), .o(n_16027) );
ao22s80 g554213 ( .a(n_15999), .b(n_4195), .c(x_out_61_29), .d(FE_OFN271_n_16028), .o(n_16029) );
ao22s80 g554214 ( .a(n_16023), .b(n_4316), .c(x_out_63_29), .d(FE_OFN196_n_5003), .o(n_16030) );
oa22f80 g554215 ( .a(FE_OFN690_n_16216), .b(FE_OFN402_n_28303), .c(n_127), .d(FE_OFN122_n_27449), .o(n_15182) );
ao22s80 g554216 ( .a(n_15890), .b(n_15992), .c(n_15889), .d(x_in_44_1), .o(n_16513) );
ao22s80 g554218 ( .a(n_15890), .b(n_15247), .c(n_15889), .d(n_11641), .o(n_16760) );
ao22s80 g554219 ( .a(n_14478), .b(x_in_7_13), .c(n_14594), .d(n_7285), .o(n_15639) );
ao22s80 g554220 ( .a(n_15035), .b(x_in_23_13), .c(n_15670), .d(n_6488), .o(n_16349) );
ao22s80 g554221 ( .a(n_15034), .b(x_in_31_13), .c(n_15280), .d(n_7291), .o(n_16352) );
ao22s80 g554222 ( .a(n_15036), .b(x_in_55_13), .c(n_15671), .d(n_7231), .o(n_16353) );
no02f80 g554270 ( .a(n_15268), .b(x_in_39_13), .o(n_15269) );
na02f80 g554271 ( .a(n_14079), .b(n_13490), .o(n_13491) );
in01f80 g554272 ( .a(n_15001), .o(n_15002) );
na02f80 g554273 ( .a(n_14589), .b(FE_OFN1174_n_4860), .o(n_15001) );
in01f80 g554274 ( .a(n_14999), .o(n_15000) );
na02f80 g554275 ( .a(n_14588), .b(FE_OFN34_n_15183), .o(n_14999) );
na02f80 g554276 ( .a(n_16011), .b(n_16010), .o(n_16021) );
no02f80 g554277 ( .a(n_14589), .b(n_13677), .o(n_15915) );
na02f80 g554278 ( .a(n_15998), .b(x_in_8_3), .o(n_16653) );
in01f80 g554279 ( .a(n_18822), .o(n_16392) );
na02f80 g554280 ( .a(n_16675), .b(x_in_6_0), .o(n_18822) );
in01f80 g554281 ( .a(n_16024), .o(n_16025) );
no02f80 g554282 ( .a(n_15998), .b(x_in_8_3), .o(n_16024) );
na02f80 g554283 ( .a(n_15268), .b(n_7213), .o(n_15922) );
na02f80 g554284 ( .a(n_15016), .b(n_784), .o(n_15677) );
in01f80 g554285 ( .a(n_18209), .o(n_16134) );
na02f80 g554286 ( .a(n_15769), .b(x_in_52_0), .o(n_18209) );
na02f80 g554287 ( .a(n_14616), .b(n_119), .o(n_15292) );
no02f80 g554288 ( .a(n_15271), .b(n_15270), .o(n_15272) );
na02f80 g554289 ( .a(n_15296), .b(n_15295), .o(n_15297) );
in01f80 g554290 ( .a(n_15338), .o(n_15339) );
na02f80 g554291 ( .a(n_15108), .b(n_14501), .o(n_15338) );
na03f80 g554292 ( .a(n_13753), .b(n_18116), .c(FE_OFN422_n_16909), .o(n_15554) );
no02f80 g554293 ( .a(n_15205), .b(n_14979), .o(n_14980) );
na02f80 g554294 ( .a(n_15660), .b(x_in_24_3), .o(n_16424) );
na02f80 g554295 ( .a(n_15434), .b(n_15638), .o(n_16217) );
na03f80 g554296 ( .a(n_15010), .b(n_18113), .c(FE_OFN421_n_16909), .o(n_16372) );
na03f80 g554297 ( .a(n_13750), .b(n_17645), .c(FE_OFN385_n_16289), .o(n_15534) );
na03f80 g554298 ( .a(n_13328), .b(n_17882), .c(n_16289), .o(n_15213) );
in01f80 g554299 ( .a(n_15994), .o(n_15995) );
na02f80 g554300 ( .a(n_14839), .b(n_15655), .o(n_15994) );
na02f80 g554301 ( .a(n_15267), .b(x_in_0_9), .o(n_16188) );
in01f80 g554302 ( .a(n_15658), .o(n_15659) );
no02f80 g554303 ( .a(n_15267), .b(x_in_0_9), .o(n_15658) );
in01f80 g554304 ( .a(n_15675), .o(n_15676) );
na02f80 g554305 ( .a(n_15275), .b(n_14506), .o(n_15675) );
na03f80 g554306 ( .a(n_14111), .b(n_17874), .c(FE_OFN382_n_16289), .o(n_15817) );
no02f80 g554307 ( .a(n_16003), .b(n_16002), .o(n_16416) );
in01f80 g554308 ( .a(n_16389), .o(n_19129) );
no02f80 g554309 ( .a(n_16011), .b(n_16010), .o(n_16389) );
in01f80 g554310 ( .a(n_18203), .o(n_16391) );
na02f80 g554311 ( .a(n_15807), .b(x_in_48_0), .o(n_18203) );
na02f80 g554312 ( .a(n_15017), .b(n_1810), .o(n_16022) );
na02f80 g554313 ( .a(n_15008), .b(n_15007), .o(n_15924) );
na02f80 g554314 ( .a(n_15282), .b(x_in_8_2), .o(n_16414) );
in01f80 g554315 ( .a(n_15680), .o(n_15681) );
no02f80 g554316 ( .a(n_15282), .b(x_in_8_2), .o(n_15680) );
in01f80 g554317 ( .a(n_18206), .o(n_16133) );
na02f80 g554318 ( .a(n_15819), .b(x_in_32_0), .o(n_18206) );
in01f80 g554319 ( .a(n_19414), .o(n_16650) );
na02f80 g554320 ( .a(n_17170), .b(x_in_20_0), .o(n_19414) );
na02f80 g554321 ( .a(n_14611), .b(n_1705), .o(n_15346) );
na02f80 g554322 ( .a(n_15283), .b(n_1599), .o(n_16034) );
in01f80 g554323 ( .a(n_18458), .o(n_16390) );
na02f80 g554324 ( .a(n_16105), .b(x_in_40_0), .o(n_18458) );
na02f80 g554325 ( .a(n_15020), .b(n_1790), .o(n_15714) );
na02f80 g554326 ( .a(n_14581), .b(n_14077), .o(n_14078) );
na02f80 g554327 ( .a(n_13761), .b(n_14080), .o(n_15254) );
na03f80 g554328 ( .a(n_13741), .b(n_17666), .c(FE_OFN383_n_16289), .o(n_16082) );
na03f80 g554329 ( .a(n_14110), .b(n_17674), .c(FE_OFN421_n_16909), .o(n_15790) );
in01f80 g554330 ( .a(n_15656), .o(n_15657) );
no02f80 g554331 ( .a(n_15264), .b(x_in_56_2), .o(n_15656) );
na03f80 g554332 ( .a(n_14109), .b(n_17671), .c(FE_OFN382_n_16289), .o(n_15853) );
na02f80 g554333 ( .a(n_14996), .b(x_in_4_9), .o(n_15899) );
in01f80 g554334 ( .a(n_15278), .o(n_15279) );
no02f80 g554335 ( .a(n_14996), .b(x_in_4_9), .o(n_15278) );
no02f80 g554336 ( .a(n_16001), .b(FE_OFN600_n_16000), .o(n_16426) );
no02f80 g554337 ( .a(n_16005), .b(n_16004), .o(n_16006) );
in01f80 g554338 ( .a(n_19737), .o(n_16388) );
na02f80 g554339 ( .a(n_17172), .b(x_in_36_0), .o(n_19737) );
na02f80 g554340 ( .a(n_15019), .b(n_1914), .o(n_16015) );
na02f80 g554341 ( .a(n_16018), .b(n_16017), .o(n_16019) );
na03f80 g554342 ( .a(n_14108), .b(n_17877), .c(FE_OFN1109_rst), .o(n_15773) );
no02f80 g554343 ( .a(n_14588), .b(n_13675), .o(n_15896) );
no02f80 g554344 ( .a(n_13786), .b(n_14080), .o(n_13787) );
in01f80 g554345 ( .a(n_15683), .o(n_15684) );
no02f80 g554346 ( .a(n_15660), .b(x_in_24_3), .o(n_15683) );
na02f80 g554347 ( .a(n_15264), .b(x_in_56_2), .o(n_16215) );
na02f80 g554348 ( .a(n_13489), .b(n_12860), .o(n_12861) );
no02f80 g554349 ( .a(n_14496), .b(x_in_1_11), .o(n_15620) );
no02f80 g554350 ( .a(n_15446), .b(n_15445), .o(n_15447) );
na02f80 g554351 ( .a(n_15458), .b(n_15457), .o(n_15459) );
no02f80 g554352 ( .a(n_15242), .b(n_10075), .o(n_15886) );
no02f80 g554353 ( .a(n_14620), .b(n_4972), .o(n_15674) );
no02f80 g554354 ( .a(n_14978), .b(n_14584), .o(n_14585) );
na02f80 g554355 ( .a(n_14991), .b(n_14460), .o(n_15592) );
no02f80 g554356 ( .a(n_15476), .b(n_15258), .o(n_15259) );
no02f80 g554357 ( .a(n_15654), .b(n_15653), .o(n_16466) );
na02f80 g554358 ( .a(n_15996), .b(n_3872), .o(n_16397) );
na02f80 g554359 ( .a(n_15999), .b(n_3870), .o(n_16401) );
na02f80 g554360 ( .a(n_16023), .b(n_3504), .o(n_16399) );
no02f80 g554361 ( .a(n_15645), .b(x_in_63_13), .o(n_16164) );
no02f80 g554362 ( .a(n_15643), .b(x_in_15_13), .o(n_16166) );
no02f80 g554363 ( .a(n_15649), .b(x_in_47_13), .o(n_16162) );
in01f80 g554364 ( .a(n_16159), .o(n_16016) );
no02f80 g554365 ( .a(n_15670), .b(x_in_23_13), .o(n_16159) );
in01f80 g554366 ( .a(n_16157), .o(n_16014) );
no02f80 g554367 ( .a(n_15671), .b(x_in_55_13), .o(n_16157) );
in01f80 g554368 ( .a(n_16155), .o(n_16020) );
no02f80 g554369 ( .a(n_15280), .b(x_in_31_13), .o(n_16155) );
in01f80 g554370 ( .a(n_15591), .o(n_15009) );
no02f80 g554371 ( .a(n_14594), .b(x_in_7_13), .o(n_15591) );
no02f80 g554372 ( .a(n_15187), .b(n_15186), .o(n_15188) );
no02f80 g554373 ( .a(n_14480), .b(n_14481), .o(n_25173) );
na02f80 g554374 ( .a(n_15185), .b(n_15184), .o(n_15875) );
no02f80 g554375 ( .a(n_15288), .b(n_15287), .o(n_16143) );
no02f80 g554376 ( .a(n_15341), .b(n_15340), .o(n_16152) );
no02f80 g554377 ( .a(n_15721), .b(n_15340), .o(n_15026) );
no02f80 g554378 ( .a(n_15663), .b(n_15662), .o(n_16138) );
no02f80 g554379 ( .a(n_15725), .b(n_15285), .o(n_15243) );
no02f80 g554380 ( .a(n_15733), .b(n_15672), .o(n_15244) );
no02f80 g554381 ( .a(n_15642), .b(n_15641), .o(n_16393) );
no02f80 g554382 ( .a(n_15727), .b(n_15287), .o(n_15256) );
na02f80 g554383 ( .a(n_14058), .b(n_14992), .o(n_15575) );
no02f80 g554384 ( .a(n_15648), .b(n_15647), .o(n_16140) );
na02f80 g554385 ( .a(n_15265), .b(x_in_1_11), .o(n_15266) );
no02f80 g554386 ( .a(n_15998), .b(n_15997), .o(n_16395) );
na02f80 g554387 ( .a(n_15667), .b(n_15997), .o(n_15668) );
no02f80 g554388 ( .a(n_15661), .b(n_15660), .o(n_16277) );
na02f80 g554389 ( .a(n_15661), .b(n_15273), .o(n_15274) );
no02f80 g554390 ( .a(n_15726), .b(n_15641), .o(n_15277) );
no02f80 g554391 ( .a(n_15673), .b(n_15672), .o(n_16147) );
no02f80 g554392 ( .a(n_15718), .b(n_15647), .o(n_15251) );
no02f80 g554393 ( .a(n_15679), .b(n_15662), .o(n_15022) );
no02f80 g554394 ( .a(n_15286), .b(n_15285), .o(n_16150) );
in01f80 g554395 ( .a(n_15293), .o(n_15294) );
na02f80 g554396 ( .a(n_15059), .b(n_14997), .o(n_15293) );
no02f80 g554397 ( .a(n_15889), .b(n_15247), .o(n_15874) );
no02f80 g554398 ( .a(n_14969), .b(n_16510), .o(n_14970) );
no02f80 g554399 ( .a(n_15229), .b(n_15228), .o(n_15230) );
no02f80 g554400 ( .a(n_15005), .b(n_8188), .o(n_15006) );
na02f80 g554401 ( .a(n_15643), .b(n_2575), .o(n_15644) );
na02f80 g554402 ( .a(n_15645), .b(n_2523), .o(n_15646) );
na02f80 g554403 ( .a(n_15649), .b(n_2448), .o(n_15650) );
no02f80 g554404 ( .a(n_15262), .b(n_15261), .o(n_15263) );
in01f80 g554405 ( .a(n_14994), .o(n_14995) );
na02f80 g554406 ( .a(n_14587), .b(n_4860), .o(n_14994) );
na02f80 g554407 ( .a(n_13378), .b(n_14081), .o(n_15579) );
na02f80 g554408 ( .a(n_14472), .b(n_14997), .o(n_14998) );
no02f80 g554409 ( .a(n_15753), .b(n_15665), .o(n_15666) );
na02f80 g554410 ( .a(n_15200), .b(n_15003), .o(n_15004) );
oa22f80 g554411 ( .a(n_12824), .b(n_8803), .c(n_3656), .d(x_in_61_14), .o(n_14082) );
no02f80 g554412 ( .a(n_15712), .b(n_15711), .o(n_15713) );
no02f80 g554413 ( .a(n_15709), .b(n_15708), .o(n_15710) );
na02f80 g554414 ( .a(n_15477), .b(n_15198), .o(n_15199) );
no02f80 g554415 ( .a(n_14459), .b(n_15011), .o(n_16588) );
in01f80 g554416 ( .a(n_15442), .o(n_15443) );
na02f80 g554417 ( .a(n_15242), .b(FE_OFN34_n_15183), .o(n_15442) );
in01f80 g554418 ( .a(n_15755), .o(n_15441) );
na02f80 g554419 ( .a(n_16686), .b(rst), .o(n_15755) );
in01f80 g554420 ( .a(n_15439), .o(n_15440) );
no02f80 g554421 ( .a(n_15185), .b(n_2022), .o(n_15439) );
in01f80 g554422 ( .a(n_16033), .o(n_16645) );
no02f80 g554423 ( .a(n_15707), .b(n_2022), .o(n_16033) );
na02f80 g554424 ( .a(n_16003), .b(FE_OFN350_n_4860), .o(n_16370) );
na02f80 g554425 ( .a(n_16001), .b(FE_OFN1174_n_4860), .o(n_16368) );
in01f80 g554426 ( .a(n_15437), .o(n_15438) );
no02f80 g554427 ( .a(n_15008), .b(FE_OFN413_n_28303), .o(n_15437) );
in01f80 g554428 ( .a(n_15705), .o(n_15706) );
na02f80 g554429 ( .a(n_15436), .b(FE_OFN1154_n_14586), .o(n_15705) );
in01f80 g554430 ( .a(n_15703), .o(n_15704) );
na02f80 g554431 ( .a(n_15435), .b(FE_OFN1113_rst), .o(n_15703) );
in01f80 g554432 ( .a(n_15701), .o(n_15702) );
no02f80 g554433 ( .a(n_15434), .b(n_2022), .o(n_15701) );
no02f80 g554434 ( .a(n_14799), .b(n_15433), .o(n_16600) );
na02f80 g554435 ( .a(n_16234), .b(n_14919), .o(n_15891) );
na02f80 g554436 ( .a(n_14761), .b(n_15432), .o(n_16339) );
no02f80 g554437 ( .a(n_14202), .b(n_11038), .o(n_15571) );
na02f80 g554438 ( .a(n_14769), .b(n_15431), .o(n_21972) );
no02f80 g554439 ( .a(n_14967), .b(n_14966), .o(n_14968) );
in01f80 g554440 ( .a(n_16084), .o(n_15700) );
no02f80 g554441 ( .a(n_15430), .b(n_15689), .o(n_16084) );
no02f80 g554442 ( .a(n_15429), .b(n_15428), .o(n_16124) );
na02f80 g554443 ( .a(n_14177), .b(n_13589), .o(n_25728) );
in01f80 g554444 ( .a(n_15180), .o(n_15181) );
na02f80 g554445 ( .a(n_14191), .b(n_14189), .o(n_15180) );
in01f80 g554446 ( .a(n_17181), .o(n_15427) );
oa12f80 g554447 ( .a(n_15039), .b(n_14120), .c(n_11750), .o(n_17181) );
na02f80 g554448 ( .a(n_14192), .b(n_14190), .o(n_15861) );
no02f80 g554449 ( .a(n_16361), .b(n_15698), .o(n_15699) );
no02f80 g554450 ( .a(n_14783), .b(n_15426), .o(n_17156) );
na02f80 g554451 ( .a(n_15177), .b(n_15176), .o(n_16121) );
na02f80 g554452 ( .a(n_14964), .b(n_15948), .o(n_14965) );
na02f80 g554453 ( .a(n_14256), .b(n_15179), .o(n_19033) );
na02f80 g554454 ( .a(n_15950), .b(n_14964), .o(n_15618) );
no02f80 g554455 ( .a(n_15989), .b(n_15428), .o(n_15178) );
no02f80 g554456 ( .a(n_13827), .b(n_11729), .o(n_14963) );
no02f80 g554457 ( .a(n_13826), .b(n_11728), .o(n_14578) );
in01f80 g554458 ( .a(n_15424), .o(n_15425) );
no02f80 g554459 ( .a(n_15177), .b(n_15176), .o(n_15424) );
no02f80 g554460 ( .a(n_15878), .b(n_15377), .o(n_15175) );
na02f80 g554461 ( .a(n_14193), .b(n_11737), .o(n_15850) );
na02f80 g554462 ( .a(n_14194), .b(n_11738), .o(n_15849) );
na02f80 g554463 ( .a(n_14755), .b(n_15423), .o(n_18085) );
na02f80 g554464 ( .a(n_14962), .b(n_14007), .o(n_15614) );
no02f80 g554465 ( .a(n_16053), .b(n_15421), .o(n_15422) );
na02f80 g554466 ( .a(n_14404), .b(n_15174), .o(n_24896) );
in01f80 g554467 ( .a(n_15419), .o(n_15420) );
no02f80 g554468 ( .a(n_14180), .b(n_9682), .o(n_15419) );
no02f80 g554469 ( .a(n_15735), .b(n_15358), .o(n_15173) );
na02f80 g554470 ( .a(n_14233), .b(n_15172), .o(n_17126) );
no02f80 g554471 ( .a(n_14763), .b(n_15418), .o(n_19057) );
in01f80 g554472 ( .a(n_15845), .o(n_15417) );
no02f80 g554473 ( .a(n_15171), .b(n_15421), .o(n_15845) );
no02f80 g554474 ( .a(n_14445), .b(n_15170), .o(n_20848) );
na02f80 g554475 ( .a(n_13996), .b(n_14961), .o(n_19694) );
no02f80 g554476 ( .a(n_14313), .b(n_15169), .o(n_15881) );
no02f80 g554477 ( .a(n_14779), .b(n_15416), .o(n_21163) );
na02f80 g554478 ( .a(n_15415), .b(n_14637), .o(n_20078) );
no02f80 g554479 ( .a(n_14777), .b(n_15414), .o(n_19359) );
no02f80 g554480 ( .a(n_14773), .b(n_15413), .o(n_16185) );
in01f80 g554481 ( .a(n_15167), .o(n_15168) );
no02f80 g554482 ( .a(n_14183), .b(n_12419), .o(n_15167) );
in01f80 g554483 ( .a(n_14959), .o(n_14960) );
na02f80 g554484 ( .a(n_13807), .b(n_11067), .o(n_14959) );
in01f80 g554485 ( .a(n_15165), .o(n_15166) );
na02f80 g554486 ( .a(n_14181), .b(n_9713), .o(n_15165) );
na02f80 g554487 ( .a(n_13998), .b(n_14958), .o(n_21952) );
na02f80 g554488 ( .a(n_15412), .b(n_14766), .o(n_19714) );
na02f80 g554489 ( .a(n_14182), .b(n_9714), .o(n_15844) );
na02f80 g554490 ( .a(n_14575), .b(n_14574), .o(n_14576) );
na02f80 g554491 ( .a(n_14437), .b(n_15164), .o(n_16317) );
in01f80 g554492 ( .a(n_15162), .o(n_15163) );
no02f80 g554493 ( .a(n_14140), .b(n_12400), .o(n_15162) );
no02f80 g554494 ( .a(n_14141), .b(n_12401), .o(n_15839) );
no02f80 g554495 ( .a(n_16048), .b(n_15694), .o(n_15411) );
in01f80 g554496 ( .a(n_14956), .o(n_14957) );
na02f80 g554497 ( .a(n_13805), .b(n_11065), .o(n_14956) );
no02f80 g554498 ( .a(n_14443), .b(n_15161), .o(n_19035) );
no02f80 g554499 ( .a(n_14767), .b(n_15410), .o(n_20868) );
na02f80 g554500 ( .a(n_14424), .b(n_15160), .o(n_22234) );
no02f80 g554501 ( .a(n_14751), .b(n_15409), .o(n_20866) );
na02f80 g554502 ( .a(n_15408), .b(n_14796), .o(n_19712) );
no02f80 g554503 ( .a(n_14753), .b(n_15407), .o(n_19055) );
na02f80 g554504 ( .a(n_14652), .b(n_15406), .o(n_18081) );
no02f80 g554505 ( .a(n_14756), .b(n_15405), .o(n_17152) );
na02f80 g554506 ( .a(n_15404), .b(n_14642), .o(n_16337) );
no02f80 g554507 ( .a(n_14668), .b(n_15403), .o(n_16207) );
in01f80 g554508 ( .a(n_15158), .o(n_15159) );
no02f80 g554509 ( .a(n_14172), .b(n_12398), .o(n_15158) );
no02f80 g554510 ( .a(n_14173), .b(n_12399), .o(n_15836) );
in01f80 g554511 ( .a(n_14954), .o(n_14955) );
na02f80 g554512 ( .a(n_13803), .b(n_11063), .o(n_14954) );
na02f80 g554513 ( .a(n_13804), .b(n_11062), .o(n_15544) );
in01f80 g554514 ( .a(n_15401), .o(n_15402) );
no02f80 g554515 ( .a(n_14171), .b(n_9667), .o(n_15401) );
no02f80 g554516 ( .a(n_14170), .b(n_9668), .o(n_15835) );
no02f80 g554517 ( .a(n_14421), .b(n_15157), .o(n_21146) );
na02f80 g554518 ( .a(n_14418), .b(n_15156), .o(n_20067) );
no02f80 g554519 ( .a(n_14416), .b(n_15155), .o(n_19346) );
na02f80 g554520 ( .a(n_15400), .b(n_14747), .o(n_21970) );
na02f80 g554521 ( .a(n_14414), .b(n_15154), .o(n_18350) );
no02f80 g554522 ( .a(n_14410), .b(n_15153), .o(n_17448) );
na02f80 g554523 ( .a(n_14408), .b(n_15152), .o(n_16586) );
no02f80 g554524 ( .a(n_14406), .b(n_15151), .o(n_15879) );
no02f80 g554525 ( .a(n_14394), .b(n_15150), .o(n_23197) );
in01f80 g554526 ( .a(n_15148), .o(n_15149) );
na02f80 g554527 ( .a(n_14168), .b(n_10575), .o(n_15148) );
na02f80 g554528 ( .a(n_14169), .b(n_10574), .o(n_15832) );
no02f80 g554529 ( .a(n_14744), .b(n_15399), .o(n_20864) );
na02f80 g554530 ( .a(n_15398), .b(n_14743), .o(n_19710) );
no02f80 g554531 ( .a(n_14740), .b(n_15397), .o(n_19053) );
na02f80 g554532 ( .a(n_14738), .b(n_15396), .o(n_18079) );
no02f80 g554533 ( .a(n_14736), .b(n_15395), .o(n_17150) );
na02f80 g554534 ( .a(n_15394), .b(n_14734), .o(n_16335) );
no02f80 g554535 ( .a(n_14733), .b(n_15393), .o(n_16202) );
in01f80 g554536 ( .a(n_15146), .o(n_15147) );
no02f80 g554537 ( .a(n_14166), .b(n_12388), .o(n_15146) );
na02f80 g554538 ( .a(n_14952), .b(n_14951), .o(n_14953) );
no02f80 g554539 ( .a(n_14167), .b(n_12389), .o(n_15829) );
in01f80 g554540 ( .a(n_14949), .o(n_14950) );
na02f80 g554541 ( .a(n_13801), .b(n_11061), .o(n_14949) );
na02f80 g554542 ( .a(n_13802), .b(n_11060), .o(n_15543) );
in01f80 g554543 ( .a(n_15391), .o(n_15392) );
no02f80 g554544 ( .a(n_14165), .b(n_9658), .o(n_15391) );
no02f80 g554545 ( .a(n_14164), .b(n_9659), .o(n_15828) );
no02f80 g554546 ( .a(n_15145), .b(n_14386), .o(n_21968) );
oa12f80 g554547 ( .a(n_12074), .b(n_14515), .c(n_13236), .o(n_15909) );
na02f80 g554548 ( .a(n_14383), .b(n_15144), .o(n_20862) );
no02f80 g554549 ( .a(n_14381), .b(n_15143), .o(n_19708) );
na02f80 g554550 ( .a(n_14379), .b(n_15142), .o(n_19051) );
no02f80 g554551 ( .a(n_14377), .b(n_15141), .o(n_18077) );
na02f80 g554552 ( .a(n_14375), .b(n_15140), .o(n_17148) );
no02f80 g554553 ( .a(n_15139), .b(n_14373), .o(n_16333) );
na02f80 g554554 ( .a(n_14371), .b(n_15138), .o(n_15908) );
na02f80 g554555 ( .a(n_14730), .b(n_15390), .o(n_22918) );
na02f80 g554556 ( .a(n_14883), .b(n_15137), .o(n_25452) );
no02f80 g554557 ( .a(n_15389), .b(n_14725), .o(n_22238) );
no02f80 g554558 ( .a(n_14359), .b(n_15136), .o(n_21956) );
na02f80 g554559 ( .a(n_15388), .b(n_14719), .o(n_21966) );
no02f80 g554560 ( .a(n_14716), .b(n_15387), .o(n_20860) );
na02f80 g554561 ( .a(n_15386), .b(n_14714), .o(n_19706) );
no02f80 g554562 ( .a(n_14712), .b(n_15385), .o(n_19049) );
na02f80 g554563 ( .a(n_14710), .b(n_15384), .o(n_18075) );
no02f80 g554564 ( .a(n_14708), .b(n_15383), .o(n_17146) );
na02f80 g554565 ( .a(n_14704), .b(n_15382), .o(n_16331) );
no02f80 g554566 ( .a(n_14701), .b(n_15381), .o(n_16195) );
in01f80 g554567 ( .a(n_15134), .o(n_15135) );
no02f80 g554568 ( .a(n_14160), .b(n_12920), .o(n_15134) );
na02f80 g554569 ( .a(n_14352), .b(n_15133), .o(n_20852) );
no02f80 g554570 ( .a(n_14161), .b(n_12921), .o(n_15826) );
no02f80 g554571 ( .a(n_14350), .b(n_15132), .o(n_19698) );
na02f80 g554572 ( .a(n_14346), .b(n_15131), .o(n_19039) );
in01f80 g554573 ( .a(n_14947), .o(n_14948) );
na02f80 g554574 ( .a(n_13799), .b(n_11059), .o(n_14947) );
no02f80 g554575 ( .a(n_14344), .b(n_15130), .o(n_18067) );
na02f80 g554576 ( .a(n_13800), .b(n_11058), .o(n_15541) );
na02f80 g554577 ( .a(n_14342), .b(n_15129), .o(n_17138) );
no02f80 g554578 ( .a(n_13971), .b(n_14946), .o(n_16321) );
in01f80 g554579 ( .a(n_15379), .o(n_15380) );
no02f80 g554580 ( .a(n_14159), .b(n_9628), .o(n_15379) );
no02f80 g554581 ( .a(n_14158), .b(n_9629), .o(n_15825) );
na02f80 g554582 ( .a(n_13968), .b(n_14945), .o(n_22907) );
no02f80 g554583 ( .a(n_15378), .b(n_15377), .o(n_16120) );
in01f80 g554584 ( .a(n_15127), .o(n_15128) );
no02f80 g554585 ( .a(n_14156), .b(n_9765), .o(n_15127) );
na02f80 g554586 ( .a(n_15376), .b(n_14693), .o(n_21964) );
no02f80 g554587 ( .a(n_14157), .b(n_9764), .o(n_15824) );
na02f80 g554588 ( .a(n_14943), .b(n_14942), .o(n_14944) );
na02f80 g554589 ( .a(n_14722), .b(n_15375), .o(n_21152) );
no02f80 g554590 ( .a(n_14643), .b(n_15374), .o(n_16171) );
no02f80 g554591 ( .a(n_15373), .b(n_14703), .o(n_20073) );
na02f80 g554592 ( .a(n_14706), .b(n_15372), .o(n_19352) );
no02f80 g554593 ( .a(n_14698), .b(n_15371), .o(n_18356) );
na02f80 g554594 ( .a(n_14696), .b(n_15370), .o(n_17454) );
no02f80 g554595 ( .a(n_14690), .b(n_15369), .o(n_20858) );
na02f80 g554596 ( .a(n_15368), .b(n_14689), .o(n_19704) );
na02f80 g554597 ( .a(n_13880), .b(n_14941), .o(n_19027) );
no02f80 g554598 ( .a(n_14686), .b(n_15367), .o(n_19047) );
na02f80 g554599 ( .a(n_14684), .b(n_15366), .o(n_18073) );
no02f80 g554600 ( .a(n_14682), .b(n_15365), .o(n_17144) );
na02f80 g554601 ( .a(n_14680), .b(n_15364), .o(n_16329) );
no02f80 g554602 ( .a(n_14679), .b(n_15363), .o(n_16189) );
in01f80 g554603 ( .a(n_15125), .o(n_15126) );
no02f80 g554604 ( .a(n_14154), .b(n_12910), .o(n_15125) );
no02f80 g554605 ( .a(n_14155), .b(n_12911), .o(n_15823) );
in01f80 g554606 ( .a(n_14939), .o(n_14940) );
na02f80 g554607 ( .a(n_13796), .b(n_11057), .o(n_14939) );
na02f80 g554608 ( .a(n_13797), .b(n_11056), .o(n_15537) );
in01f80 g554609 ( .a(n_15361), .o(n_15362) );
no02f80 g554610 ( .a(n_14153), .b(n_9624), .o(n_15361) );
na02f80 g554611 ( .a(n_14676), .b(n_15360), .o(n_23201) );
no02f80 g554612 ( .a(n_14152), .b(n_9625), .o(n_15822) );
no02f80 g554613 ( .a(n_15697), .b(n_15696), .o(n_16381) );
no02f80 g554614 ( .a(n_15359), .b(n_15358), .o(n_16116) );
in01f80 g554615 ( .a(n_14937), .o(n_14938) );
na02f80 g554616 ( .a(n_14569), .b(n_14568), .o(n_14937) );
na02f80 g554617 ( .a(n_13963), .b(n_14936), .o(n_21942) );
na02f80 g554618 ( .a(n_14608), .b(n_15124), .o(n_15815) );
in01f80 g554619 ( .a(n_15813), .o(n_15123) );
no02f80 g554620 ( .a(n_14935), .b(n_15121), .o(n_15813) );
no02f80 g554621 ( .a(n_15730), .b(n_15121), .o(n_15122) );
in01f80 g554622 ( .a(n_15356), .o(n_15357) );
no02f80 g554623 ( .a(n_14175), .b(n_9626), .o(n_15356) );
na02f80 g554624 ( .a(n_15355), .b(n_14726), .o(n_21962) );
no02f80 g554625 ( .a(n_14184), .b(n_12420), .o(n_15851) );
no02f80 g554626 ( .a(n_13960), .b(n_14934), .o(n_20838) );
na02f80 g554627 ( .a(n_13958), .b(n_14933), .o(n_19684) );
no02f80 g554628 ( .a(n_13956), .b(n_14932), .o(n_19025) );
na02f80 g554629 ( .a(n_14671), .b(n_15354), .o(n_18053) );
no02f80 g554630 ( .a(n_13954), .b(n_14931), .o(n_17124) );
na02f80 g554631 ( .a(n_14330), .b(n_15120), .o(n_16309) );
no02f80 g554632 ( .a(n_13952), .b(n_14930), .o(n_22893) );
in01f80 g554633 ( .a(n_15118), .o(n_15119) );
na02f80 g554634 ( .a(n_14150), .b(n_9790), .o(n_15118) );
na02f80 g554635 ( .a(n_14230), .b(n_15117), .o(n_15865) );
na02f80 g554636 ( .a(n_14151), .b(n_9791), .o(n_15809) );
no02f80 g554637 ( .a(n_13947), .b(n_14929), .o(n_24444) );
na02f80 g554638 ( .a(n_14927), .b(n_14926), .o(n_14928) );
in01f80 g554639 ( .a(n_18497), .o(n_15353) );
oa12f80 g554640 ( .a(n_15040), .b(n_14118), .c(n_11751), .o(n_18497) );
no02f80 g554641 ( .a(n_15695), .b(n_15694), .o(n_16384) );
in01f80 g554642 ( .a(n_16122), .o(n_15693) );
no02f80 g554643 ( .a(n_15352), .b(n_15698), .o(n_16122) );
na02f80 g554644 ( .a(n_14217), .b(n_15116), .o(n_20854) );
oa12f80 g554645 ( .a(n_13734), .b(n_14835), .c(n_15457), .o(n_15956) );
in01f80 g554646 ( .a(n_14573), .o(n_15628) );
ao12f80 g554647 ( .a(n_12294), .b(n_14488), .c(n_12959), .o(n_14573) );
na02f80 g554648 ( .a(n_14660), .b(n_14659), .o(n_18916) );
no02f80 g554649 ( .a(n_13878), .b(n_14925), .o(n_18055) );
na02f80 g554650 ( .a(n_14441), .b(n_15115), .o(n_18063) );
ao12f80 g554651 ( .a(n_13024), .b(n_13143), .c(n_12308), .o(n_14924) );
no02f80 g554652 ( .a(n_15290), .b(n_16032), .o(n_22236) );
no02f80 g554653 ( .a(n_15351), .b(n_14656), .o(n_17964) );
na02f80 g554654 ( .a(n_15350), .b(n_14654), .o(n_21150) );
no02f80 g554655 ( .a(n_14306), .b(n_15114), .o(n_20069) );
na02f80 g554656 ( .a(n_15113), .b(n_14304), .o(n_19348) );
no02f80 g554657 ( .a(n_14302), .b(n_15112), .o(n_18352) );
na02f80 g554658 ( .a(n_15111), .b(n_14301), .o(n_17450) );
na02f80 g554659 ( .a(n_15110), .b(n_14299), .o(n_23199) );
no02f80 g554660 ( .a(n_14296), .b(n_15109), .o(n_24163) );
no02f80 g554661 ( .a(n_14903), .b(n_14902), .o(n_15759) );
no02f80 g554662 ( .a(n_16042), .b(n_15696), .o(n_15349) );
in01f80 g554663 ( .a(n_14922), .o(n_14923) );
na02f80 g554664 ( .a(n_13784), .b(n_13010), .o(n_14922) );
no02f80 g554665 ( .a(n_14439), .b(n_15107), .o(n_17134) );
na02f80 g554666 ( .a(n_13785), .b(n_13011), .o(n_15493) );
no02f80 g554667 ( .a(n_14289), .b(n_15106), .o(n_25612) );
in01f80 g554668 ( .a(n_14572), .o(n_15248) );
na02f80 g554669 ( .a(n_14076), .b(n_14565), .o(n_14572) );
no02f80 g554670 ( .a(n_14174), .b(n_9627), .o(n_15838) );
no02f80 g554671 ( .a(n_13987), .b(n_14921), .o(n_22903) );
na02f80 g554672 ( .a(n_14919), .b(n_15944), .o(n_14920) );
na02f80 g554673 ( .a(n_13806), .b(n_11064), .o(n_15545) );
no02f80 g554674 ( .a(n_14179), .b(n_9683), .o(n_15843) );
na02f80 g554675 ( .a(n_13867), .b(n_14918), .o(n_17140) );
no02f80 g554676 ( .a(n_14231), .b(n_15105), .o(n_16311) );
no02f80 g554677 ( .a(n_13981), .b(n_14917), .o(n_24173) );
no02f80 g554678 ( .a(n_14673), .b(n_15348), .o(n_18071) );
na02f80 g554679 ( .a(n_14771), .b(n_15347), .o(n_16593) );
no02f80 g554680 ( .a(n_14261), .b(n_15104), .o(n_21950) );
oa12f80 g554681 ( .a(n_11010), .b(n_14571), .c(n_12138), .o(n_15633) );
no02f80 g554682 ( .a(n_15264), .b(n_13119), .o(n_15789) );
na02f80 g554683 ( .a(n_15264), .b(n_15102), .o(n_15103) );
in01f80 g554684 ( .a(n_15961), .o(n_14916) );
na02f80 g554685 ( .a(FE_OFN1029_n_14570), .b(n_14966), .o(n_15961) );
na02f80 g554686 ( .a(n_14258), .b(n_15101), .o(n_20846) );
no02f80 g554687 ( .a(n_13922), .b(n_14915), .o(n_19692) );
na02f80 g554688 ( .a(n_14602), .b(n_15100), .o(n_15827) );
no02f80 g554689 ( .a(n_14254), .b(n_15099), .o(n_18061) );
oa12f80 g554690 ( .a(n_15027), .b(n_16004), .c(n_14095), .o(n_16445) );
no02f80 g554691 ( .a(n_14250), .b(n_15098), .o(n_16315) );
na02f80 g554692 ( .a(n_13916), .b(n_14914), .o(n_22901) );
in01f80 g554693 ( .a(n_15096), .o(n_15097) );
no02f80 g554694 ( .a(n_14144), .b(n_9770), .o(n_15096) );
no02f80 g554695 ( .a(n_14145), .b(n_9769), .o(n_15785) );
no02f80 g554696 ( .a(n_15691), .b(n_16232), .o(n_15692) );
na02f80 g554697 ( .a(n_14252), .b(n_15095), .o(n_17132) );
no02f80 g554698 ( .a(n_14569), .b(n_14568), .o(n_15546) );
no02f80 g554699 ( .a(n_14204), .b(n_11044), .o(n_15507) );
no02f80 g554700 ( .a(n_14205), .b(n_11045), .o(n_15847) );
no02f80 g554701 ( .a(n_13904), .b(n_14913), .o(n_21948) );
no02f80 g554702 ( .a(n_16243), .b(n_15691), .o(n_16408) );
na02f80 g554703 ( .a(n_13902), .b(n_14912), .o(n_20844) );
no02f80 g554704 ( .a(n_14247), .b(n_15094), .o(n_18059) );
no02f80 g554705 ( .a(n_13900), .b(n_14911), .o(n_19690) );
na02f80 g554706 ( .a(n_13898), .b(n_14910), .o(n_19031) );
na02f80 g554707 ( .a(n_14245), .b(n_15093), .o(n_17130) );
no02f80 g554708 ( .a(n_14243), .b(n_15092), .o(n_16313) );
no02f80 g554709 ( .a(n_14566), .b(n_14565), .o(n_14567) );
na02f80 g554710 ( .a(n_13892), .b(n_14909), .o(n_22899) );
na02f80 g554711 ( .a(n_14563), .b(n_14562), .o(n_14564) );
in01f80 g554712 ( .a(n_15090), .o(n_15091) );
no02f80 g554713 ( .a(n_14142), .b(n_9749), .o(n_15090) );
no02f80 g554714 ( .a(n_14143), .b(n_9748), .o(n_15778) );
no02f80 g554715 ( .a(n_14195), .b(n_11680), .o(n_15498) );
no02f80 g554716 ( .a(n_14196), .b(n_11681), .o(n_15775) );
no02f80 g554717 ( .a(n_14635), .b(n_15345), .o(n_17463) );
no02f80 g554718 ( .a(n_13885), .b(n_14908), .o(n_21944) );
ao12f80 g554719 ( .a(n_12531), .b(n_14561), .c(n_11586), .o(n_15632) );
na02f80 g554720 ( .a(n_14322), .b(n_15089), .o(n_22909) );
na02f80 g554721 ( .a(n_14781), .b(n_15344), .o(n_22243) );
no02f80 g554722 ( .a(n_14203), .b(n_11039), .o(n_15837) );
na02f80 g554723 ( .a(n_13882), .b(n_14907), .o(n_20840) );
no02f80 g554724 ( .a(n_13973), .b(n_14906), .o(n_19686) );
na02f80 g554725 ( .a(n_13872), .b(n_14905), .o(n_22895) );
in01f80 g554726 ( .a(n_15087), .o(n_15088) );
no02f80 g554727 ( .a(n_14138), .b(n_9747), .o(n_15087) );
no02f80 g554728 ( .a(n_14139), .b(n_9746), .o(n_15772) );
no02f80 g554729 ( .a(n_14760), .b(n_15343), .o(n_16168) );
no02f80 g554730 ( .a(n_14197), .b(n_11685), .o(n_15485) );
no02f80 g554731 ( .a(n_14198), .b(n_11686), .o(n_15762) );
na02f80 g554732 ( .a(n_13808), .b(n_11066), .o(n_15549) );
na02f80 g554733 ( .a(n_14215), .b(n_15086), .o(n_19043) );
no02f80 g554734 ( .a(n_16066), .b(n_15689), .o(n_15690) );
no02f80 g554735 ( .a(n_14223), .b(n_15085), .o(n_21958) );
na02f80 g554736 ( .a(n_14775), .b(n_15342), .o(n_18361) );
no02f80 g554737 ( .a(n_14287), .b(n_15084), .o(n_19700) );
no02f80 g554738 ( .a(n_13858), .b(n_14904), .o(n_16325) );
in01f80 g554739 ( .a(n_15082), .o(n_15083) );
na02f80 g554740 ( .a(n_14903), .b(n_14902), .o(n_15082) );
na02f80 g554741 ( .a(n_14178), .b(n_13588), .o(n_15840) );
oa12f80 g554742 ( .a(n_13215), .b(n_15270), .c(n_14447), .o(n_15960) );
oa12f80 g554743 ( .a(n_13663), .b(n_14789), .c(n_15295), .o(n_15959) );
oa12f80 g554744 ( .a(n_12674), .b(n_14075), .c(n_12673), .o(n_15606) );
oa12f80 g554745 ( .a(n_12845), .b(n_14560), .c(n_11088), .o(n_16186) );
ao12f80 g554746 ( .a(n_11086), .b(n_14559), .c(n_12841), .o(n_16169) );
ao12f80 g554747 ( .a(n_10605), .b(n_32732), .c(n_14073), .o(n_14982) );
oa12f80 g554748 ( .a(n_13334), .b(n_14558), .c(n_11773), .o(n_16203) );
ao12f80 g554749 ( .a(n_12551), .b(n_14557), .c(n_13728), .o(n_16196) );
in01f80 g554750 ( .a(n_14901), .o(n_15958) );
oa12f80 g554751 ( .a(n_12125), .b(n_14537), .c(n_10992), .o(n_14901) );
ao12f80 g554752 ( .a(n_11080), .b(n_14556), .c(n_12844), .o(n_16190) );
oa12f80 g554753 ( .a(n_11473), .b(n_14900), .c(n_12461), .o(n_15957) );
ao12f80 g554754 ( .a(n_11047), .b(n_14554), .c(FE_OFN1244_n_12940), .o(n_14555) );
ao12f80 g554755 ( .a(n_11456), .b(n_14072), .c(n_12447), .o(n_15246) );
ao12f80 g554756 ( .a(n_14084), .b(n_16017), .c(n_15024), .o(n_16468) );
oa12f80 g554757 ( .a(n_12846), .b(n_14553), .c(n_11084), .o(n_16208) );
ao12f80 g554758 ( .a(n_14524), .b(n_14552), .c(n_11418), .o(n_15627) );
ao12f80 g554759 ( .a(n_14071), .b(n_14531), .c(n_12315), .o(n_15626) );
ao12f80 g554760 ( .a(n_14538), .b(n_14551), .c(n_12374), .o(n_15625) );
oa12f80 g554761 ( .a(n_13607), .b(n_15445), .c(n_14798), .o(n_16242) );
oa12f80 g554762 ( .a(n_10344), .b(n_14899), .c(n_8830), .o(n_15954) );
oa12f80 g554763 ( .a(n_13848), .b(n_14898), .c(n_10153), .o(n_15953) );
ao12f80 g554764 ( .a(n_10942), .b(n_14528), .c(n_12096), .o(n_15630) );
ao12f80 g554765 ( .a(n_11042), .b(n_14550), .c(n_12807), .o(n_15882) );
ao12f80 g554766 ( .a(n_13230), .b(n_14461), .c(n_15261), .o(n_15631) );
ao12f80 g554767 ( .a(n_11721), .b(n_14897), .c(n_12793), .o(n_15952) );
ao12f80 g554768 ( .a(n_10659), .b(n_14070), .c(n_11837), .o(n_15245) );
ao12f80 g554769 ( .a(n_14529), .b(n_14549), .c(n_12329), .o(n_15624) );
ao12f80 g554770 ( .a(n_14526), .b(n_14548), .c(n_11048), .o(n_15623) );
oa12f80 g554771 ( .a(n_9533), .b(n_14547), .c(n_8322), .o(n_15629) );
oa12f80 g554772 ( .a(n_11461), .b(n_14069), .c(n_12448), .o(n_15582) );
oa12f80 g554773 ( .a(n_12349), .b(n_14546), .c(n_13107), .o(n_15866) );
in01f80 g554774 ( .a(n_16444), .o(n_23062) );
no02f80 g554775 ( .a(n_14465), .b(x_in_5_15), .o(n_16444) );
oa12f80 g554776 ( .a(n_14535), .b(n_14545), .c(n_11392), .o(n_15622) );
in01f80 g554777 ( .a(n_16804), .o(n_15081) );
oa12f80 g554778 ( .a(n_14618), .b(n_14896), .c(n_14617), .o(n_16804) );
ao12f80 g554779 ( .a(n_13825), .b(n_13798), .c(n_12815), .o(n_15539) );
in01f80 g554780 ( .a(n_15336), .o(n_15337) );
ao12f80 g554781 ( .a(n_14398), .b(n_14397), .c(n_14396), .o(n_15336) );
oa12f80 g554782 ( .a(n_14429), .b(n_14428), .c(FE_OFN1085_n_14427), .o(n_15766) );
ao12f80 g554783 ( .a(n_13995), .b(n_13994), .c(n_13993), .o(n_15531) );
in01f80 g554784 ( .a(n_15079), .o(n_15080) );
oa12f80 g554785 ( .a(n_14013), .b(n_14012), .c(n_14011), .o(n_15079) );
in01f80 g554786 ( .a(n_15687), .o(n_15688) );
ao12f80 g554787 ( .a(n_14794), .b(n_14793), .c(n_14792), .o(n_15687) );
in01f80 g554788 ( .a(n_15334), .o(n_15335) );
ao12f80 g554789 ( .a(n_14457), .b(n_14456), .c(n_14455), .o(n_15334) );
oa12f80 g554790 ( .a(n_14005), .b(n_14004), .c(n_14003), .o(n_15548) );
in01f80 g554791 ( .a(n_14894), .o(n_14895) );
oa12f80 g554792 ( .a(n_13411), .b(n_13410), .c(n_13409), .o(n_14894) );
ao12f80 g554793 ( .a(n_13446), .b(n_13445), .c(n_13444), .o(n_15949) );
in01f80 g554794 ( .a(n_15332), .o(n_15333) );
ao12f80 g554795 ( .a(n_14454), .b(n_14453), .c(n_14452), .o(n_15332) );
oa12f80 g554796 ( .a(n_14451), .b(n_14450), .c(n_14449), .o(n_15804) );
in01f80 g554797 ( .a(n_14892), .o(n_14893) );
oa12f80 g554798 ( .a(n_13443), .b(n_13442), .c(n_13441), .o(n_14892) );
ao12f80 g554799 ( .a(n_13440), .b(n_13439), .c(FE_OFN957_n_13438), .o(n_15217) );
in01f80 g554800 ( .a(n_14890), .o(n_14891) );
oa12f80 g554801 ( .a(n_13423), .b(n_13422), .c(FE_OFN953_n_13421), .o(n_14890) );
in01f80 g554802 ( .a(n_16699), .o(n_15686) );
oa12f80 g554803 ( .a(n_14809), .b(n_14808), .c(n_14807), .o(n_16699) );
in01f80 g554804 ( .a(n_14888), .o(n_14889) );
oa12f80 g554805 ( .a(n_13437), .b(n_13436), .c(n_13435), .o(n_14888) );
ao12f80 g554806 ( .a(n_14047), .b(n_14046), .c(x_in_7_12), .o(n_14887) );
oa22f80 g554807 ( .a(n_13604), .b(FE_OFN170_n_22948), .c(n_1561), .d(n_27449), .o(n_15078) );
oa22f80 g554808 ( .a(n_12569), .b(FE_OFN239_n_4162), .c(n_621), .d(FE_OFN74_n_27012), .o(n_14544) );
ao12f80 g554809 ( .a(n_14831), .b(n_14830), .c(x_in_23_12), .o(n_15331) );
oa12f80 g554810 ( .a(n_14031), .b(n_14550), .c(n_14030), .o(n_16387) );
ao12f80 g554811 ( .a(n_13452), .b(n_13451), .c(n_13450), .o(n_15223) );
oa12f80 g554812 ( .a(n_13914), .b(n_13913), .c(n_13912), .o(n_15488) );
oa22f80 g554813 ( .a(n_12568), .b(FE_OFN307_n_3069), .c(n_576), .d(FE_OFN355_n_4860), .o(n_14543) );
oa22f80 g554814 ( .a(FE_OFN857_n_12565), .b(n_27933), .c(n_1734), .d(FE_OFN64_n_27012), .o(n_14542) );
ao12f80 g554815 ( .a(n_14823), .b(n_14822), .c(x_in_47_12), .o(n_15330) );
oa12f80 g554816 ( .a(n_14815), .b(n_15329), .c(x_in_5_14), .o(n_16177) );
oa22f80 g554817 ( .a(n_12564), .b(FE_OFN303_n_3069), .c(n_369), .d(FE_OFN69_n_27012), .o(n_14541) );
in01f80 g554818 ( .a(n_16135), .o(n_15077) );
oa22f80 g554819 ( .a(n_14559), .b(n_13304), .c(n_12731), .d(n_13305), .o(n_16135) );
oa22f80 g554820 ( .a(n_12567), .b(n_28597), .c(n_227), .d(n_27449), .o(n_14540) );
ao12f80 g554821 ( .a(n_14827), .b(n_14826), .c(x_in_63_12), .o(n_15328) );
in01f80 g554822 ( .a(n_15940), .o(n_16532) );
ao12f80 g554823 ( .a(n_14064), .b(n_14063), .c(n_14062), .o(n_15940) );
in01f80 g554824 ( .a(n_15075), .o(n_15076) );
oa12f80 g554825 ( .a(n_14010), .b(n_14009), .c(n_14008), .o(n_15075) );
ao12f80 g554826 ( .a(n_14027), .b(n_14026), .c(n_15868), .o(n_14886) );
in01f80 g554827 ( .a(n_16148), .o(n_15074) );
oa22f80 g554828 ( .a(n_14553), .b(n_13341), .c(n_12803), .d(n_13342), .o(n_16148) );
oa12f80 g554829 ( .a(n_14483), .b(n_14897), .c(n_14482), .o(n_16374) );
in01f80 g554830 ( .a(n_15072), .o(n_15073) );
ao12f80 g554831 ( .a(n_13979), .b(n_13978), .c(n_13977), .o(n_15072) );
in01f80 g554832 ( .a(n_16145), .o(n_15327) );
oa22f80 g554833 ( .a(n_13751), .b(n_14558), .c(n_13752), .d(n_12790), .o(n_16145) );
ao12f80 g554834 ( .a(n_14045), .b(n_14044), .c(x_in_27_13), .o(n_14885) );
oa12f80 g554835 ( .a(n_14883), .b(n_13353), .c(n_13352), .o(n_14884) );
ao12f80 g554836 ( .a(n_13449), .b(n_13448), .c(n_13447), .o(n_15219) );
oa12f80 g554837 ( .a(n_14516), .b(n_14515), .c(n_14514), .o(n_15907) );
ao12f80 g554838 ( .a(n_14804), .b(n_14803), .c(n_14802), .o(n_15326) );
in01f80 g554839 ( .a(n_15325), .o(n_16916) );
oa12f80 g554840 ( .a(n_14513), .b(n_14512), .c(n_14511), .o(n_15325) );
oa12f80 g554841 ( .a(n_13855), .b(n_14882), .c(n_14881), .o(n_15598) );
in01f80 g554842 ( .a(n_16194), .o(n_15685) );
oa22f80 g554843 ( .a(n_14106), .b(n_14557), .c(n_14107), .d(n_12764), .o(n_16194) );
oa12f80 g554844 ( .a(n_13171), .b(n_14551), .c(n_14538), .o(n_14539) );
oa12f80 g554845 ( .a(n_13970), .b(n_14880), .c(n_14879), .o(n_15596) );
in01f80 g554846 ( .a(n_16382), .o(n_15324) );
oa12f80 g554847 ( .a(n_14498), .b(n_14551), .c(n_14497), .o(n_16382) );
in01f80 g554848 ( .a(n_16151), .o(n_15071) );
oa22f80 g554849 ( .a(n_14560), .b(n_13329), .c(n_12808), .d(n_13330), .o(n_16151) );
in01f80 g554850 ( .a(n_15069), .o(n_15070) );
ao12f80 g554851 ( .a(n_14002), .b(n_14001), .c(n_14000), .o(n_15069) );
ao12f80 g554852 ( .a(n_14829), .b(n_14828), .c(x_in_15_12), .o(n_15323) );
in01f80 g554853 ( .a(n_16141), .o(n_15068) );
oa22f80 g554854 ( .a(n_14556), .b(n_13320), .c(n_12757), .d(n_13321), .o(n_16141) );
in01f80 g554855 ( .a(n_16137), .o(n_14878) );
oa22f80 g554856 ( .a(n_14537), .b(n_12549), .c(n_12758), .d(n_12550), .o(n_16137) );
oa12f80 g554857 ( .a(n_14068), .b(n_14067), .c(x_in_1_10), .o(n_15611) );
in01f80 g554858 ( .a(n_16225), .o(n_16425) );
ao12f80 g554859 ( .a(n_14508), .b(n_14900), .c(n_14507), .o(n_16225) );
ao12f80 g554860 ( .a(n_13967), .b(n_13966), .c(n_13965), .o(n_24883) );
oa12f80 g554861 ( .a(n_13962), .b(n_14877), .c(n_14876), .o(n_15586) );
in01f80 g554862 ( .a(n_14874), .o(n_14875) );
oa12f80 g554863 ( .a(n_13426), .b(n_13425), .c(n_13424), .o(n_14874) );
ao12f80 g554864 ( .a(n_12456), .b(n_14545), .c(n_14535), .o(n_14536) );
ao12f80 g554865 ( .a(n_13420), .b(n_14534), .c(n_14533), .o(n_15226) );
in01f80 g554866 ( .a(n_16379), .o(n_15067) );
oa12f80 g554867 ( .a(n_14023), .b(n_14545), .c(n_14022), .o(n_16379) );
in01f80 g554868 ( .a(n_15529), .o(n_16453) );
oa12f80 g554869 ( .a(n_14060), .b(n_14554), .c(n_14059), .o(n_15529) );
in01f80 g554870 ( .a(n_15065), .o(n_15066) );
ao12f80 g554871 ( .a(n_13951), .b(n_13950), .c(n_13949), .o(n_15065) );
in01f80 g554872 ( .a(FE_OFN897_n_15930), .o(n_16480) );
ao12f80 g554873 ( .a(n_14020), .b(n_14547), .c(n_14019), .o(n_15930) );
ao12f80 g554874 ( .a(n_14825), .b(n_14824), .c(x_in_55_12), .o(n_15322) );
na03f80 g554875 ( .a(n_14073), .b(n_14049), .c(n_12260), .o(n_15064) );
in01f80 g554876 ( .a(n_16394), .o(n_15321) );
oa12f80 g554877 ( .a(n_14489), .b(n_14488), .c(n_14487), .o(n_16394) );
in01f80 g554878 ( .a(n_16705), .o(n_16182) );
ao12f80 g554879 ( .a(n_14504), .b(n_14503), .c(n_14502), .o(n_16705) );
oa12f80 g554880 ( .a(n_13102), .b(n_14531), .c(n_14071), .o(n_14532) );
in01f80 g554881 ( .a(n_15063), .o(n_16535) );
oa12f80 g554882 ( .a(n_14043), .b(n_14042), .c(n_14041), .o(n_15063) );
oa12f80 g554883 ( .a(n_14039), .b(n_14038), .c(n_14037), .o(n_15528) );
in01f80 g554884 ( .a(n_14872), .o(n_14873) );
ao12f80 g554885 ( .a(n_13480), .b(n_13479), .c(n_13478), .o(n_14872) );
in01f80 g554886 ( .a(n_15061), .o(n_15062) );
oa12f80 g554887 ( .a(n_14036), .b(n_14035), .c(n_14034), .o(n_15061) );
in01f80 g554888 ( .a(n_14870), .o(n_14871) );
ao12f80 g554889 ( .a(n_13477), .b(n_13476), .c(n_13475), .o(n_14870) );
in01f80 g554890 ( .a(n_14868), .o(n_14869) );
oa12f80 g554891 ( .a(n_13474), .b(n_13473), .c(n_13472), .o(n_14868) );
in01f80 g554892 ( .a(n_14866), .o(n_14867) );
ao12f80 g554893 ( .a(n_13486), .b(n_13485), .c(n_13484), .o(n_14866) );
in01f80 g554894 ( .a(n_15871), .o(n_15873) );
oa22f80 g554895 ( .a(n_32732), .b(n_12142), .c(n_14048), .d(n_12141), .o(n_15871) );
in01f80 g554896 ( .a(n_15798), .o(n_16663) );
oa12f80 g554897 ( .a(n_14471), .b(n_14898), .c(n_14470), .o(n_15798) );
oa12f80 g554898 ( .a(n_13936), .b(n_13935), .c(n_13934), .o(n_15516) );
ao12f80 g554899 ( .a(n_13941), .b(n_13940), .c(n_13939), .o(n_15514) );
in01f80 g554900 ( .a(n_15536), .o(n_16455) );
oa12f80 g554901 ( .a(n_14025), .b(n_14069), .c(n_14024), .o(n_15536) );
in01f80 g554902 ( .a(n_14864), .o(n_14865) );
ao12f80 g554903 ( .a(n_13471), .b(n_13470), .c(n_13469), .o(n_14864) );
ao12f80 g554904 ( .a(n_14658), .b(n_13523), .c(n_12888), .o(n_15060) );
in01f80 g554905 ( .a(n_15057), .o(n_15058) );
oa12f80 g554906 ( .a(n_13931), .b(n_13930), .c(n_13929), .o(n_15057) );
in01f80 g554907 ( .a(n_15489), .o(n_16441) );
oa12f80 g554908 ( .a(n_14066), .b(n_14065), .c(n_14075), .o(n_15489) );
ao12f80 g554909 ( .a(n_14033), .b(n_14032), .c(x_in_43_14), .o(n_14863) );
in01f80 g554910 ( .a(n_14861), .o(n_14862) );
ao12f80 g554911 ( .a(n_13434), .b(n_13433), .c(n_13432), .o(n_14861) );
in01f80 g554912 ( .a(n_15056), .o(n_16222) );
oa12f80 g554913 ( .a(n_14056), .b(n_14072), .c(n_14055), .o(n_15056) );
in01f80 g554914 ( .a(n_15319), .o(n_15320) );
ao12f80 g554915 ( .a(n_14284), .b(n_14283), .c(n_14282), .o(n_15319) );
oa12f80 g554916 ( .a(n_13466), .b(n_13488), .c(n_13465), .o(n_15241) );
in01f80 g554917 ( .a(n_15317), .o(n_15318) );
oa12f80 g554918 ( .a(n_14280), .b(n_14279), .c(n_14278), .o(n_15317) );
ao22s80 g554919 ( .a(n_14896), .b(n_12572), .c(n_13522), .d(x_in_24_1), .o(n_15869) );
in01f80 g554920 ( .a(n_14859), .o(n_14860) );
oa12f80 g554921 ( .a(n_13483), .b(n_13482), .c(n_13481), .o(n_14859) );
in01f80 g554922 ( .a(n_15315), .o(n_15316) );
ao12f80 g554923 ( .a(n_14270), .b(n_14269), .c(n_14268), .o(n_15315) );
in01f80 g554924 ( .a(n_15313), .o(n_15314) );
oa12f80 g554925 ( .a(n_14264), .b(n_14263), .c(n_14262), .o(n_15313) );
in01f80 g554926 ( .a(n_15862), .o(n_16212) );
ao12f80 g554927 ( .a(n_14468), .b(n_14467), .c(n_14466), .o(n_15862) );
ao12f80 g554928 ( .a(n_13416), .b(n_13415), .c(n_13414), .o(n_15212) );
in01f80 g554929 ( .a(n_15787), .o(n_15055) );
oa12f80 g554930 ( .a(n_13921), .b(n_14571), .c(n_13920), .o(n_15787) );
oa12f80 g554931 ( .a(n_13116), .b(n_14549), .c(n_14529), .o(n_14530) );
in01f80 g554932 ( .a(n_14858), .o(n_15935) );
oa22f80 g554933 ( .a(n_14528), .b(n_12533), .c(n_12718), .d(n_12532), .o(n_14858) );
in01f80 g554934 ( .a(n_16112), .o(n_15312) );
oa12f80 g554935 ( .a(n_14476), .b(n_14549), .c(n_14475), .o(n_16112) );
oa12f80 g554936 ( .a(n_13911), .b(n_13910), .c(n_13909), .o(n_16233) );
in01f80 g554937 ( .a(n_15053), .o(n_15054) );
oa12f80 g554938 ( .a(n_13908), .b(n_13907), .c(n_13906), .o(n_15053) );
in01f80 g554939 ( .a(n_15900), .o(n_15311) );
oa12f80 g554940 ( .a(n_14493), .b(n_14492), .c(n_14491), .o(n_15900) );
in01f80 g554941 ( .a(n_14857), .o(n_15937) );
oa12f80 g554942 ( .a(n_13468), .b(n_14070), .c(n_13467), .o(n_14857) );
oa12f80 g554943 ( .a(n_12222), .b(n_14548), .c(n_14526), .o(n_14527) );
in01f80 g554944 ( .a(n_15051), .o(n_15052) );
oa12f80 g554945 ( .a(n_13897), .b(n_13896), .c(n_13895), .o(n_15051) );
oa12f80 g554946 ( .a(n_13894), .b(n_14856), .c(n_14855), .o(n_15584) );
in01f80 g554947 ( .a(n_16118), .o(n_15310) );
oa12f80 g554948 ( .a(n_14474), .b(n_14548), .c(n_14473), .o(n_16118) );
in01f80 g554949 ( .a(n_16219), .o(n_16702) );
ao12f80 g554950 ( .a(n_14485), .b(n_14899), .c(n_14484), .o(n_16219) );
in01f80 g554951 ( .a(n_15049), .o(n_15050) );
oa12f80 g554952 ( .a(n_14016), .b(n_14015), .c(n_14014), .o(n_15049) );
in01f80 g554953 ( .a(n_14853), .o(n_14854) );
ao12f80 g554954 ( .a(n_13408), .b(n_13407), .c(n_13406), .o(n_14853) );
in01f80 g554955 ( .a(n_14851), .o(n_14852) );
oa12f80 g554956 ( .a(n_13464), .b(n_13463), .c(n_13462), .o(n_14851) );
in01f80 g554957 ( .a(n_15047), .o(n_15048) );
oa12f80 g554958 ( .a(n_13891), .b(n_13890), .c(n_13889), .o(n_15047) );
in01f80 g554959 ( .a(n_14849), .o(n_14850) );
ao12f80 g554960 ( .a(n_13461), .b(n_13460), .c(n_13459), .o(n_14849) );
in01f80 g554961 ( .a(n_14847), .o(n_14848) );
oa12f80 g554962 ( .a(n_13458), .b(n_13457), .c(n_13456), .o(n_14847) );
in01f80 g554963 ( .a(n_15308), .o(n_15309) );
oa12f80 g554964 ( .a(n_14242), .b(n_14241), .c(n_14240), .o(n_15308) );
in01f80 g554965 ( .a(n_15306), .o(n_15307) );
oa12f80 g554966 ( .a(n_14239), .b(n_14238), .c(n_14237), .o(n_15306) );
ao12f80 g554967 ( .a(n_13455), .b(n_13454), .c(n_13453), .o(n_15210) );
in01f80 g554968 ( .a(n_14845), .o(n_14846) );
oa12f80 g554969 ( .a(n_13402), .b(n_13401), .c(n_13400), .o(n_14845) );
ao12f80 g554970 ( .a(n_13888), .b(n_13887), .c(n_13886), .o(n_15491) );
in01f80 g554971 ( .a(n_14843), .o(n_14844) );
ao12f80 g554972 ( .a(n_13419), .b(n_13418), .c(n_13417), .o(n_14843) );
in01f80 g554973 ( .a(n_15600), .o(n_15897) );
ao12f80 g554974 ( .a(n_14053), .b(n_14561), .c(n_14052), .o(n_15600) );
oa12f80 g554975 ( .a(n_14464), .b(n_14463), .c(n_14546), .o(n_16117) );
in01f80 g554976 ( .a(n_15045), .o(n_15046) );
oa12f80 g554977 ( .a(n_13871), .b(n_13870), .c(n_13869), .o(n_15045) );
ao12f80 g554978 ( .a(n_13431), .b(n_13430), .c(n_13429), .o(n_15207) );
ao12f80 g554979 ( .a(n_14821), .b(n_14820), .c(x_in_31_12), .o(n_15305) );
in01f80 g554980 ( .a(n_15303), .o(n_15304) );
ao12f80 g554981 ( .a(n_14228), .b(n_14227), .c(n_14226), .o(n_15303) );
in01f80 g554982 ( .a(n_15043), .o(n_15044) );
oa12f80 g554983 ( .a(n_13866), .b(n_13865), .c(n_13864), .o(n_15043) );
in01f80 g554984 ( .a(n_15301), .o(n_15302) );
ao12f80 g554985 ( .a(n_14275), .b(n_14274), .c(FE_OFN1081_n_14273), .o(n_15301) );
oa12f80 g554986 ( .a(n_12433), .b(n_14552), .c(n_14524), .o(n_14525) );
ao12f80 g554987 ( .a(n_13405), .b(n_13404), .c(n_13403), .o(n_15945) );
in01f80 g554988 ( .a(n_15299), .o(n_15300) );
oa12f80 g554989 ( .a(n_14221), .b(n_14220), .c(n_14219), .o(n_15299) );
in01f80 g554990 ( .a(n_15041), .o(n_15042) );
ao12f80 g554991 ( .a(n_13861), .b(n_13860), .c(n_13859), .o(n_15041) );
oa22f80 g554992 ( .a(FE_OFN979_n_12566), .b(n_27933), .c(n_1315), .d(FE_OFN68_n_27012), .o(n_14523) );
in01f80 g554993 ( .a(n_14841), .o(n_14842) );
ao12f80 g554994 ( .a(n_13395), .b(n_13394), .c(n_13393), .o(n_14841) );
in01f80 g554995 ( .a(FE_OFN628_n_15605), .o(n_15916) );
ao12f80 g554996 ( .a(n_14051), .b(n_14552), .c(n_14050), .o(n_15605) );
in01f80 g554997 ( .a(n_16114), .o(n_15298) );
oa12f80 g554998 ( .a(n_14518), .b(n_14531), .c(n_14517), .o(n_16114) );
oa22f80 g554999 ( .a(n_12680), .b(FE_OFN300_n_3069), .c(n_1877), .d(FE_OFN91_n_27449), .o(n_14522) );
oa22f80 g555000 ( .a(n_12672), .b(FE_OFN7_n_28597), .c(n_1774), .d(FE_OFN78_n_27012), .o(n_14521) );
oa22f80 g555001 ( .a(n_12578), .b(FE_OFN411_n_28303), .c(n_1160), .d(FE_OFN335_n_4860), .o(n_14520) );
oa22f80 g555002 ( .a(n_12677), .b(FE_OFN7_n_28597), .c(n_1128), .d(FE_OFN336_n_4860), .o(n_14519) );
ao22s80 g555003 ( .a(n_13225), .b(n_11393), .c(x_out_55_19), .d(n_16656), .o(n_14840) );
na02f80 g555025 ( .a(n_14067), .b(x_in_1_10), .o(n_14068) );
na02f80 g555026 ( .a(n_14054), .b(x_in_4_8), .o(n_15108) );
na02f80 g555027 ( .a(n_15040), .b(n_14119), .o(n_15709) );
na02f80 g555028 ( .a(n_15039), .b(n_14121), .o(n_15712) );
na02f80 g555029 ( .a(n_14065), .b(n_14075), .o(n_14066) );
na02f80 g555030 ( .a(n_14531), .b(n_14517), .o(n_14518) );
no02f80 g555031 ( .a(n_14063), .b(n_14062), .o(n_14064) );
na02f80 g555032 ( .a(n_13488), .b(n_13487), .o(n_14992) );
na02f80 g555033 ( .a(n_14515), .b(n_14514), .o(n_14516) );
na02f80 g555034 ( .a(n_14512), .b(n_14511), .o(n_14513) );
na02f80 g555035 ( .a(n_14510), .b(n_14509), .o(n_15655) );
in01f80 g555036 ( .a(n_14838), .o(n_14839) );
no02f80 g555037 ( .a(n_14510), .b(n_14509), .o(n_14838) );
no02f80 g555038 ( .a(n_14900), .b(n_14507), .o(n_14508) );
na02f80 g555039 ( .a(n_14061), .b(x_in_0_8), .o(n_15275) );
in01f80 g555040 ( .a(n_14505), .o(n_14506) );
no02f80 g555041 ( .a(n_14061), .b(x_in_0_8), .o(n_14505) );
in01f80 g555042 ( .a(n_15037), .o(n_15038) );
na02f80 g555043 ( .a(n_14837), .b(n_13745), .o(n_15037) );
na02f80 g555044 ( .a(n_14554), .b(n_14059), .o(n_14060) );
in01f80 g555045 ( .a(n_14057), .o(n_14058) );
no02f80 g555046 ( .a(n_13488), .b(n_13487), .o(n_14057) );
no02f80 g555047 ( .a(n_14836), .b(n_13737), .o(n_22889) );
no02f80 g555048 ( .a(n_13735), .b(n_14835), .o(n_15458) );
na02f80 g555049 ( .a(n_14072), .b(n_14055), .o(n_14056) );
no02f80 g555050 ( .a(n_14503), .b(n_14502), .o(n_14504) );
in01f80 g555051 ( .a(n_14500), .o(n_14501) );
no02f80 g555052 ( .a(n_14054), .b(x_in_4_8), .o(n_14500) );
in01f80 g555053 ( .a(n_14833), .o(n_14834) );
na02f80 g555054 ( .a(n_14499), .b(n_13300), .o(n_14833) );
no02f80 g555055 ( .a(n_14561), .b(n_14052), .o(n_14053) );
no02f80 g555056 ( .a(n_14552), .b(n_14050), .o(n_14051) );
na02f80 g555057 ( .a(n_14551), .b(n_14497), .o(n_14498) );
in01f80 g555058 ( .a(n_14496), .o(n_15265) );
na02f80 g555059 ( .a(n_14067), .b(n_260), .o(n_14496) );
na02f80 g555060 ( .a(n_14048), .b(n_11372), .o(n_14049) );
no02f80 g555061 ( .a(n_13485), .b(n_13484), .o(n_13486) );
no02f80 g555062 ( .a(n_13310), .b(n_14477), .o(n_14495) );
na02f80 g555063 ( .a(n_13311), .b(n_14494), .o(n_16868) );
no02f80 g555064 ( .a(n_13717), .b(n_14832), .o(n_23845) );
no02f80 g555065 ( .a(n_14830), .b(x_in_23_12), .o(n_14831) );
no02f80 g555066 ( .a(n_14828), .b(x_in_15_12), .o(n_14829) );
no02f80 g555067 ( .a(n_14826), .b(x_in_63_12), .o(n_14827) );
no02f80 g555068 ( .a(n_14824), .b(x_in_55_12), .o(n_14825) );
no02f80 g555069 ( .a(n_14822), .b(x_in_47_12), .o(n_14823) );
no02f80 g555070 ( .a(n_14820), .b(x_in_31_12), .o(n_14821) );
no02f80 g555071 ( .a(n_14046), .b(x_in_7_12), .o(n_14047) );
na02f80 g555072 ( .a(n_13482), .b(n_13481), .o(n_13483) );
no02f80 g555073 ( .a(n_14044), .b(x_in_27_13), .o(n_14045) );
na02f80 g555074 ( .a(n_14042), .b(n_14041), .o(n_14043) );
na02f80 g555075 ( .a(n_14492), .b(n_14491), .o(n_14493) );
na02f80 g555076 ( .a(n_14040), .b(n_15186), .o(n_14991) );
na02f80 g555077 ( .a(n_14038), .b(n_14037), .o(n_14039) );
no02f80 g555078 ( .a(n_13479), .b(n_13478), .o(n_13480) );
na02f80 g555079 ( .a(n_14035), .b(n_14034), .o(n_14036) );
no02f80 g555080 ( .a(n_13476), .b(n_13475), .o(n_13477) );
na02f80 g555081 ( .a(n_13473), .b(n_13472), .o(n_13474) );
in01f80 g555082 ( .a(n_14818), .o(n_14819) );
na02f80 g555083 ( .a(n_14490), .b(n_13276), .o(n_14818) );
na02f80 g555084 ( .a(n_14488), .b(n_14487), .o(n_14489) );
no02f80 g555085 ( .a(n_13470), .b(n_13469), .o(n_13471) );
no02f80 g555086 ( .a(n_14032), .b(x_in_43_14), .o(n_14033) );
na02f80 g555087 ( .a(n_14550), .b(n_14030), .o(n_14031) );
in01f80 g555088 ( .a(n_14816), .o(n_14817) );
na02f80 g555089 ( .a(n_13274), .b(n_14486), .o(n_14816) );
na02f80 g555090 ( .a(n_15329), .b(x_in_5_14), .o(n_14815) );
no02f80 g555091 ( .a(n_14899), .b(n_14484), .o(n_14485) );
na02f80 g555092 ( .a(n_14897), .b(n_14482), .o(n_14483) );
in01f80 g555093 ( .a(n_15645), .o(n_16023) );
na02f80 g555094 ( .a(n_14826), .b(n_8206), .o(n_15645) );
in01f80 g555095 ( .a(n_15643), .o(n_15996) );
na02f80 g555096 ( .a(n_14828), .b(n_7338), .o(n_15643) );
in01f80 g555097 ( .a(n_15671), .o(n_15036) );
na02f80 g555098 ( .a(n_14824), .b(n_7278), .o(n_15671) );
in01f80 g555099 ( .a(n_15670), .o(n_15035) );
na02f80 g555100 ( .a(n_14830), .b(n_7323), .o(n_15670) );
na02f80 g555101 ( .a(n_14070), .b(n_13467), .o(n_13468) );
in01f80 g555102 ( .a(n_15649), .o(n_15999) );
na02f80 g555103 ( .a(n_14822), .b(n_7247), .o(n_15649) );
in01f80 g555104 ( .a(n_15280), .o(n_15034) );
na02f80 g555105 ( .a(n_14820), .b(n_6753), .o(n_15280) );
in01f80 g555106 ( .a(n_14481), .o(n_25819) );
no02f80 g555107 ( .a(n_14029), .b(n_14028), .o(n_14481) );
in01f80 g555108 ( .a(n_14479), .o(n_14480) );
na02f80 g555109 ( .a(n_14029), .b(n_14028), .o(n_14479) );
in01f80 g555110 ( .a(n_14594), .o(n_14478) );
na02f80 g555111 ( .a(n_14046), .b(n_7340), .o(n_14594) );
na02f80 g555112 ( .a(n_13488), .b(n_11856), .o(n_15661) );
na02f80 g555113 ( .a(n_13488), .b(n_13465), .o(n_13466) );
in01f80 g555114 ( .a(n_15032), .o(n_15033) );
na02f80 g555115 ( .a(n_14814), .b(n_13702), .o(n_15032) );
no02f80 g555116 ( .a(n_14477), .b(n_16297), .o(n_15971) );
na02f80 g555117 ( .a(n_14549), .b(n_14475), .o(n_14476) );
na02f80 g555118 ( .a(n_14548), .b(n_14473), .o(n_14474) );
in01f80 g555119 ( .a(n_14472), .o(n_15059) );
na02f80 g555120 ( .a(n_14044), .b(n_7229), .o(n_14472) );
na02f80 g555121 ( .a(n_14898), .b(n_14470), .o(n_14471) );
na02f80 g555122 ( .a(n_15031), .b(x_in_42_1), .o(n_16069) );
no02f80 g555123 ( .a(n_15031), .b(x_in_42_1), .o(n_16068) );
no02f80 g555124 ( .a(n_14812), .b(x_in_58_1), .o(n_15736) );
na02f80 g555125 ( .a(n_14813), .b(x_in_2_1), .o(n_16067) );
no02f80 g555126 ( .a(n_14813), .b(x_in_2_1), .o(n_16065) );
na02f80 g555127 ( .a(n_14812), .b(x_in_58_1), .o(n_15737) );
na02f80 g555128 ( .a(n_15029), .b(x_in_10_1), .o(n_16059) );
na02f80 g555129 ( .a(n_15682), .b(x_in_34_1), .o(n_16644) );
no02f80 g555130 ( .a(n_15682), .b(x_in_34_1), .o(n_16643) );
na02f80 g555131 ( .a(n_14811), .b(x_in_16_1), .o(n_15747) );
no02f80 g555132 ( .a(n_14811), .b(x_in_16_1), .o(n_15746) );
no02f80 g555133 ( .a(n_14469), .b(x_in_18_1), .o(n_15743) );
na02f80 g555134 ( .a(n_14469), .b(x_in_18_1), .o(n_15744) );
na02f80 g555135 ( .a(n_15030), .b(x_in_50_1), .o(n_16062) );
no02f80 g555136 ( .a(n_15030), .b(x_in_50_1), .o(n_16061) );
no02f80 g555137 ( .a(n_15029), .b(x_in_10_1), .o(n_16058) );
na02f80 g555138 ( .a(n_15028), .b(x_in_26_1), .o(n_16057) );
no02f80 g555139 ( .a(n_15028), .b(x_in_26_1), .o(n_16056) );
no02f80 g555140 ( .a(n_14100), .b(n_14810), .o(n_22582) );
no02f80 g555141 ( .a(n_14467), .b(n_14466), .o(n_14468) );
no02f80 g555142 ( .a(n_14026), .b(n_15868), .o(n_14027) );
na02f80 g555143 ( .a(n_14808), .b(n_14807), .o(n_14809) );
na02f80 g555144 ( .a(n_14032), .b(n_7311), .o(n_15005) );
no02f80 g555145 ( .a(n_13690), .b(x_in_5_14), .o(n_14465) );
na02f80 g555146 ( .a(n_14069), .b(n_14024), .o(n_14025) );
na02f80 g555147 ( .a(n_14463), .b(n_14546), .o(n_14464) );
no02f80 g555148 ( .a(n_14462), .b(n_12930), .o(n_23405) );
na02f80 g555149 ( .a(n_14545), .b(n_14022), .o(n_14023) );
na02f80 g555150 ( .a(n_12704), .b(n_14021), .o(n_22741) );
no02f80 g555151 ( .a(n_14547), .b(n_14019), .o(n_14020) );
na02f80 g555152 ( .a(n_14096), .b(n_15027), .o(n_16005) );
no02f80 g555153 ( .a(n_13529), .b(n_9539), .o(n_15753) );
na02f80 g555154 ( .a(n_14461), .b(n_13231), .o(n_15262) );
na02f80 g555155 ( .a(n_14093), .b(n_14806), .o(n_23572) );
na02f80 g555156 ( .a(n_14040), .b(n_14460), .o(n_15187) );
na02f80 g555157 ( .a(n_13681), .b(n_14805), .o(n_23190) );
no02f80 g555158 ( .a(n_14803), .b(n_14802), .o(n_14804) );
na02f80 g555159 ( .a(n_14801), .b(n_13679), .o(n_23489) );
in01f80 g555160 ( .a(n_14458), .o(n_14459) );
na02f80 g555161 ( .a(n_14018), .b(n_14017), .o(n_14458) );
no02f80 g555162 ( .a(n_14018), .b(n_14017), .o(n_15011) );
in01f80 g555163 ( .a(n_14799), .o(n_14800) );
no02f80 g555164 ( .a(n_13546), .b(n_10744), .o(n_14799) );
no02f80 g555165 ( .a(n_13547), .b(n_10745), .o(n_15433) );
na02f80 g555166 ( .a(n_14015), .b(n_14014), .o(n_14016) );
na02f80 g555167 ( .a(n_13463), .b(n_13462), .o(n_13464) );
no02f80 g555168 ( .a(n_13460), .b(n_13459), .o(n_13461) );
na02f80 g555169 ( .a(n_13457), .b(n_13456), .o(n_13458) );
no02f80 g555170 ( .a(n_13454), .b(n_13453), .o(n_13455) );
na02f80 g555171 ( .a(n_13938), .b(n_13937), .o(n_15111) );
no02f80 g555172 ( .a(n_13606), .b(n_14798), .o(n_15446) );
in01f80 g555173 ( .a(n_14796), .o(n_14797) );
na02f80 g555174 ( .a(n_13584), .b(n_11724), .o(n_14796) );
na02f80 g555175 ( .a(n_14012), .b(n_14011), .o(n_14013) );
no02f80 g555176 ( .a(n_13657), .b(n_14795), .o(n_15607) );
no02f80 g555177 ( .a(n_13451), .b(n_13450), .o(n_13452) );
no02f80 g555178 ( .a(n_13983), .b(n_13982), .o(n_15157) );
no02f80 g555179 ( .a(n_14793), .b(n_14792), .o(n_14794) );
no02f80 g555180 ( .a(n_13392), .b(n_13391), .o(n_14904) );
na02f80 g555181 ( .a(n_14009), .b(n_14008), .o(n_14010) );
no02f80 g555182 ( .a(n_14456), .b(n_14455), .o(n_14457) );
in01f80 g555183 ( .a(n_14006), .o(n_14007) );
no02f80 g555184 ( .a(n_13428), .b(n_13427), .o(n_14006) );
na02f80 g555185 ( .a(n_14004), .b(n_14003), .o(n_14005) );
na02f80 g555186 ( .a(n_13413), .b(n_13412), .o(n_15950) );
na02f80 g555187 ( .a(n_13672), .b(n_14791), .o(n_23214) );
no02f80 g555188 ( .a(n_13448), .b(n_13447), .o(n_13449) );
no02f80 g555189 ( .a(n_13445), .b(n_13444), .o(n_13446) );
no02f80 g555190 ( .a(n_14453), .b(n_14452), .o(n_14454) );
na02f80 g555191 ( .a(n_14450), .b(n_14449), .o(n_14451) );
oa12f80 g555192 ( .a(FE_OFN396_n_14720), .b(n_1431), .c(FE_OFN364_n_4860), .o(n_14790) );
no02f80 g555193 ( .a(n_14001), .b(n_14000), .o(n_14002) );
no02f80 g555194 ( .a(n_13664), .b(n_14789), .o(n_15296) );
na02f80 g555195 ( .a(n_13442), .b(n_13441), .o(n_13443) );
no02f80 g555196 ( .a(n_13666), .b(n_14788), .o(n_16602) );
na02f80 g555197 ( .a(n_13668), .b(n_14787), .o(n_17465) );
no02f80 g555198 ( .a(n_13670), .b(n_14786), .o(n_18364) );
na02f80 g555199 ( .a(n_13219), .b(n_14448), .o(n_21165) );
no03m80 g555200 ( .a(x_in_39_11), .b(n_14595), .c(x_in_39_12), .o(n_15268) );
in01f80 g555201 ( .a(n_13998), .o(n_13999) );
na02f80 g555202 ( .a(n_12678), .b(n_12323), .o(n_13998) );
no02f80 g555203 ( .a(n_13863), .b(n_13862), .o(n_15085) );
no02f80 g555204 ( .a(n_13439), .b(FE_OFN957_n_13438), .o(n_13440) );
no02f80 g555205 ( .a(n_13214), .b(n_14447), .o(n_15271) );
oa12f80 g555206 ( .a(n_12535), .b(n_14807), .c(n_13718), .o(n_15205) );
na02f80 g555207 ( .a(n_13609), .b(n_14785), .o(n_19362) );
in01f80 g555208 ( .a(n_14445), .o(n_14446) );
no02f80 g555209 ( .a(n_13079), .b(n_10163), .o(n_14445) );
na02f80 g555210 ( .a(n_12679), .b(n_12324), .o(n_14958) );
no02f80 g555211 ( .a(n_13080), .b(n_10162), .o(n_15170) );
na02f80 g555212 ( .a(n_13436), .b(n_13435), .o(n_13437) );
in01f80 g555213 ( .a(n_13996), .o(n_13997) );
na02f80 g555214 ( .a(n_12675), .b(n_11735), .o(n_13996) );
in01f80 g555215 ( .a(n_14783), .o(n_14784) );
no02f80 g555216 ( .a(n_13590), .b(n_12402), .o(n_14783) );
in01f80 g555217 ( .a(n_14443), .o(n_14444) );
no02f80 g555218 ( .a(n_13033), .b(n_11069), .o(n_14443) );
no02f80 g555219 ( .a(n_13994), .b(n_13993), .o(n_13995) );
no02f80 g555220 ( .a(n_13433), .b(n_13432), .o(n_13434) );
in01f80 g555221 ( .a(n_14441), .o(n_14442) );
na02f80 g555222 ( .a(n_13086), .b(n_11733), .o(n_14441) );
in01f80 g555223 ( .a(n_14439), .o(n_14440) );
no02f80 g555224 ( .a(n_12989), .b(n_11051), .o(n_14439) );
na02f80 g555225 ( .a(n_13087), .b(n_11734), .o(n_15115) );
oa12f80 g555226 ( .a(n_13990), .b(n_108), .c(FE_OFN350_n_4860), .o(n_13992) );
in01f80 g555227 ( .a(n_14781), .o(n_14782) );
na02f80 g555228 ( .a(n_13602), .b(n_12886), .o(n_14781) );
no02f80 g555229 ( .a(n_12990), .b(n_11050), .o(n_15107) );
in01f80 g555230 ( .a(n_14437), .o(n_14438) );
na02f80 g555231 ( .a(n_12991), .b(n_11731), .o(n_14437) );
oa12f80 g555232 ( .a(n_13990), .b(n_382), .c(FE_OFN136_n_27449), .o(n_13991) );
na02f80 g555233 ( .a(n_13603), .b(n_12887), .o(n_15344) );
in01f80 g555234 ( .a(n_14779), .o(n_14780) );
no02f80 g555235 ( .a(n_13532), .b(n_12417), .o(n_14779) );
no02f80 g555236 ( .a(n_13533), .b(n_12418), .o(n_15416) );
na02f80 g555237 ( .a(n_14214), .b(n_14213), .o(n_15415) );
oa12f80 g555238 ( .a(FE_OFN379_n_13985), .b(n_1902), .c(n_28607), .o(n_13989) );
no02f80 g555239 ( .a(n_13944), .b(n_13943), .o(n_15169) );
in01f80 g555240 ( .a(n_14777), .o(n_14778) );
no02f80 g555241 ( .a(n_13600), .b(n_12414), .o(n_14777) );
in01f80 g555242 ( .a(n_14775), .o(n_14776) );
na02f80 g555243 ( .a(n_13598), .b(n_11739), .o(n_14775) );
in01f80 g555244 ( .a(n_14773), .o(n_14774) );
no02f80 g555245 ( .a(n_13596), .b(n_9085), .o(n_14773) );
in01f80 g555246 ( .a(n_13987), .o(n_13988) );
no02f80 g555247 ( .a(n_12666), .b(n_10161), .o(n_13987) );
in01f80 g555248 ( .a(n_14771), .o(n_14772) );
na02f80 g555249 ( .a(n_13516), .b(n_12427), .o(n_14771) );
no02f80 g555250 ( .a(n_12667), .b(n_10160), .o(n_14921) );
oa12f80 g555251 ( .a(FE_OFN379_n_13985), .b(n_1856), .c(n_28928), .o(n_13986) );
no02f80 g555252 ( .a(n_13430), .b(n_13429), .o(n_13431) );
oa12f80 g555253 ( .a(FE_OFN377_n_14285), .b(n_1753), .c(FE_OFN93_n_27449), .o(n_14436) );
na02f80 g555254 ( .a(n_13599), .b(n_11740), .o(n_15342) );
in01f80 g555255 ( .a(n_14769), .o(n_14770) );
na02f80 g555256 ( .a(n_13582), .b(n_12347), .o(n_14769) );
in01f80 g555257 ( .a(n_14767), .o(n_14768) );
no02f80 g555258 ( .a(n_13514), .b(n_12404), .o(n_14767) );
na02f80 g555259 ( .a(n_13583), .b(n_12348), .o(n_15431) );
no02f80 g555260 ( .a(n_13515), .b(n_12405), .o(n_15410) );
na02f80 g555261 ( .a(n_14435), .b(n_14434), .o(n_15412) );
in01f80 g555262 ( .a(n_14765), .o(n_14766) );
no02f80 g555263 ( .a(n_14435), .b(n_14434), .o(n_14765) );
na02f80 g555264 ( .a(n_13428), .b(n_13427), .o(n_14962) );
na02f80 g555265 ( .a(n_14431), .b(n_14430), .o(n_15423) );
in01f80 g555266 ( .a(n_14763), .o(n_14764) );
no02f80 g555267 ( .a(n_13592), .b(n_12386), .o(n_14763) );
no02f80 g555268 ( .a(n_13591), .b(n_12403), .o(n_15426) );
in01f80 g555269 ( .a(n_14761), .o(n_14762) );
na02f80 g555270 ( .a(n_13586), .b(n_11766), .o(n_14761) );
na02f80 g555271 ( .a(n_13587), .b(n_11767), .o(n_15432) );
no02f80 g555272 ( .a(n_14433), .b(n_14432), .o(n_15343) );
no02f80 g555273 ( .a(n_13097), .b(n_11483), .o(n_15477) );
in01f80 g555274 ( .a(n_14759), .o(n_14760) );
na02f80 g555275 ( .a(n_14433), .b(n_14432), .o(n_14759) );
oa12f80 g555276 ( .a(n_14694), .b(n_1107), .c(FE_OFN89_n_27449), .o(n_14758) );
na02f80 g555277 ( .a(n_12676), .b(n_11736), .o(n_14961) );
in01f80 g555278 ( .a(n_14756), .o(n_14757) );
no02f80 g555279 ( .a(n_13580), .b(n_12406), .o(n_14756) );
no02f80 g555280 ( .a(n_14324), .b(n_14323), .o(n_15403) );
in01f80 g555281 ( .a(n_14754), .o(n_14755) );
no02f80 g555282 ( .a(n_14431), .b(n_14430), .o(n_14754) );
oa12f80 g555283 ( .a(n_13924), .b(n_125), .c(FE_OFN116_n_27449), .o(n_13984) );
na02f80 g555284 ( .a(n_14428), .b(FE_OFN1085_n_14427), .o(n_14429) );
no02f80 g555285 ( .a(n_14423), .b(n_14422), .o(n_15409) );
na02f80 g555286 ( .a(n_13585), .b(n_11725), .o(n_15408) );
in01f80 g555287 ( .a(n_14752), .o(n_14753) );
na02f80 g555288 ( .a(n_14358), .b(n_14357), .o(n_14752) );
in01f80 g555289 ( .a(n_14424), .o(n_14425) );
na02f80 g555290 ( .a(n_13031), .b(n_11406), .o(n_14424) );
in01f80 g555291 ( .a(n_14750), .o(n_14751) );
na02f80 g555292 ( .a(n_14423), .b(n_14422), .o(n_14750) );
na02f80 g555293 ( .a(n_14749), .b(n_13653), .o(n_16319) );
in01f80 g555294 ( .a(n_14420), .o(n_14421) );
na02f80 g555295 ( .a(n_13983), .b(n_13982), .o(n_14420) );
no02f80 g555296 ( .a(n_14212), .b(n_14211), .o(n_15345) );
na02f80 g555297 ( .a(n_14236), .b(n_14235), .o(n_15404) );
in01f80 g555298 ( .a(n_14418), .o(n_14419) );
na02f80 g555299 ( .a(n_13077), .b(n_9704), .o(n_14418) );
na02f80 g555300 ( .a(n_13078), .b(n_9705), .o(n_15156) );
in01f80 g555301 ( .a(n_14416), .o(n_14417) );
no02f80 g555302 ( .a(n_13073), .b(n_10564), .o(n_14416) );
no02f80 g555303 ( .a(n_13074), .b(n_10565), .o(n_15155) );
in01f80 g555304 ( .a(n_14414), .o(n_14415) );
na02f80 g555305 ( .a(n_13071), .b(n_10581), .o(n_14414) );
no02f80 g555306 ( .a(n_13204), .b(n_14413), .o(n_17136) );
na02f80 g555307 ( .a(n_13072), .b(n_10580), .o(n_15154) );
na02f80 g555308 ( .a(n_14412), .b(n_13202), .o(n_18065) );
in01f80 g555309 ( .a(n_14410), .o(n_14411) );
no02f80 g555310 ( .a(n_13069), .b(n_9738), .o(n_14410) );
no02f80 g555311 ( .a(n_13070), .b(n_9737), .o(n_15153) );
in01f80 g555312 ( .a(n_14408), .o(n_14409) );
na02f80 g555313 ( .a(n_13067), .b(n_11722), .o(n_14408) );
na02f80 g555314 ( .a(n_14294), .b(n_14293), .o(n_15406) );
na02f80 g555315 ( .a(n_13068), .b(n_11723), .o(n_15152) );
in01f80 g555316 ( .a(n_14406), .o(n_14407) );
no02f80 g555317 ( .a(n_13065), .b(n_11036), .o(n_14406) );
no02f80 g555318 ( .a(n_13200), .b(n_14405), .o(n_19037) );
no02f80 g555319 ( .a(n_13066), .b(n_11035), .o(n_15151) );
in01f80 g555320 ( .a(n_14403), .o(n_14404) );
no02f80 g555321 ( .a(n_13919), .b(n_13918), .o(n_14403) );
oa12f80 g555322 ( .a(FE_OFN393_n_14663), .b(n_1756), .c(FE_OFN93_n_27449), .o(n_14748) );
na02f80 g555323 ( .a(n_13650), .b(n_14402), .o(n_19696) );
na02f80 g555324 ( .a(n_14401), .b(n_14400), .o(n_15400) );
in01f80 g555325 ( .a(n_14746), .o(n_14747) );
no02f80 g555326 ( .a(n_14401), .b(n_14400), .o(n_14746) );
in01f80 g555327 ( .a(n_14744), .o(n_14745) );
no02f80 g555328 ( .a(n_13578), .b(n_12396), .o(n_14744) );
no02f80 g555329 ( .a(n_13579), .b(n_12397), .o(n_15399) );
na02f80 g555330 ( .a(n_14393), .b(n_14392), .o(n_15398) );
no02f80 g555331 ( .a(n_13648), .b(n_14399), .o(n_20850) );
no02f80 g555332 ( .a(n_14397), .b(n_14396), .o(n_14398) );
in01f80 g555333 ( .a(n_14394), .o(n_14395) );
no02f80 g555334 ( .a(n_13063), .b(n_9700), .o(n_14394) );
in01f80 g555335 ( .a(n_14742), .o(n_14743) );
no02f80 g555336 ( .a(n_14393), .b(n_14392), .o(n_14742) );
in01f80 g555337 ( .a(n_14740), .o(n_14741) );
no02f80 g555338 ( .a(n_13576), .b(n_12394), .o(n_14740) );
no02f80 g555339 ( .a(n_13577), .b(n_12395), .o(n_15397) );
in01f80 g555340 ( .a(n_14738), .o(n_14739) );
na02f80 g555341 ( .a(n_13574), .b(n_12392), .o(n_14738) );
na02f80 g555342 ( .a(n_13425), .b(n_13424), .o(n_13426) );
no02f80 g555343 ( .a(n_13064), .b(n_9699), .o(n_15150) );
na02f80 g555344 ( .a(n_13575), .b(n_12393), .o(n_15396) );
in01f80 g555345 ( .a(n_14736), .o(n_14737) );
no02f80 g555346 ( .a(n_13572), .b(n_12390), .o(n_14736) );
no02f80 g555347 ( .a(n_13573), .b(n_12391), .o(n_15395) );
in01f80 g555348 ( .a(n_14734), .o(n_14735) );
na02f80 g555349 ( .a(n_13570), .b(n_11764), .o(n_14734) );
na02f80 g555350 ( .a(n_13197), .b(n_14391), .o(n_21954) );
na02f80 g555351 ( .a(n_13571), .b(n_11765), .o(n_15394) );
no02f80 g555352 ( .a(n_14390), .b(n_14389), .o(n_15393) );
in01f80 g555353 ( .a(n_14732), .o(n_14733) );
na02f80 g555354 ( .a(n_14390), .b(n_14389), .o(n_14732) );
in01f80 g555355 ( .a(n_13980), .o(n_13981) );
na02f80 g555356 ( .a(n_13397), .b(n_13396), .o(n_13980) );
no02f80 g555357 ( .a(n_13601), .b(n_12415), .o(n_15414) );
no02f80 g555358 ( .a(n_13978), .b(n_13977), .o(n_13979) );
no02f80 g555359 ( .a(n_13646), .b(n_14388), .o(n_22905) );
na02f80 g555360 ( .a(n_14387), .b(n_13196), .o(n_23861) );
na02f80 g555361 ( .a(n_13061), .b(n_10482), .o(n_14883) );
na02f80 g555362 ( .a(n_13062), .b(n_10483), .o(n_15137) );
no02f80 g555363 ( .a(n_13976), .b(n_13975), .o(n_15145) );
na02f80 g555364 ( .a(n_14088), .b(n_15025), .o(n_25631) );
in01f80 g555365 ( .a(n_14385), .o(n_14386) );
na02f80 g555366 ( .a(n_13976), .b(n_13975), .o(n_14385) );
in01f80 g555367 ( .a(n_14383), .o(n_14384) );
na02f80 g555368 ( .a(n_13059), .b(n_11747), .o(n_14383) );
na02f80 g555369 ( .a(n_13060), .b(n_11748), .o(n_15144) );
in01f80 g555370 ( .a(n_14381), .o(n_14382) );
no02f80 g555371 ( .a(n_13057), .b(n_11710), .o(n_14381) );
no02f80 g555372 ( .a(n_13058), .b(n_11711), .o(n_15143) );
in01f80 g555373 ( .a(n_14379), .o(n_14380) );
na02f80 g555374 ( .a(n_13055), .b(n_11745), .o(n_14379) );
na02f80 g555375 ( .a(n_13056), .b(n_11746), .o(n_15142) );
in01f80 g555376 ( .a(n_14377), .o(n_14378) );
no02f80 g555377 ( .a(n_13053), .b(n_11708), .o(n_14377) );
no02f80 g555378 ( .a(n_13054), .b(n_11709), .o(n_15141) );
in01f80 g555379 ( .a(n_14375), .o(n_14376) );
na02f80 g555380 ( .a(n_13051), .b(n_11743), .o(n_14375) );
na02f80 g555381 ( .a(n_13052), .b(n_11744), .o(n_15140) );
in01f80 g555382 ( .a(n_14373), .o(n_14374) );
no02f80 g555383 ( .a(n_13049), .b(n_11752), .o(n_14373) );
no02f80 g555384 ( .a(n_13050), .b(n_11753), .o(n_15139) );
in01f80 g555385 ( .a(n_14371), .o(n_14372) );
na02f80 g555386 ( .a(n_13047), .b(n_9772), .o(n_14371) );
na02f80 g555387 ( .a(n_13048), .b(n_9773), .o(n_15138) );
in01f80 g555388 ( .a(n_13973), .o(n_13974) );
no02f80 g555389 ( .a(n_12592), .b(n_9722), .o(n_13973) );
in01f80 g555390 ( .a(n_14730), .o(n_14731) );
na02f80 g555391 ( .a(n_13568), .b(n_11706), .o(n_14730) );
na02f80 g555392 ( .a(n_13569), .b(n_11707), .o(n_15390) );
no02f80 g555393 ( .a(n_13642), .b(n_14729), .o(n_23874) );
na02f80 g555394 ( .a(n_14728), .b(n_13645), .o(n_16160) );
no02f80 g555395 ( .a(n_13177), .b(n_14370), .o(n_17035) );
na02f80 g555396 ( .a(n_14369), .b(n_13179), .o(n_17962) );
no02f80 g555397 ( .a(n_13182), .b(n_14368), .o(n_18914) );
na02f80 g555398 ( .a(n_13184), .b(n_14367), .o(n_19933) );
no02f80 g555399 ( .a(n_13186), .b(n_14366), .o(n_20730) );
na02f80 g555400 ( .a(n_13188), .b(n_14365), .o(n_21839) );
no02f80 g555401 ( .a(n_13190), .b(n_14364), .o(n_22779) );
na02f80 g555402 ( .a(n_14363), .b(n_13192), .o(n_23741) );
oa12f80 g555403 ( .a(FE_OFN375_n_14224), .b(n_1543), .c(FE_OFN134_n_27449), .o(n_14362) );
no02f80 g555404 ( .a(n_13194), .b(n_14361), .o(n_24743) );
oa12f80 g555405 ( .a(n_12464), .b(n_12099), .c(n_12562), .o(n_15476) );
no02f80 g555406 ( .a(n_14355), .b(n_14354), .o(n_15389) );
in01f80 g555407 ( .a(n_14359), .o(n_14360) );
no02f80 g555408 ( .a(n_13045), .b(n_10579), .o(n_14359) );
in01f80 g555409 ( .a(n_14726), .o(n_14727) );
na02f80 g555410 ( .a(n_13594), .b(n_12321), .o(n_14726) );
no02f80 g555411 ( .a(n_14358), .b(n_14357), .o(n_15407) );
na02f80 g555412 ( .a(n_13172), .b(n_14356), .o(n_23839) );
in01f80 g555413 ( .a(n_14724), .o(n_14725) );
na02f80 g555414 ( .a(n_14355), .b(n_14354), .o(n_14724) );
in01f80 g555415 ( .a(n_14352), .o(n_14353) );
na02f80 g555416 ( .a(n_13043), .b(n_10588), .o(n_14352) );
in01f80 g555417 ( .a(n_14722), .o(n_14723) );
na02f80 g555418 ( .a(n_13564), .b(n_12383), .o(n_14722) );
no02f80 g555419 ( .a(n_13046), .b(n_10578), .o(n_15136) );
oa12f80 g555420 ( .a(FE_OFN396_n_14720), .b(n_1363), .c(FE_OFN134_n_27449), .o(n_14721) );
na02f80 g555421 ( .a(n_13044), .b(n_10589), .o(n_15133) );
in01f80 g555422 ( .a(n_14350), .o(n_14351) );
no02f80 g555423 ( .a(n_13041), .b(n_10583), .o(n_14350) );
na02f80 g555424 ( .a(n_14349), .b(n_14348), .o(n_15388) );
na02f80 g555425 ( .a(n_13565), .b(n_12384), .o(n_15375) );
no02f80 g555426 ( .a(n_14341), .b(n_14340), .o(n_15373) );
no02f80 g555427 ( .a(n_13042), .b(n_10582), .o(n_15132) );
in01f80 g555428 ( .a(n_14718), .o(n_14719) );
no02f80 g555429 ( .a(n_14349), .b(n_14348), .o(n_14718) );
in01f80 g555430 ( .a(n_14346), .o(n_14347) );
na02f80 g555431 ( .a(n_13039), .b(n_10590), .o(n_14346) );
in01f80 g555432 ( .a(n_14716), .o(n_14717) );
no02f80 g555433 ( .a(n_13566), .b(n_12381), .o(n_14716) );
no02f80 g555434 ( .a(n_13567), .b(n_12382), .o(n_15387) );
in01f80 g555435 ( .a(n_14714), .o(n_14715) );
na02f80 g555436 ( .a(n_13562), .b(n_12379), .o(n_14714) );
na02f80 g555437 ( .a(n_13040), .b(n_10591), .o(n_15131) );
in01f80 g555438 ( .a(n_14344), .o(n_14345) );
no02f80 g555439 ( .a(n_13037), .b(n_10595), .o(n_14344) );
na02f80 g555440 ( .a(n_13563), .b(n_12380), .o(n_15386) );
in01f80 g555441 ( .a(n_14712), .o(n_14713) );
no02f80 g555442 ( .a(n_13560), .b(n_12377), .o(n_14712) );
no02f80 g555443 ( .a(n_13561), .b(n_12378), .o(n_15385) );
in01f80 g555444 ( .a(n_14710), .o(n_14711) );
na02f80 g555445 ( .a(n_13558), .b(n_12375), .o(n_14710) );
no02f80 g555446 ( .a(n_13038), .b(n_10594), .o(n_15130) );
in01f80 g555447 ( .a(n_14342), .o(n_14343) );
na02f80 g555448 ( .a(n_13035), .b(n_10592), .o(n_14342) );
na02f80 g555449 ( .a(n_13559), .b(n_12376), .o(n_15384) );
in01f80 g555450 ( .a(n_14708), .o(n_14709) );
no02f80 g555451 ( .a(n_13556), .b(n_12924), .o(n_14708) );
in01f80 g555452 ( .a(n_14706), .o(n_14707) );
na02f80 g555453 ( .a(n_13552), .b(n_12901), .o(n_14706) );
no02f80 g555454 ( .a(n_13557), .b(n_12925), .o(n_15383) );
in01f80 g555455 ( .a(n_14704), .o(n_14705) );
na02f80 g555456 ( .a(n_13554), .b(n_11762), .o(n_14704) );
in01f80 g555457 ( .a(n_14702), .o(n_14703) );
na02f80 g555458 ( .a(n_14341), .b(n_14340), .o(n_14702) );
na02f80 g555459 ( .a(n_13036), .b(n_10593), .o(n_15129) );
in01f80 g555460 ( .a(n_13971), .o(n_13972) );
no02f80 g555461 ( .a(n_12668), .b(n_9631), .o(n_13971) );
na02f80 g555462 ( .a(n_13555), .b(n_11763), .o(n_15382) );
no02f80 g555463 ( .a(n_14339), .b(n_14338), .o(n_15381) );
in01f80 g555464 ( .a(n_14700), .o(n_14701) );
na02f80 g555465 ( .a(n_14339), .b(n_14338), .o(n_14700) );
no02f80 g555466 ( .a(n_12669), .b(n_9630), .o(n_14946) );
na02f80 g555467 ( .a(n_13553), .b(n_12902), .o(n_15372) );
in01f80 g555468 ( .a(n_14698), .o(n_14699) );
no02f80 g555469 ( .a(n_13550), .b(n_12922), .o(n_14698) );
in01f80 g555470 ( .a(n_14696), .o(n_14697) );
na02f80 g555471 ( .a(n_13548), .b(n_12918), .o(n_14696) );
no02f80 g555472 ( .a(n_13551), .b(n_12923), .o(n_15371) );
na02f80 g555473 ( .a(n_14880), .b(n_14879), .o(n_13970) );
na02f80 g555474 ( .a(n_13422), .b(FE_OFN953_n_13421), .o(n_13423) );
na02f80 g555475 ( .a(n_13549), .b(n_12919), .o(n_15370) );
in01f80 g555476 ( .a(n_13968), .o(n_13969) );
na02f80 g555477 ( .a(n_12662), .b(n_10584), .o(n_13968) );
na02f80 g555478 ( .a(n_12663), .b(n_10585), .o(n_14945) );
oa12f80 g555479 ( .a(n_14694), .b(n_679), .c(FE_OFN89_n_27449), .o(n_14695) );
na02f80 g555480 ( .a(n_14337), .b(n_14336), .o(n_15376) );
in01f80 g555481 ( .a(n_14692), .o(n_14693) );
no02f80 g555482 ( .a(n_14337), .b(n_14336), .o(n_14692) );
in01f80 g555483 ( .a(n_14690), .o(n_14691) );
no02f80 g555484 ( .a(n_13544), .b(n_12916), .o(n_14690) );
no02f80 g555485 ( .a(n_13545), .b(n_12917), .o(n_15369) );
na02f80 g555486 ( .a(n_14335), .b(n_14334), .o(n_15368) );
in01f80 g555487 ( .a(n_14688), .o(n_14689) );
no02f80 g555488 ( .a(n_14335), .b(n_14334), .o(n_14688) );
in01f80 g555489 ( .a(n_14686), .o(n_14687) );
no02f80 g555490 ( .a(n_13542), .b(n_12914), .o(n_14686) );
no02f80 g555491 ( .a(n_13543), .b(n_12915), .o(n_15367) );
in01f80 g555492 ( .a(n_14684), .o(n_14685) );
na02f80 g555493 ( .a(n_13540), .b(n_12912), .o(n_14684) );
na02f80 g555494 ( .a(n_13541), .b(n_12913), .o(n_15366) );
in01f80 g555495 ( .a(n_14682), .o(n_14683) );
no02f80 g555496 ( .a(n_13538), .b(n_12408), .o(n_14682) );
no02f80 g555497 ( .a(n_13539), .b(n_12409), .o(n_15365) );
in01f80 g555498 ( .a(n_14680), .o(n_14681) );
na02f80 g555499 ( .a(n_13536), .b(n_11760), .o(n_14680) );
na02f80 g555500 ( .a(n_13537), .b(n_11761), .o(n_15364) );
no02f80 g555501 ( .a(n_14333), .b(n_14332), .o(n_15363) );
in01f80 g555502 ( .a(n_14678), .o(n_14679) );
na02f80 g555503 ( .a(n_14333), .b(n_14332), .o(n_14678) );
in01f80 g555504 ( .a(n_14676), .o(n_14677) );
na02f80 g555505 ( .a(n_13534), .b(FE_OFN1194_n_12908), .o(n_14676) );
na02f80 g555506 ( .a(n_13535), .b(n_12909), .o(n_15360) );
no02f80 g555507 ( .a(n_13638), .b(n_14675), .o(n_24168) );
no02f80 g555508 ( .a(n_13966), .b(n_13965), .o(n_13967) );
in01f80 g555509 ( .a(n_14673), .o(n_14674) );
no02f80 g555510 ( .a(n_13512), .b(n_9779), .o(n_14673) );
in01f80 g555511 ( .a(n_13963), .o(n_13964) );
na02f80 g555512 ( .a(n_12658), .b(n_9788), .o(n_13963) );
na02f80 g555513 ( .a(n_14877), .b(n_14876), .o(n_13962) );
na02f80 g555514 ( .a(n_12659), .b(n_9789), .o(n_14936) );
in01f80 g555515 ( .a(n_13960), .o(n_13961) );
no02f80 g555516 ( .a(n_12656), .b(n_9795), .o(n_13960) );
no02f80 g555517 ( .a(n_12657), .b(n_9794), .o(n_14934) );
in01f80 g555518 ( .a(n_13958), .o(n_13959) );
na02f80 g555519 ( .a(n_12654), .b(n_10568), .o(n_13958) );
na02f80 g555520 ( .a(n_12655), .b(n_10569), .o(n_14933) );
in01f80 g555521 ( .a(n_13956), .o(n_13957) );
no02f80 g555522 ( .a(n_12652), .b(n_10607), .o(n_13956) );
no02f80 g555523 ( .a(n_12653), .b(n_10606), .o(n_14932) );
in01f80 g555524 ( .a(n_14671), .o(n_14672) );
na02f80 g555525 ( .a(n_13530), .b(n_10567), .o(n_14671) );
na02f80 g555526 ( .a(n_13531), .b(n_10566), .o(n_15354) );
in01f80 g555527 ( .a(n_13954), .o(n_13955) );
no02f80 g555528 ( .a(n_12650), .b(n_10613), .o(n_13954) );
no02f80 g555529 ( .a(n_12651), .b(n_10614), .o(n_14931) );
in01f80 g555530 ( .a(n_14330), .o(n_14331) );
na02f80 g555531 ( .a(n_13027), .b(n_10363), .o(n_14330) );
na02f80 g555532 ( .a(n_13028), .b(n_10362), .o(n_15120) );
na02f80 g555533 ( .a(n_13946), .b(n_13945), .o(n_15089) );
no02f80 g555534 ( .a(n_13166), .b(n_14329), .o(n_22510) );
no02f80 g555535 ( .a(n_14534), .b(n_14533), .o(n_13420) );
in01f80 g555536 ( .a(n_13952), .o(n_13953) );
no02f80 g555537 ( .a(n_12648), .b(n_10611), .o(n_13952) );
no02f80 g555538 ( .a(n_12649), .b(n_10612), .o(n_14930) );
na02f80 g555539 ( .a(n_13636), .b(n_14670), .o(n_21491) );
no02f80 g555540 ( .a(n_13165), .b(n_14328), .o(n_20398) );
na02f80 g555541 ( .a(n_13162), .b(n_14327), .o(n_19590) );
no02f80 g555542 ( .a(n_13160), .b(n_14326), .o(n_18612) );
na02f80 g555543 ( .a(n_14083), .b(n_15024), .o(n_16018) );
na02f80 g555544 ( .a(n_13634), .b(n_14669), .o(n_23492) );
no02f80 g555545 ( .a(n_13950), .b(n_13949), .o(n_13951) );
in01f80 g555546 ( .a(n_13947), .o(n_13948) );
no02f80 g555547 ( .a(n_12644), .b(n_11470), .o(n_13947) );
no02f80 g555548 ( .a(n_12645), .b(n_12356), .o(n_14929) );
na02f80 g555549 ( .a(n_13595), .b(n_12322), .o(n_15355) );
na02f80 g555550 ( .a(n_13632), .b(n_14325), .o(n_25175) );
in01f80 g555551 ( .a(n_14667), .o(n_14668) );
na02f80 g555552 ( .a(n_14324), .b(n_14323), .o(n_14667) );
oa12f80 g555553 ( .a(n_14638), .b(n_419), .c(FE_OFN119_n_27449), .o(n_14666) );
na02f80 g555554 ( .a(n_13032), .b(n_11405), .o(n_15160) );
in01f80 g555555 ( .a(n_14321), .o(n_14322) );
no02f80 g555556 ( .a(n_13946), .b(n_13945), .o(n_14321) );
oa12f80 g555557 ( .a(FE_OFN393_n_14663), .b(n_1572), .c(FE_OFN355_n_4860), .o(n_14664) );
na02f80 g555558 ( .a(n_13629), .b(n_14662), .o(n_15603) );
no02f80 g555559 ( .a(n_14320), .b(n_13147), .o(n_16596) );
na02f80 g555560 ( .a(n_13149), .b(n_14319), .o(n_17461) );
no02f80 g555561 ( .a(n_14318), .b(n_13151), .o(n_18359) );
na02f80 g555562 ( .a(n_13153), .b(n_14317), .o(n_19356) );
no02f80 g555563 ( .a(n_13155), .b(n_14316), .o(n_20076) );
in01f80 g555564 ( .a(n_14660), .o(n_14661) );
na02f80 g555565 ( .a(n_14311), .b(n_14310), .o(n_14660) );
na02f80 g555566 ( .a(n_13157), .b(n_14315), .o(n_21156) );
no02f80 g555567 ( .a(n_13159), .b(n_14314), .o(n_22240) );
na02f80 g555568 ( .a(n_15023), .b(n_14087), .o(n_24442) );
in01f80 g555569 ( .a(n_14312), .o(n_14313) );
na02f80 g555570 ( .a(n_13944), .b(n_13943), .o(n_14312) );
in01f80 g555571 ( .a(n_14658), .o(n_14659) );
no02f80 g555572 ( .a(n_14311), .b(n_14310), .o(n_14658) );
in01f80 g555573 ( .a(n_14656), .o(n_14657) );
no02f80 g555574 ( .a(n_13527), .b(n_12410), .o(n_14656) );
no02f80 g555575 ( .a(n_13528), .b(n_12411), .o(n_15351) );
na02f80 g555576 ( .a(n_14309), .b(n_14308), .o(n_16270) );
oa12f80 g555577 ( .a(n_13876), .b(n_349), .c(FE_OFN101_n_27449), .o(n_13942) );
in01f80 g555578 ( .a(n_15290), .o(n_15291) );
no02f80 g555579 ( .a(n_14592), .b(n_10599), .o(n_15290) );
no02f80 g555580 ( .a(n_14593), .b(n_10598), .o(n_16032) );
in01f80 g555581 ( .a(n_14654), .o(n_14655) );
na02f80 g555582 ( .a(n_13525), .b(n_9761), .o(n_14654) );
na02f80 g555583 ( .a(n_13526), .b(n_9760), .o(n_15350) );
in01f80 g555584 ( .a(n_14306), .o(n_14307) );
no02f80 g555585 ( .a(n_13021), .b(n_11758), .o(n_14306) );
no02f80 g555586 ( .a(n_13940), .b(n_13939), .o(n_13941) );
no02f80 g555587 ( .a(n_13022), .b(n_11759), .o(n_15114) );
in01f80 g555588 ( .a(n_14304), .o(n_14305) );
na02f80 g555589 ( .a(n_13019), .b(n_9759), .o(n_14304) );
na02f80 g555590 ( .a(n_13020), .b(n_9758), .o(n_15113) );
in01f80 g555591 ( .a(n_14302), .o(n_14303) );
no02f80 g555592 ( .a(n_13017), .b(n_11411), .o(n_14302) );
no02f80 g555593 ( .a(n_13018), .b(n_11412), .o(n_15112) );
in01f80 g555594 ( .a(n_14300), .o(n_14301) );
no02f80 g555595 ( .a(n_13938), .b(n_13937), .o(n_14300) );
na02f80 g555596 ( .a(n_13935), .b(n_13934), .o(n_13936) );
na02f80 g555597 ( .a(n_13933), .b(n_13932), .o(n_15110) );
in01f80 g555598 ( .a(n_14298), .o(n_14299) );
no02f80 g555599 ( .a(n_13933), .b(n_13932), .o(n_14298) );
no02f80 g555600 ( .a(n_13597), .b(n_11090), .o(n_15413) );
in01f80 g555601 ( .a(n_14296), .o(n_14297) );
no02f80 g555602 ( .a(n_13015), .b(n_11754), .o(n_14296) );
no02f80 g555603 ( .a(n_13016), .b(n_11755), .o(n_15109) );
na02f80 g555604 ( .a(n_13138), .b(n_14295), .o(n_24881) );
na02f80 g555605 ( .a(n_13654), .b(n_14653), .o(n_15581) );
in01f80 g555606 ( .a(n_14651), .o(n_14652) );
no02f80 g555607 ( .a(n_14294), .b(n_14293), .o(n_14651) );
no02f80 g555608 ( .a(n_13221), .b(n_14292), .o(n_22245) );
na02f80 g555609 ( .a(n_13524), .b(n_12889), .o(n_19935) );
na02f80 g555610 ( .a(n_13930), .b(n_13929), .o(n_13931) );
no02f80 g555611 ( .a(n_24513), .b(n_14291), .o(n_23833) );
in01f80 g555612 ( .a(n_14289), .o(n_14290) );
no02f80 g555613 ( .a(n_13095), .b(n_13928), .o(n_14289) );
no02f80 g555614 ( .a(n_13096), .b(n_10389), .o(n_15106) );
in01f80 g555615 ( .a(n_14287), .o(n_14288) );
no02f80 g555616 ( .a(n_12964), .b(n_10359), .o(n_14287) );
oa12f80 g555617 ( .a(FE_OFN377_n_14285), .b(n_1519), .c(FE_OFN93_n_27449), .o(n_14286) );
no02f80 g555618 ( .a(n_14283), .b(n_14282), .o(n_14284) );
ao12f80 g555619 ( .a(n_12063), .b(n_13301), .c(n_10843), .o(n_14581) );
na02f80 g555620 ( .a(n_14281), .b(n_13122), .o(n_24523) );
na02f80 g555621 ( .a(n_14279), .b(n_14278), .o(n_14280) );
na02f80 g555622 ( .a(n_13875), .b(n_13874), .o(n_15117) );
no02f80 g555623 ( .a(n_13927), .b(n_13926), .o(n_15104) );
no02f80 g555624 ( .a(n_13418), .b(n_13417), .o(n_13419) );
na02f80 g555625 ( .a(n_13626), .b(n_14650), .o(n_17107) );
no02f80 g555626 ( .a(n_13131), .b(n_14277), .o(n_18034) );
na02f80 g555627 ( .a(n_14276), .b(n_13129), .o(n_19006) );
no02f80 g555628 ( .a(n_14274), .b(FE_OFN1081_n_14273), .o(n_14275) );
no02f80 g555629 ( .a(n_13127), .b(n_14272), .o(n_20018) );
na02f80 g555630 ( .a(n_13623), .b(n_14271), .o(n_20822) );
no02f80 g555631 ( .a(n_14269), .b(n_14268), .o(n_14270) );
no02f80 g555632 ( .a(n_13125), .b(n_14267), .o(n_21926) );
na02f80 g555633 ( .a(n_13621), .b(n_14266), .o(n_22875) );
no02f80 g555634 ( .a(n_13619), .b(n_14265), .o(n_23837) );
na02f80 g555635 ( .a(n_13617), .b(n_14649), .o(n_26226) );
na02f80 g555636 ( .a(n_14263), .b(n_14262), .o(n_14264) );
in01f80 g555637 ( .a(n_14260), .o(n_14261) );
na02f80 g555638 ( .a(n_13927), .b(n_13926), .o(n_14260) );
in01f80 g555639 ( .a(n_14258), .o(n_14259) );
na02f80 g555640 ( .a(n_12999), .b(n_9762), .o(n_14258) );
no02f80 g555641 ( .a(n_13399), .b(n_13398), .o(n_14908) );
oa12f80 g555642 ( .a(n_13924), .b(n_313), .c(FE_OFN353_n_4860), .o(n_13925) );
na02f80 g555643 ( .a(n_13000), .b(n_9763), .o(n_15101) );
in01f80 g555644 ( .a(n_13922), .o(n_13923) );
no02f80 g555645 ( .a(n_12622), .b(n_9757), .o(n_13922) );
no02f80 g555646 ( .a(n_12623), .b(n_9756), .o(n_14915) );
in01f80 g555647 ( .a(n_14256), .o(n_14257) );
na02f80 g555648 ( .a(n_12997), .b(n_9754), .o(n_14256) );
na02f80 g555649 ( .a(n_12998), .b(n_9755), .o(n_15179) );
in01f80 g555650 ( .a(n_14254), .o(n_14255) );
no02f80 g555651 ( .a(n_12995), .b(n_9753), .o(n_14254) );
no02f80 g555652 ( .a(n_12996), .b(n_9752), .o(n_15099) );
no02f80 g555653 ( .a(n_13415), .b(n_13414), .o(n_13416) );
in01f80 g555654 ( .a(n_14252), .o(n_14253) );
na02f80 g555655 ( .a(n_12993), .b(n_9750), .o(n_14252) );
na02f80 g555656 ( .a(n_14571), .b(n_13920), .o(n_13921) );
na02f80 g555657 ( .a(n_12994), .b(n_9751), .o(n_15095) );
in01f80 g555658 ( .a(n_14250), .o(n_14251) );
no02f80 g555659 ( .a(n_13088), .b(n_12330), .o(n_14250) );
no02f80 g555660 ( .a(n_13089), .b(n_12331), .o(n_15098) );
no02f80 g555661 ( .a(n_13217), .b(n_14249), .o(n_20080) );
na02f80 g555662 ( .a(n_13919), .b(n_13918), .o(n_15174) );
no02f80 g555663 ( .a(n_14648), .b(n_14647), .o(n_16243) );
in01f80 g555664 ( .a(n_15021), .o(n_15691) );
na02f80 g555665 ( .a(n_14648), .b(n_14647), .o(n_15021) );
in01f80 g555666 ( .a(n_13916), .o(n_13917) );
na02f80 g555667 ( .a(n_12620), .b(n_9766), .o(n_13916) );
na02f80 g555668 ( .a(n_12621), .b(n_9767), .o(n_14914) );
in01f80 g555669 ( .a(n_13915), .o(n_14964) );
no02f80 g555670 ( .a(n_13413), .b(n_13412), .o(n_13915) );
na02f80 g555671 ( .a(n_13517), .b(n_12428), .o(n_15347) );
na02f80 g555672 ( .a(n_13913), .b(n_13912), .o(n_13914) );
na02f80 g555673 ( .a(n_13910), .b(n_13909), .o(n_13911) );
na02f80 g555674 ( .a(n_13907), .b(n_13906), .o(n_13908) );
na02f80 g555675 ( .a(n_13410), .b(n_13409), .o(n_13411) );
na02f80 g555676 ( .a(n_13615), .b(n_14646), .o(n_20457) );
in01f80 g555677 ( .a(n_13904), .o(n_13905) );
no02f80 g555678 ( .a(n_12660), .b(n_9717), .o(n_13904) );
no02f80 g555679 ( .a(n_12661), .b(n_9716), .o(n_14913) );
in01f80 g555680 ( .a(n_13902), .o(n_13903) );
na02f80 g555681 ( .a(n_12611), .b(n_9729), .o(n_13902) );
na02f80 g555682 ( .a(n_12612), .b(n_9730), .o(n_14912) );
in01f80 g555683 ( .a(n_13900), .o(n_13901) );
no02f80 g555684 ( .a(n_12609), .b(n_10573), .o(n_13900) );
no02f80 g555685 ( .a(n_12610), .b(n_10572), .o(n_14911) );
in01f80 g555686 ( .a(n_13898), .o(n_13899) );
na02f80 g555687 ( .a(n_12607), .b(n_9727), .o(n_13898) );
na02f80 g555688 ( .a(n_12608), .b(n_9728), .o(n_14910) );
in01f80 g555689 ( .a(n_14247), .o(n_14248) );
no02f80 g555690 ( .a(n_13075), .b(n_9736), .o(n_14247) );
no02f80 g555691 ( .a(n_13076), .b(n_9735), .o(n_15094) );
in01f80 g555692 ( .a(n_14245), .o(n_14246) );
na02f80 g555693 ( .a(n_12987), .b(n_9725), .o(n_14245) );
na02f80 g555694 ( .a(n_13896), .b(n_13895), .o(n_13897) );
na02f80 g555695 ( .a(n_12988), .b(n_9726), .o(n_15093) );
in01f80 g555696 ( .a(n_14243), .o(n_14244) );
no02f80 g555697 ( .a(n_12985), .b(n_12325), .o(n_14243) );
no02f80 g555698 ( .a(n_12986), .b(n_12326), .o(n_15092) );
na02f80 g555699 ( .a(n_13612), .b(n_14645), .o(n_23574) );
na02f80 g555700 ( .a(n_14856), .b(n_14855), .o(n_13894) );
in01f80 g555701 ( .a(n_13892), .o(n_13893) );
na02f80 g555702 ( .a(n_12603), .b(n_9743), .o(n_13892) );
na02f80 g555703 ( .a(n_12604), .b(n_9744), .o(n_14909) );
no02f80 g555704 ( .a(n_13034), .b(n_11068), .o(n_15161) );
no02f80 g555705 ( .a(n_13407), .b(n_13406), .o(n_13408) );
no02f80 g555706 ( .a(n_13593), .b(n_12387), .o(n_15418) );
na02f80 g555707 ( .a(n_13890), .b(n_13889), .o(n_13891) );
na02f80 g555708 ( .a(n_12992), .b(n_11732), .o(n_15164) );
na02f80 g555709 ( .a(n_14241), .b(n_14240), .o(n_14242) );
na02f80 g555710 ( .a(n_14238), .b(n_14237), .o(n_14239) );
in01f80 g555711 ( .a(n_14643), .o(n_14644) );
no02f80 g555712 ( .a(n_13518), .b(n_12247), .o(n_14643) );
no02f80 g555713 ( .a(n_13519), .b(n_12248), .o(n_15374) );
no02f80 g555714 ( .a(n_13404), .b(n_13403), .o(n_13405) );
na02f80 g555715 ( .a(n_13401), .b(n_13400), .o(n_13402) );
no02f80 g555716 ( .a(n_13887), .b(n_13886), .o(n_13888) );
in01f80 g555717 ( .a(n_14641), .o(n_14642) );
no02f80 g555718 ( .a(n_14236), .b(n_14235), .o(n_14641) );
in01f80 g555719 ( .a(n_13884), .o(n_13885) );
na02f80 g555720 ( .a(n_13399), .b(n_13398), .o(n_13884) );
in01f80 g555721 ( .a(n_13882), .o(n_13883) );
na02f80 g555722 ( .a(n_12594), .b(n_9723), .o(n_13882) );
na02f80 g555723 ( .a(n_12595), .b(n_9724), .o(n_14907) );
no02f80 g555724 ( .a(n_12593), .b(n_9721), .o(n_14906) );
in01f80 g555725 ( .a(n_13880), .o(n_13881) );
na02f80 g555726 ( .a(n_12590), .b(n_11408), .o(n_13880) );
na02f80 g555727 ( .a(n_12591), .b(n_11407), .o(n_14941) );
in01f80 g555728 ( .a(n_13878), .o(n_13879) );
no02f80 g555729 ( .a(n_12588), .b(n_9732), .o(n_13878) );
no02f80 g555730 ( .a(n_12589), .b(n_9731), .o(n_14925) );
in01f80 g555731 ( .a(n_14233), .o(n_14234) );
na02f80 g555732 ( .a(n_12973), .b(n_9739), .o(n_14233) );
na02f80 g555733 ( .a(n_12974), .b(n_9740), .o(n_15172) );
in01f80 g555734 ( .a(n_14231), .o(n_14232) );
no02f80 g555735 ( .a(n_12971), .b(n_12319), .o(n_14231) );
oa12f80 g555736 ( .a(n_13876), .b(n_1124), .c(FE_OFN101_n_27449), .o(n_13877) );
no02f80 g555737 ( .a(n_12972), .b(n_12320), .o(n_15105) );
in01f80 g555738 ( .a(n_14229), .o(n_14230) );
no02f80 g555739 ( .a(n_13875), .b(n_13874), .o(n_14229) );
in01f80 g555740 ( .a(n_13872), .o(n_13873) );
na02f80 g555741 ( .a(n_12584), .b(n_9741), .o(n_13872) );
na02f80 g555742 ( .a(n_12585), .b(n_9742), .o(n_14905) );
na02f80 g555743 ( .a(n_13870), .b(n_13869), .o(n_13871) );
no02f80 g555744 ( .a(n_13581), .b(n_12407), .o(n_15405) );
in01f80 g555745 ( .a(n_13867), .o(n_13868) );
na02f80 g555746 ( .a(n_12573), .b(n_9733), .o(n_13867) );
no02f80 g555747 ( .a(n_14227), .b(n_14226), .o(n_14228) );
na02f80 g555748 ( .a(n_13611), .b(n_14640), .o(n_20461) );
oa12f80 g555749 ( .a(FE_OFN375_n_14224), .b(n_678), .c(FE_OFN134_n_27449), .o(n_14225) );
na02f80 g555750 ( .a(n_13865), .b(n_13864), .o(n_13866) );
in01f80 g555751 ( .a(n_14222), .o(n_14223) );
na02f80 g555752 ( .a(n_13863), .b(n_13862), .o(n_14222) );
na02f80 g555753 ( .a(n_14220), .b(n_14219), .o(n_14221) );
oa12f80 g555754 ( .a(n_14638), .b(n_578), .c(FE_OFN1111_rst), .o(n_14639) );
no02f80 g555755 ( .a(n_13397), .b(n_13396), .o(n_14917) );
in01f80 g555756 ( .a(n_14217), .o(n_14218) );
na02f80 g555757 ( .a(n_12966), .b(n_10563), .o(n_14217) );
na02f80 g555758 ( .a(n_12967), .b(n_10562), .o(n_15116) );
no02f80 g555759 ( .a(n_13860), .b(n_13859), .o(n_13861) );
no02f80 g555760 ( .a(n_12965), .b(n_10358), .o(n_15084) );
in01f80 g555761 ( .a(n_14215), .o(n_14216) );
na02f80 g555762 ( .a(n_12962), .b(n_10602), .o(n_14215) );
in01f80 g555763 ( .a(n_14636), .o(n_14637) );
no02f80 g555764 ( .a(n_14214), .b(n_14213), .o(n_14636) );
in01f80 g555765 ( .a(n_14634), .o(n_14635) );
na02f80 g555766 ( .a(n_14212), .b(n_14211), .o(n_14634) );
na02f80 g555767 ( .a(n_12963), .b(n_10603), .o(n_15086) );
no02f80 g555768 ( .a(n_13394), .b(n_13393), .o(n_13395) );
no02f80 g555769 ( .a(n_13513), .b(n_9778), .o(n_15348) );
na02f80 g555770 ( .a(n_12574), .b(n_9734), .o(n_14918) );
in01f80 g555771 ( .a(n_13857), .o(n_13858) );
na02f80 g555772 ( .a(n_13392), .b(n_13391), .o(n_13857) );
na02f80 g555773 ( .a(n_13390), .b(n_13389), .o(n_16234) );
in01f80 g555774 ( .a(n_18500), .o(n_14210) );
oa12f80 g555775 ( .a(n_13746), .b(n_12538), .c(n_11749), .o(n_18500) );
in01f80 g555776 ( .a(n_13856), .o(n_14919) );
no02f80 g555777 ( .a(n_13390), .b(n_13389), .o(n_13856) );
na02f80 g555778 ( .a(n_14882), .b(n_14881), .o(n_13855) );
oa12f80 g555779 ( .a(n_13853), .b(n_1188), .c(FE_OFN134_n_27449), .o(n_13854) );
in01f80 g555780 ( .a(n_13388), .o(n_14976) );
oa12f80 g555781 ( .a(n_3271), .b(n_12858), .c(n_2181), .o(n_13388) );
oa12f80 g555782 ( .a(n_13853), .b(n_452), .c(FE_OFN134_n_27449), .o(n_13852) );
in01f80 g555783 ( .a(n_13851), .o(n_15194) );
oa12f80 g555784 ( .a(n_10969), .b(n_13366), .c(n_9201), .o(n_13851) );
in01f80 g555785 ( .a(n_13387), .o(n_14974) );
oa12f80 g555786 ( .a(n_2704), .b(n_12856), .c(n_2188), .o(n_13387) );
in01f80 g555787 ( .a(n_13850), .o(n_15196) );
oa12f80 g555788 ( .a(n_10996), .b(n_13370), .c(n_9197), .o(n_13850) );
oa12f80 g555789 ( .a(n_14632), .b(n_3), .c(FE_OFN116_n_27449), .o(n_14633) );
oa12f80 g555790 ( .a(n_14630), .b(n_1490), .c(FE_OFN1112_rst), .o(n_14631) );
oa12f80 g555791 ( .a(n_14628), .b(n_1248), .c(FE_OFN1106_rst), .o(n_14629) );
oa12f80 g555792 ( .a(n_14208), .b(n_50), .c(FE_OFN358_n_4860), .o(n_14209) );
oa12f80 g555793 ( .a(n_13224), .b(n_225), .c(FE_OFN113_n_27449), .o(n_13849) );
oa12f80 g555794 ( .a(n_14208), .b(n_1066), .c(FE_OFN77_n_27012), .o(n_14207) );
oa12f80 g555795 ( .a(n_14632), .b(n_591), .c(FE_OFN1143_n_27012), .o(n_14627) );
oa12f80 g555796 ( .a(n_14628), .b(n_593), .c(FE_OFN324_n_4860), .o(n_14626) );
oa12f80 g555797 ( .a(n_14624), .b(n_861), .c(FE_OFN134_n_27449), .o(n_14625) );
oa12f80 g555798 ( .a(n_14630), .b(n_295), .c(n_29261), .o(n_14623) );
oa12f80 g555799 ( .a(n_14624), .b(n_206), .c(FE_OFN1174_n_4860), .o(n_14622) );
oa22f80 g555800 ( .a(n_12850), .b(n_11501), .c(n_12849), .d(n_11102), .o(n_14588) );
oa12f80 g555801 ( .a(FE_OFN548_n_10452), .b(n_11377), .c(n_6372), .o(n_13489) );
ao12f80 g555802 ( .a(n_3869), .b(n_12242), .c(n_6443), .o(n_14079) );
oa12f80 g555803 ( .a(n_10151), .b(n_13257), .c(n_10152), .o(n_13848) );
oa22f80 g555804 ( .a(n_12848), .b(n_11538), .c(n_12847), .d(n_11101), .o(n_14589) );
oa12f80 g555805 ( .a(n_9559), .b(n_13377), .c(n_8388), .o(n_14978) );
in01f80 g555806 ( .a(n_13846), .o(n_13847) );
ao22s80 g555807 ( .a(n_13386), .b(n_7931), .c(n_8845), .d(n_9302), .o(n_13846) );
in01f80 g555808 ( .a(FE_OFN690_n_16216), .o(n_14206) );
ao22s80 g555809 ( .a(n_13278), .b(n_8829), .c(n_11769), .d(n_13277), .o(n_16216) );
in01f80 g555810 ( .a(FE_OFN895_n_15923), .o(n_13845) );
ao22s80 g555811 ( .a(n_12835), .b(n_8363), .c(n_11078), .d(n_12834), .o(n_15923) );
oa12f80 g555812 ( .a(n_12082), .b(n_14502), .c(n_13258), .o(n_15200) );
in01f80 g555813 ( .a(n_13843), .o(n_13844) );
ao22s80 g555814 ( .a(n_11357), .b(n_12636), .c(n_14037), .d(n_12635), .o(n_13843) );
in01f80 g555815 ( .a(n_13841), .o(n_13842) );
ao22s80 g555816 ( .a(n_11358), .b(n_12633), .c(n_14034), .d(n_12634), .o(n_13841) );
ao12f80 g555817 ( .a(n_14621), .b(n_11301), .c(n_11300), .o(n_15654) );
ao22s80 g555818 ( .a(n_13385), .b(n_7881), .c(n_8849), .d(n_8848), .o(n_15530) );
oa22f80 g555819 ( .a(n_11322), .b(n_13895), .c(n_12605), .d(n_12606), .o(n_14563) );
in01f80 g555820 ( .a(n_13839), .o(n_13840) );
oa22f80 g555821 ( .a(n_11299), .b(n_13934), .c(n_12630), .d(x_in_33_5), .o(n_13839) );
oa22f80 g555822 ( .a(n_14595), .b(n_3208), .c(n_14596), .d(x_in_39_12), .o(n_14620) );
in01f80 g555823 ( .a(n_13837), .o(n_13838) );
oa22f80 g555824 ( .a(n_13384), .b(n_7004), .c(n_8450), .d(n_8449), .o(n_13837) );
oa12f80 g555825 ( .a(n_12703), .b(n_12647), .c(n_12646), .o(n_14927) );
in01f80 g555826 ( .a(n_13835), .o(n_13836) );
oa22f80 g555827 ( .a(n_13383), .b(n_6466), .c(n_8446), .d(n_8445), .o(n_13835) );
in01f80 g555828 ( .a(n_13833), .o(n_13834) );
oa22f80 g555829 ( .a(n_13382), .b(n_6972), .c(n_8505), .d(n_8504), .o(n_13833) );
oa22f80 g555830 ( .a(n_13381), .b(n_6965), .c(n_8507), .d(n_8506), .o(n_15487) );
in01f80 g555831 ( .a(n_13831), .o(n_13832) );
oa22f80 g555832 ( .a(n_13380), .b(n_6949), .c(n_8487), .d(n_8486), .o(n_13831) );
oa22f80 g555833 ( .a(n_11219), .b(n_13912), .c(n_12642), .d(n_12643), .o(n_14575) );
in01f80 g555834 ( .a(n_14204), .o(n_14205) );
ao12f80 g555835 ( .a(n_12702), .b(n_12617), .c(n_12616), .o(n_14204) );
in01f80 g555836 ( .a(n_14202), .o(n_14203) );
ao22s80 g555837 ( .a(n_12059), .b(n_13993), .c(n_12695), .d(n_12696), .o(n_14202) );
oa12f80 g555838 ( .a(n_12701), .b(n_12671), .c(n_12670), .o(n_14952) );
in01f80 g555839 ( .a(n_16696), .o(n_14619) );
oa12f80 g555840 ( .a(n_14201), .b(n_14200), .c(n_14146), .o(n_16696) );
in01f80 g555841 ( .a(n_16906), .o(n_14199) );
oa12f80 g555842 ( .a(n_11054), .b(n_13830), .c(n_11053), .o(n_16906) );
oa12f80 g555843 ( .a(n_14618), .b(n_14617), .c(n_13007), .o(n_15754) );
in01f80 g555844 ( .a(n_14197), .o(n_14198) );
ao12f80 g555845 ( .a(n_12700), .b(n_12583), .c(n_12582), .o(n_14197) );
in01f80 g555846 ( .a(n_14195), .o(n_14196) );
ao12f80 g555847 ( .a(n_12699), .b(n_12600), .c(n_12599), .o(n_14195) );
in01f80 g555848 ( .a(n_13828), .o(n_13829) );
ao22s80 g555849 ( .a(n_11203), .b(n_13450), .c(n_12196), .d(n_12197), .o(n_13828) );
in01f80 g555850 ( .a(n_14193), .o(n_14194) );
oa12f80 g555851 ( .a(n_12698), .b(n_12597), .c(n_12596), .o(n_14193) );
in01f80 g555852 ( .a(n_13826), .o(n_13827) );
oa22f80 g555853 ( .a(n_11197), .b(n_14011), .c(n_12687), .d(n_12688), .o(n_13826) );
no02f80 g555854 ( .a(n_12816), .b(n_14942), .o(n_13825) );
in01f80 g555855 ( .a(n_13823), .o(n_13824) );
ao22s80 g555856 ( .a(n_13379), .b(n_7725), .c(n_8520), .d(n_8519), .o(n_13823) );
in01f80 g555857 ( .a(n_13821), .o(n_13822) );
oa12f80 g555858 ( .a(n_12216), .b(n_12198), .c(n_10226), .o(n_13821) );
in01f80 g555859 ( .a(n_13378), .o(n_14587) );
ao22s80 g555860 ( .a(n_12239), .b(n_10860), .c(n_12238), .d(n_10165), .o(n_13378) );
ao12f80 g555861 ( .a(n_12215), .b(n_12205), .c(n_10220), .o(n_15206) );
in01f80 g555862 ( .a(n_13819), .o(n_13820) );
ao12f80 g555863 ( .a(n_12214), .b(n_12199), .c(n_10216), .o(n_13819) );
in01f80 g555864 ( .a(n_13817), .o(n_13818) );
oa12f80 g555865 ( .a(n_12213), .b(n_12194), .c(n_10212), .o(n_13817) );
in01f80 g555866 ( .a(FE_OFN1029_n_14570), .o(n_14967) );
ao22s80 g555867 ( .a(n_11073), .b(n_10346), .c(n_13377), .d(n_10347), .o(n_14570) );
in01f80 g555868 ( .a(n_14191), .o(n_14192) );
oa12f80 g555869 ( .a(n_12694), .b(n_13094), .c(n_13093), .o(n_14191) );
in01f80 g555870 ( .a(n_14189), .o(n_14190) );
oa12f80 g555871 ( .a(n_12728), .b(n_12727), .c(n_12726), .o(n_14189) );
in01f80 g555872 ( .a(n_15667), .o(n_15998) );
ao12f80 g555873 ( .a(n_13733), .b(n_13732), .c(n_13731), .o(n_15667) );
in01f80 g555874 ( .a(n_16105), .o(n_15020) );
oa12f80 g555875 ( .a(n_13696), .b(n_13695), .c(n_13694), .o(n_16105) );
in01f80 g555876 ( .a(n_17172), .o(n_15019) );
oa12f80 g555877 ( .a(n_13699), .b(n_13698), .c(n_13697), .o(n_17172) );
ao12f80 g555878 ( .a(n_13250), .b(n_13249), .c(n_15228), .o(n_14188) );
in01f80 g555879 ( .a(n_15769), .o(n_14616) );
oa12f80 g555880 ( .a(n_13349), .b(n_13348), .c(n_13347), .o(n_15769) );
in01f80 g555881 ( .a(n_13815), .o(n_13816) );
ao12f80 g555882 ( .a(n_12207), .b(n_12185), .c(FE_OFN480_n_12184), .o(n_13815) );
in01f80 g555883 ( .a(n_13813), .o(n_13814) );
oa22f80 g555884 ( .a(n_11172), .b(n_14003), .c(n_12682), .d(n_12683), .o(n_13813) );
oa22f80 g555885 ( .a(n_11169), .b(n_13441), .c(n_12191), .d(n_8502), .o(n_15218) );
in01f80 g555886 ( .a(n_13811), .o(n_13812) );
oa12f80 g555887 ( .a(n_12206), .b(n_12202), .c(FE_OFN1186_n_12201), .o(n_13811) );
in01f80 g555888 ( .a(n_14186), .o(n_14187) );
oa12f80 g555889 ( .a(n_12689), .b(n_9601), .c(FE_OFN1272_n_9600), .o(n_14186) );
ao12f80 g555890 ( .a(n_13083), .b(n_13085), .c(n_13084), .o(n_15177) );
ao12f80 g555891 ( .a(n_12753), .b(n_12752), .c(n_12751), .o(n_15176) );
oa22f80 g555892 ( .a(n_11149), .b(FE_OFN953_n_13421), .c(n_12200), .d(n_8503), .o(n_15216) );
in01f80 g555893 ( .a(n_14614), .o(n_14615) );
ao12f80 g555894 ( .a(n_12981), .b(n_13030), .c(n_13029), .o(n_14614) );
in01f80 g555895 ( .a(n_13809), .o(n_13810) );
ao12f80 g555896 ( .a(n_12208), .b(n_12146), .c(n_12147), .o(n_13809) );
ao12f80 g555897 ( .a(n_13253), .b(n_13252), .c(n_13251), .o(n_14185) );
in01f80 g555898 ( .a(n_15430), .o(n_16066) );
oa12f80 g555899 ( .a(n_13758), .b(n_13757), .c(n_13756), .o(n_15430) );
in01f80 g555900 ( .a(n_14183), .o(n_14184) );
ao12f80 g555901 ( .a(n_12813), .b(n_12812), .c(n_12811), .o(n_14183) );
in01f80 g555902 ( .a(n_13807), .o(n_13808) );
oa12f80 g555903 ( .a(n_12234), .b(n_12233), .c(n_13376), .o(n_13807) );
in01f80 g555904 ( .a(n_14181), .o(n_14182) );
oa12f80 g555905 ( .a(n_12713), .b(n_13381), .c(n_12712), .o(n_14181) );
in01f80 g555906 ( .a(n_15989), .o(n_15429) );
ao12f80 g555907 ( .a(n_13295), .b(n_13294), .c(n_13293), .o(n_15989) );
in01f80 g555908 ( .a(n_14179), .o(n_14180) );
oa22f80 g555909 ( .a(n_11795), .b(n_10146), .c(n_13376), .d(n_10147), .o(n_14179) );
oa12f80 g555910 ( .a(n_12190), .b(n_12187), .c(FE_OFN1254_n_12186), .o(n_14568) );
oa12f80 g555911 ( .a(n_12232), .b(n_12231), .c(n_13375), .o(n_14569) );
in01f80 g555912 ( .a(n_14177), .o(n_14178) );
oa22f80 g555913 ( .a(n_12000), .b(n_10143), .c(n_13375), .d(n_10144), .o(n_14177) );
ao12f80 g555914 ( .a(n_13137), .b(n_13136), .c(FE_OFN817_n_13135), .o(n_14176) );
oa22f80 g555915 ( .a(n_10209), .b(n_13409), .c(n_12203), .d(n_12204), .o(n_15547) );
in01f80 g555916 ( .a(n_15718), .o(n_15648) );
ao12f80 g555917 ( .a(n_13337), .b(n_13336), .c(n_13335), .o(n_15718) );
in01f80 g555918 ( .a(n_15018), .o(n_16035) );
oa12f80 g555919 ( .a(n_13727), .b(n_13726), .c(n_13725), .o(n_15018) );
in01f80 g555920 ( .a(n_13805), .o(n_13806) );
oa12f80 g555921 ( .a(n_12236), .b(n_12235), .c(FE_OFN989_n_13374), .o(n_13805) );
in01f80 g555922 ( .a(n_14174), .o(n_14175) );
oa22f80 g555923 ( .a(n_11990), .b(n_10140), .c(FE_OFN989_n_13374), .d(n_10141), .o(n_14174) );
in01f80 g555924 ( .a(n_15721), .o(n_15341) );
ao12f80 g555925 ( .a(n_13346), .b(n_13345), .c(n_13344), .o(n_15721) );
ao22s80 g555926 ( .a(n_12858), .b(n_3703), .c(n_10173), .d(n_3702), .o(n_12859) );
in01f80 g555927 ( .a(n_15725), .o(n_15286) );
ao12f80 g555928 ( .a(n_13340), .b(n_13339), .c(n_13338), .o(n_15725) );
in01f80 g555929 ( .a(n_14172), .o(n_14173) );
ao12f80 g555930 ( .a(n_12802), .b(n_12801), .c(FE_OFN572_n_12800), .o(n_14172) );
in01f80 g555931 ( .a(n_13803), .o(n_13804) );
oa12f80 g555932 ( .a(n_12230), .b(n_12229), .c(n_13373), .o(n_13803) );
in01f80 g555933 ( .a(n_14170), .o(n_14171) );
oa22f80 g555934 ( .a(n_11967), .b(FE_OFN574_n_10137), .c(n_13373), .d(n_10138), .o(n_14170) );
in01f80 g555935 ( .a(n_15352), .o(n_16361) );
oa12f80 g555936 ( .a(n_13684), .b(n_13683), .c(n_13682), .o(n_15352) );
in01f80 g555937 ( .a(n_14168), .o(n_14169) );
oa12f80 g555938 ( .a(n_12792), .b(n_13386), .c(n_12791), .o(n_14168) );
in01f80 g555939 ( .a(n_15733), .o(n_15673) );
ao12f80 g555940 ( .a(n_13333), .b(n_13332), .c(n_13331), .o(n_15733) );
in01f80 g555941 ( .a(n_14166), .o(n_14167) );
ao12f80 g555942 ( .a(n_12789), .b(n_12788), .c(n_12787), .o(n_14166) );
in01f80 g555943 ( .a(n_13801), .o(n_13802) );
oa12f80 g555944 ( .a(n_12228), .b(n_12227), .c(n_13372), .o(n_13801) );
in01f80 g555945 ( .a(n_14164), .o(n_14165) );
oa22f80 g555946 ( .a(n_11942), .b(n_10134), .c(n_13372), .d(n_10135), .o(n_14164) );
in01f80 g555947 ( .a(n_14935), .o(n_15730) );
oa12f80 g555948 ( .a(n_12853), .b(n_12852), .c(n_12851), .o(n_14935) );
in01f80 g555949 ( .a(n_15707), .o(n_15284) );
ao12f80 g555950 ( .a(n_14105), .b(n_14104), .c(n_14103), .o(n_15707) );
in01f80 g555951 ( .a(n_15185), .o(n_14613) );
ao12f80 g555952 ( .a(n_13284), .b(n_13283), .c(n_13282), .o(n_15185) );
oa12f80 g555953 ( .a(n_14117), .b(n_14116), .c(n_14115), .o(n_16003) );
in01f80 g555954 ( .a(n_16008), .o(n_16415) );
ao12f80 g555955 ( .a(n_13749), .b(n_13748), .c(n_13747), .o(n_16008) );
in01f80 g555956 ( .a(n_14162), .o(n_14163) );
ao12f80 g555957 ( .a(n_12686), .b(n_12691), .c(n_12690), .o(n_14162) );
ao22s80 g555958 ( .a(n_13370), .b(n_11620), .c(n_11077), .d(n_11619), .o(n_13371) );
in01f80 g555959 ( .a(n_15726), .o(n_15642) );
ao12f80 g555960 ( .a(n_13324), .b(n_13323), .c(n_13322), .o(n_15726) );
in01f80 g555961 ( .a(n_14160), .o(n_14161) );
ao12f80 g555962 ( .a(n_12763), .b(n_12762), .c(FE_OFN1216_n_12761), .o(n_14160) );
in01f80 g555963 ( .a(n_13799), .o(n_13800) );
oa12f80 g555964 ( .a(n_12226), .b(n_12225), .c(FE_OFN1218_n_13369), .o(n_13799) );
in01f80 g555965 ( .a(n_14158), .o(n_14159) );
oa22f80 g555966 ( .a(n_11899), .b(n_11032), .c(FE_OFN1218_n_13369), .d(n_11033), .o(n_14158) );
in01f80 g555967 ( .a(n_16048), .o(n_15695) );
ao12f80 g555968 ( .a(n_13705), .b(n_13704), .c(n_13703), .o(n_16048) );
in01f80 g555969 ( .a(n_14156), .o(n_14157) );
ao12f80 g555970 ( .a(n_12760), .b(n_13380), .c(n_12759), .o(n_14156) );
oa12f80 g555971 ( .a(n_12818), .b(n_13798), .c(n_12817), .o(n_14943) );
in01f80 g555972 ( .a(n_15727), .o(n_15288) );
ao12f80 g555973 ( .a(n_13319), .b(n_13318), .c(n_13317), .o(n_15727) );
in01f80 g555974 ( .a(n_14154), .o(n_14155) );
ao12f80 g555975 ( .a(n_12756), .b(n_12755), .c(FE_OFN1276_n_12754), .o(n_14154) );
in01f80 g555976 ( .a(n_15679), .o(n_15663) );
ao12f80 g555977 ( .a(n_13316), .b(n_13315), .c(n_13314), .o(n_15679) );
in01f80 g555978 ( .a(n_13796), .o(n_13797) );
oa12f80 g555979 ( .a(n_12224), .b(n_12223), .c(n_13368), .o(n_13796) );
in01f80 g555980 ( .a(n_14152), .o(n_14153) );
oa22f80 g555981 ( .a(n_11869), .b(n_11029), .c(n_13368), .d(n_11030), .o(n_14152) );
oa12f80 g555982 ( .a(n_14114), .b(n_14113), .c(n_14112), .o(n_16001) );
oa12f80 g555983 ( .a(n_13266), .b(n_13265), .c(x_in_1_9), .o(n_15267) );
ao22s80 g555984 ( .a(n_13366), .b(n_11608), .c(n_11079), .d(n_11607), .o(n_13367) );
in01f80 g555985 ( .a(n_13364), .o(n_13365) );
oa22f80 g555986 ( .a(n_10200), .b(n_13453), .c(n_12153), .d(n_12152), .o(n_13364) );
in01f80 g555987 ( .a(n_13761), .o(n_13786) );
ao12f80 g555988 ( .a(n_10326), .b(n_11377), .c(n_10325), .o(n_13761) );
in01f80 g555989 ( .a(n_15807), .o(n_15017) );
oa12f80 g555990 ( .a(n_13721), .b(n_13720), .c(n_13719), .o(n_15807) );
in01f80 g555991 ( .a(n_16042), .o(n_15697) );
ao12f80 g555992 ( .a(n_13740), .b(n_13739), .c(n_13738), .o(n_16042) );
in01f80 g555993 ( .a(n_14150), .o(n_14151) );
oa12f80 g555994 ( .a(n_12748), .b(n_13379), .c(n_12747), .o(n_14150) );
in01f80 g555995 ( .a(n_15008), .o(n_14612) );
ao12f80 g555996 ( .a(n_13234), .b(n_13233), .c(n_13232), .o(n_15008) );
in01f80 g555997 ( .a(n_14148), .o(n_14149) );
ao12f80 g555998 ( .a(n_12681), .b(n_9623), .c(n_9622), .o(n_14148) );
ao22s80 g555999 ( .a(n_12856), .b(n_4067), .c(n_10174), .d(n_4066), .o(n_12857) );
oa12f80 g556000 ( .a(n_13706), .b(n_13760), .c(n_14102), .o(n_15282) );
oa12f80 g556001 ( .a(n_13245), .b(n_13244), .c(n_13243), .o(n_15242) );
ao22s80 g556002 ( .a(n_13830), .b(n_12312), .c(n_12896), .d(x_in_8_1), .o(n_15229) );
in01f80 g556003 ( .a(n_17170), .o(n_15283) );
oa12f80 g556004 ( .a(n_14099), .b(n_14098), .c(n_14097), .o(n_17170) );
in01f80 g556005 ( .a(n_15715), .o(n_15885) );
ao12f80 g556006 ( .a(n_13715), .b(n_13714), .c(n_13713), .o(n_15715) );
in01f80 g556007 ( .a(n_16675), .o(n_15016) );
oa12f80 g556008 ( .a(n_13724), .b(n_13723), .c(n_13722), .o(n_16675) );
in01f80 g556009 ( .a(n_15819), .o(n_14611) );
oa12f80 g556010 ( .a(n_13240), .b(n_13239), .c(n_14147), .o(n_15819) );
ao22s80 g556011 ( .a(n_11242), .b(n_13478), .c(n_12177), .d(n_12178), .o(n_15527) );
in01f80 g556012 ( .a(n_13794), .o(n_13795) );
oa12f80 g556013 ( .a(n_12219), .b(n_12176), .c(x_in_33_9), .o(n_13794) );
in01f80 g556014 ( .a(n_13792), .o(n_13793) );
ao22s80 g556015 ( .a(n_11251), .b(n_13472), .c(n_12174), .d(n_12175), .o(n_13792) );
in01f80 g556016 ( .a(n_13790), .o(n_13791) );
oa12f80 g556017 ( .a(n_12220), .b(n_12173), .c(x_in_33_7), .o(n_13790) );
in01f80 g556018 ( .a(n_13788), .o(n_13789) );
ao22s80 g556019 ( .a(n_11249), .b(n_13481), .c(n_12171), .d(n_12172), .o(n_13788) );
in01f80 g556020 ( .a(n_15889), .o(n_15890) );
oa12f80 g556021 ( .a(n_13264), .b(n_13263), .c(n_13262), .o(n_15889) );
ao12f80 g556022 ( .a(n_13142), .b(n_13141), .c(n_13140), .o(n_21790) );
oa12f80 g556023 ( .a(n_13281), .b(n_13280), .c(n_13279), .o(n_16686) );
in01f80 g556024 ( .a(n_14076), .o(n_14566) );
ao22s80 g556025 ( .a(n_10164), .b(n_6469), .c(n_12242), .d(n_6468), .o(n_14076) );
in01f80 g556026 ( .a(n_13784), .o(n_13785) );
oa12f80 g556027 ( .a(n_12218), .b(n_12183), .c(n_12697), .o(n_13784) );
in01f80 g556028 ( .a(n_14609), .o(n_14610) );
oa12f80 g556029 ( .a(n_13092), .b(n_13091), .c(FE_OFN1190_n_13090), .o(n_14609) );
in01f80 g556030 ( .a(n_14608), .o(n_15436) );
ao12f80 g556031 ( .a(n_13238), .b(n_13237), .c(n_14147), .o(n_14608) );
in01f80 g556032 ( .a(n_14606), .o(n_14607) );
oa12f80 g556033 ( .a(n_13006), .b(n_13004), .c(FE_OFN1198_n_13003), .o(n_14606) );
in01f80 g556034 ( .a(n_15273), .o(n_15660) );
ao12f80 g556035 ( .a(n_13303), .b(n_13302), .c(n_13301), .o(n_15273) );
in01f80 g556036 ( .a(n_14604), .o(n_14605) );
ao12f80 g556037 ( .a(n_13005), .b(n_13002), .c(n_13001), .o(n_14604) );
in01f80 g556038 ( .a(n_13362), .o(n_13363) );
oa22f80 g556039 ( .a(n_10190), .b(n_13414), .c(n_12166), .d(n_12165), .o(n_13362) );
oa22f80 g556040 ( .a(n_11122), .b(n_13909), .c(n_12618), .d(n_12619), .o(n_15211) );
oa12f80 g556041 ( .a(n_13287), .b(n_13286), .c(n_13285), .o(n_15264) );
in01f80 g556042 ( .a(n_15461), .o(n_14603) );
ao12f80 g556043 ( .a(n_13118), .b(n_14146), .c(n_13117), .o(n_15461) );
in01f80 g556044 ( .a(n_14602), .o(n_15435) );
ao12f80 g556045 ( .a(n_13327), .b(n_13326), .c(n_13325), .o(n_14602) );
in01f80 g556046 ( .a(n_14144), .o(n_14145) );
ao12f80 g556047 ( .a(n_12717), .b(n_13384), .c(n_12716), .o(n_14144) );
in01f80 g556048 ( .a(n_13782), .o(n_13783) );
oa22f80 g556049 ( .a(n_11113), .b(n_13939), .c(n_12632), .d(n_12631), .o(n_13782) );
in01f80 g556050 ( .a(n_15434), .o(n_15015) );
ao12f80 g556051 ( .a(n_13689), .b(n_13688), .c(n_13687), .o(n_15434) );
in01f80 g556052 ( .a(n_15878), .o(n_15378) );
ao12f80 g556053 ( .a(n_13292), .b(n_13291), .c(n_13290), .o(n_15878) );
in01f80 g556054 ( .a(n_13780), .o(n_13781) );
oa12f80 g556055 ( .a(n_12162), .b(n_12161), .c(n_12160), .o(n_13780) );
in01f80 g556056 ( .a(n_14142), .o(n_14143) );
ao12f80 g556057 ( .a(n_12711), .b(n_13383), .c(n_12710), .o(n_14142) );
in01f80 g556058 ( .a(n_13778), .o(n_13779) );
ao12f80 g556059 ( .a(n_12212), .b(n_12159), .c(FE_OFN779_n_12158), .o(n_13778) );
in01f80 g556060 ( .a(n_13360), .o(n_13361) );
oa22f80 g556061 ( .a(n_10185), .b(n_13459), .c(n_12156), .d(n_12157), .o(n_13360) );
in01f80 g556062 ( .a(n_14140), .o(n_14141) );
ao12f80 g556063 ( .a(n_12806), .b(n_12805), .c(FE_OFN987_n_12804), .o(n_14140) );
in01f80 g556064 ( .a(n_13776), .o(n_13777) );
ao12f80 g556065 ( .a(n_12211), .b(n_12155), .c(n_12154), .o(n_13776) );
in01f80 g556066 ( .a(n_14600), .o(n_14601) );
oa12f80 g556067 ( .a(n_12982), .b(n_12977), .c(n_12978), .o(n_14600) );
ao12f80 g556068 ( .a(n_12151), .b(n_12210), .c(n_12209), .o(n_15490) );
in01f80 g556069 ( .a(n_16899), .o(n_16011) );
oa12f80 g556070 ( .a(n_13693), .b(n_13692), .c(n_13691), .o(n_16899) );
in01f80 g556071 ( .a(n_15171), .o(n_16053) );
oa12f80 g556072 ( .a(n_13298), .b(n_13297), .c(n_13296), .o(n_15171) );
in01f80 g556073 ( .a(n_14138), .o(n_14139) );
ao12f80 g556074 ( .a(n_12709), .b(n_13382), .c(n_12708), .o(n_14138) );
ao12f80 g556075 ( .a(n_14092), .b(n_14091), .c(n_14090), .o(n_15014) );
in01f80 g556076 ( .a(n_14136), .o(n_14137) );
ao12f80 g556077 ( .a(n_12615), .b(n_12638), .c(n_12637), .o(n_14136) );
in01f80 g556078 ( .a(n_14134), .o(n_14135) );
oa12f80 g556079 ( .a(n_12581), .b(n_12984), .c(n_12983), .o(n_14134) );
in01f80 g556080 ( .a(n_14598), .o(n_14599) );
ao12f80 g556081 ( .a(n_12970), .b(n_12969), .c(n_12968), .o(n_14598) );
ao12f80 g556082 ( .a(n_12838), .b(n_12840), .c(n_12854), .o(n_13775) );
in01f80 g556083 ( .a(n_14132), .o(n_14133) );
oa12f80 g556084 ( .a(n_12577), .b(n_12576), .c(n_12575), .o(n_14132) );
in01f80 g556085 ( .a(n_13773), .o(n_13774) );
oa12f80 g556086 ( .a(n_12182), .b(n_12164), .c(n_12163), .o(n_13773) );
in01f80 g556087 ( .a(n_13771), .o(n_13772) );
oa22f80 g556088 ( .a(n_11167), .b(FE_OFN957_n_13438), .c(n_12148), .d(n_8485), .o(n_13771) );
in01f80 g556089 ( .a(n_15012), .o(n_15013) );
oa12f80 g556090 ( .a(n_13605), .b(n_13521), .c(FE_OFN482_n_13520), .o(n_15012) );
ao12f80 g556091 ( .a(n_13248), .b(n_13247), .c(n_13246), .o(n_14131) );
in01f80 g556092 ( .a(n_15735), .o(n_15359) );
ao12f80 g556093 ( .a(n_13256), .b(n_13255), .c(n_13254), .o(n_15735) );
oa12f80 g556094 ( .a(n_12707), .b(n_13385), .c(n_12706), .o(n_14903) );
oa22f80 g556095 ( .a(n_11661), .b(n_28597), .c(n_83), .d(FE_OFN91_n_27449), .o(n_13359) );
oa22f80 g556096 ( .a(n_11660), .b(FE_OFN234_n_4162), .c(n_1359), .d(FE_OFN1109_rst), .o(n_13358) );
oa22f80 g556097 ( .a(n_11659), .b(FE_OFN296_n_3069), .c(n_1592), .d(FE_OFN62_n_27012), .o(n_13357) );
oa22f80 g556098 ( .a(n_11730), .b(FE_OFN257_n_4280), .c(n_274), .d(FE_OFN1115_rst), .o(n_13770) );
oa22f80 g556099 ( .a(n_11658), .b(n_29033), .c(n_1771), .d(FE_OFN1121_rst), .o(n_13356) );
ao22s80 g556100 ( .a(n_14146), .b(n_13769), .c(n_12719), .d(x_in_56_1), .o(n_14969) );
oa22f80 g556101 ( .a(n_9362), .b(FE_OFN224_n_21642), .c(n_1202), .d(FE_OFN92_n_27449), .o(n_12241) );
oa22f80 g556102 ( .a(n_11049), .b(FE_OFN247_n_4162), .c(n_1502), .d(FE_OFN134_n_27449), .o(n_13355) );
oa22f80 g556103 ( .a(n_12903), .b(FE_OFN406_n_28303), .c(n_948), .d(FE_OFN1120_rst), .o(n_14130) );
oa22f80 g556104 ( .a(n_12854), .b(n_4162), .c(n_975), .d(FE_OFN129_n_27449), .o(n_12855) );
oa22f80 g556105 ( .a(n_10132), .b(FE_OFN260_n_4280), .c(n_1960), .d(FE_OFN127_n_27449), .o(n_12240) );
oa22f80 g556106 ( .a(FE_OFN811_n_12878), .b(n_21076), .c(n_414), .d(FE_OFN324_n_4860), .o(n_14129) );
oa22f80 g556107 ( .a(n_12364), .b(FE_OFN170_n_22948), .c(n_601), .d(n_29617), .o(n_13768) );
oa22f80 g556108 ( .a(n_12872), .b(FE_OFN256_n_4280), .c(n_1491), .d(FE_OFN69_n_27012), .o(n_14128) );
oa22f80 g556109 ( .a(FE_OFN532_n_12317), .b(n_21076), .c(n_157), .d(FE_OFN336_n_4860), .o(n_13767) );
oa22f80 g556110 ( .a(n_12077), .b(n_13241), .c(n_13242), .d(x_in_5_13), .o(n_14996) );
ao22s80 g556111 ( .a(n_12076), .b(x_in_43_13), .c(n_12826), .d(n_7274), .o(n_13766) );
ao22s80 g556112 ( .a(n_12090), .b(x_in_7_11), .c(n_12831), .d(n_7336), .o(n_13765) );
ao22s80 g556113 ( .a(n_12079), .b(x_in_27_12), .c(n_12828), .d(n_7402), .o(n_13764) );
ao22s80 g556114 ( .a(n_12527), .b(x_in_23_11), .c(n_13711), .d(n_7296), .o(n_14127) );
ao22s80 g556115 ( .a(n_12529), .b(x_in_15_11), .c(n_13710), .d(n_7334), .o(n_14126) );
ao22s80 g556116 ( .a(n_12525), .b(x_in_47_11), .c(n_13708), .d(n_7245), .o(n_14125) );
ao22s80 g556117 ( .a(n_12524), .b(x_in_31_11), .c(n_13707), .d(n_7298), .o(n_14124) );
ao22s80 g556118 ( .a(n_12528), .b(x_in_63_11), .c(n_13712), .d(n_7308), .o(n_14123) );
ao22s80 g556119 ( .a(n_12526), .b(x_in_55_11), .c(n_13709), .d(n_7332), .o(n_14122) );
ao22s80 g556120 ( .a(n_14596), .b(x_in_39_11), .c(n_14595), .d(n_7317), .o(n_14597) );
in01f80 g556121 ( .a(n_13354), .o(n_13763) );
ao22s80 g556122 ( .a(n_13353), .b(n_13352), .c(n_13351), .d(n_13350), .o(n_13354) );
na02f80 g556142 ( .a(n_13348), .b(n_13347), .o(n_13349) );
na02f80 g556143 ( .a(n_12852), .b(n_12851), .o(n_12853) );
na02f80 g556144 ( .a(FE_OFN600_n_16000), .b(FE_OFN29_n_13676), .o(n_13853) );
na02f80 g556145 ( .a(n_12850), .b(n_12849), .o(n_14561) );
na02f80 g556146 ( .a(n_12848), .b(n_12847), .o(n_14552) );
na02f80 g556147 ( .a(n_13760), .b(x_in_8_2), .o(n_15039) );
in01f80 g556148 ( .a(n_14120), .o(n_14121) );
no02f80 g556149 ( .a(n_13760), .b(x_in_8_2), .o(n_14120) );
na03f80 g556150 ( .a(n_11624), .b(n_17657), .c(FE_OFN384_n_16289), .o(n_13985) );
in01f80 g556151 ( .a(n_18116), .o(n_14813) );
na02f80 g556152 ( .a(n_15689), .b(x_in_2_0), .o(n_18116) );
na02f80 g556153 ( .a(n_13759), .b(x_in_38_2), .o(n_15040) );
in01f80 g556154 ( .a(n_14118), .o(n_14119) );
no02f80 g556155 ( .a(n_13759), .b(x_in_38_2), .o(n_14118) );
na03f80 g556156 ( .a(n_11656), .b(n_17663), .c(FE_OFN385_n_16289), .o(n_13990) );
na02f80 g556157 ( .a(n_13757), .b(n_13756), .o(n_13758) );
no02f80 g556158 ( .a(n_13345), .b(n_13344), .o(n_13346) );
in01f80 g556159 ( .a(n_13754), .o(n_13755) );
na02f80 g556160 ( .a(n_13343), .b(n_12116), .o(n_13754) );
in01f80 g556161 ( .a(n_18113), .o(n_15682) );
na02f80 g556162 ( .a(n_15698), .b(x_in_34_0), .o(n_18113) );
in01f80 g556163 ( .a(n_13341), .o(n_13342) );
na02f80 g556164 ( .a(n_11085), .b(n_12846), .o(n_13341) );
no02f80 g556165 ( .a(n_13339), .b(n_13338), .o(n_13340) );
no02f80 g556166 ( .a(n_13336), .b(n_13335), .o(n_13337) );
na03f80 g556167 ( .a(n_11655), .b(n_17654), .c(FE_OFN419_n_16909), .o(n_14663) );
na02f80 g556168 ( .a(n_12416), .b(n_884), .o(n_13753) );
in01f80 g556169 ( .a(n_13751), .o(n_13752) );
na02f80 g556170 ( .a(n_11774), .b(n_13334), .o(n_13751) );
no02f80 g556171 ( .a(n_13332), .b(n_13331), .o(n_13333) );
in01f80 g556172 ( .a(n_13329), .o(n_13330) );
na02f80 g556173 ( .a(n_11089), .b(n_12845), .o(n_13329) );
in01f80 g556174 ( .a(n_17645), .o(n_14811) );
na02f80 g556175 ( .a(n_15121), .b(x_in_16_0), .o(n_17645) );
na02f80 g556176 ( .a(n_12385), .b(n_844), .o(n_13750) );
na02f80 g556177 ( .a(n_14116), .b(n_14115), .o(n_14117) );
no02f80 g556178 ( .a(n_13748), .b(n_13747), .o(n_13749) );
na03f80 g556179 ( .a(n_17642), .b(n_11652), .c(FE_OFN382_n_16289), .o(n_14224) );
in01f80 g556180 ( .a(n_17882), .o(n_14469) );
na02f80 g556181 ( .a(n_15694), .b(x_in_18_0), .o(n_17882) );
na02f80 g556182 ( .a(n_11703), .b(n_503), .o(n_13328) );
no02f80 g556183 ( .a(n_13326), .b(n_13325), .o(n_13327) );
na03f80 g556184 ( .a(n_11649), .b(n_17651), .c(FE_OFN422_n_16909), .o(n_14720) );
na02f80 g556185 ( .a(n_13746), .b(n_12539), .o(n_14803) );
no02f80 g556186 ( .a(n_13323), .b(n_13322), .o(n_13324) );
na03f80 g556187 ( .a(n_11646), .b(n_17648), .c(n_16289), .o(n_14694) );
in01f80 g556188 ( .a(n_13320), .o(n_13321) );
na02f80 g556189 ( .a(n_11081), .b(n_12844), .o(n_13320) );
no02f80 g556190 ( .a(n_13318), .b(n_13317), .o(n_13319) );
no02f80 g556191 ( .a(n_13315), .b(n_13314), .o(n_13316) );
na02f80 g556192 ( .a(n_14113), .b(n_14112), .o(n_14114) );
na02f80 g556193 ( .a(n_13313), .b(x_in_0_7), .o(n_14837) );
in01f80 g556194 ( .a(n_13744), .o(n_13745) );
no02f80 g556195 ( .a(n_13313), .b(x_in_0_7), .o(n_13744) );
in01f80 g556196 ( .a(n_13742), .o(n_13743) );
na02f80 g556197 ( .a(n_13312), .b(n_12124), .o(n_13742) );
in01f80 g556198 ( .a(n_17874), .o(n_15030) );
na02f80 g556199 ( .a(n_15696), .b(x_in_50_0), .o(n_17874) );
na02f80 g556200 ( .a(n_13499), .b(n_1616), .o(n_14111) );
na02f80 g556201 ( .a(n_13730), .b(n_13729), .o(n_13741) );
no02f80 g556202 ( .a(n_13739), .b(n_13738), .o(n_13740) );
na02f80 g556203 ( .a(n_12843), .b(n_12842), .o(n_14494) );
in01f80 g556204 ( .a(n_13310), .o(n_13311) );
no02f80 g556205 ( .a(n_12843), .b(n_12842), .o(n_13310) );
na03f80 g556206 ( .a(n_11642), .b(n_17639), .c(FE_OFN383_n_16289), .o(n_14638) );
no02f80 g556207 ( .a(n_13309), .b(n_13308), .o(n_14836) );
in01f80 g556208 ( .a(n_13736), .o(n_13737) );
na02f80 g556209 ( .a(n_13309), .b(n_13308), .o(n_13736) );
in01f80 g556210 ( .a(n_13734), .o(n_13735) );
na02f80 g556211 ( .a(n_13307), .b(n_13306), .o(n_13734) );
no02f80 g556212 ( .a(n_13307), .b(n_13306), .o(n_14835) );
no02f80 g556213 ( .a(n_13732), .b(n_13731), .o(n_13733) );
in01f80 g556214 ( .a(n_13304), .o(n_13305) );
na02f80 g556215 ( .a(n_11087), .b(n_12841), .o(n_13304) );
na03f80 g556216 ( .a(n_12289), .b(n_15868), .c(FE_OFN383_n_16289), .o(n_14285) );
no02f80 g556217 ( .a(n_13302), .b(n_13301), .o(n_13303) );
in01f80 g556218 ( .a(n_14812), .o(n_17666) );
no02f80 g556219 ( .a(n_13730), .b(n_13729), .o(n_14812) );
in01f80 g556220 ( .a(n_17674), .o(n_15029) );
na02f80 g556221 ( .a(n_15428), .b(x_in_10_0), .o(n_17674) );
na02f80 g556222 ( .a(n_13496), .b(n_373), .o(n_14110) );
na03f80 g556223 ( .a(n_11612), .b(n_16510), .c(FE_OFN382_n_16289), .o(n_13924) );
no02f80 g556224 ( .a(n_12840), .b(n_11027), .o(n_14080) );
in01f80 g556225 ( .a(n_17671), .o(n_15031) );
na02f80 g556226 ( .a(n_15377), .b(x_in_42_0), .o(n_17671) );
na02f80 g556227 ( .a(n_12928), .b(n_1903), .o(n_14109) );
na02f80 g556228 ( .a(n_12839), .b(x_in_4_7), .o(n_14499) );
in01f80 g556229 ( .a(n_13299), .o(n_13300) );
no02f80 g556230 ( .a(n_12839), .b(x_in_4_7), .o(n_13299) );
in01f80 g556231 ( .a(n_17877), .o(n_15028) );
na02f80 g556232 ( .a(n_15421), .b(x_in_26_0), .o(n_17877) );
na02f80 g556233 ( .a(n_13493), .b(n_497), .o(n_14108) );
na03f80 g556234 ( .a(n_11643), .b(n_17660), .c(FE_OFN421_n_16909), .o(n_13876) );
na02f80 g556235 ( .a(n_14590), .b(n_1266), .o(n_15010) );
no02f80 g556236 ( .a(n_12840), .b(n_12854), .o(n_12838) );
in01f80 g556237 ( .a(n_14106), .o(n_14107) );
na02f80 g556238 ( .a(n_13728), .b(n_12552), .o(n_14106) );
no02f80 g556239 ( .a(n_11377), .b(n_10325), .o(n_10326) );
na02f80 g556240 ( .a(n_13297), .b(n_13296), .o(n_13298) );
na02f80 g556241 ( .a(n_13726), .b(n_13725), .o(n_13727) );
no02f80 g556242 ( .a(n_12110), .b(x_in_1_9), .o(n_14067) );
na02f80 g556243 ( .a(n_13723), .b(n_13722), .o(n_13724) );
no02f80 g556244 ( .a(n_13294), .b(n_13293), .o(n_13295) );
no02f80 g556245 ( .a(n_13291), .b(n_13290), .o(n_13292) );
no02f80 g556246 ( .a(n_14104), .b(n_14103), .o(n_14105) );
na02f80 g556247 ( .a(n_13720), .b(n_13719), .o(n_13721) );
no02f80 g556248 ( .a(n_12536), .b(n_13718), .o(n_14808) );
no02f80 g556249 ( .a(n_13289), .b(n_13288), .o(n_14832) );
in01f80 g556250 ( .a(n_13716), .o(n_13717) );
na02f80 g556251 ( .a(n_13289), .b(n_13288), .o(n_13716) );
na02f80 g556252 ( .a(n_13286), .b(n_13285), .o(n_13287) );
no02f80 g556253 ( .a(n_13283), .b(n_13282), .o(n_13284) );
no02f80 g556254 ( .a(n_13714), .b(n_13713), .o(n_13715) );
na02f80 g556255 ( .a(n_13280), .b(n_13279), .o(n_13281) );
no02f80 g556256 ( .a(n_13278), .b(n_13277), .o(n_14899) );
na02f80 g556257 ( .a(n_12837), .b(n_12836), .o(n_14490) );
in01f80 g556258 ( .a(n_13275), .o(n_13276) );
no02f80 g556259 ( .a(n_12837), .b(n_12836), .o(n_13275) );
no02f80 g556260 ( .a(n_12835), .b(n_12834), .o(n_14547) );
in01f80 g556261 ( .a(n_13273), .o(n_13274) );
no02f80 g556262 ( .a(n_12833), .b(n_12832), .o(n_13273) );
na02f80 g556263 ( .a(n_12833), .b(n_12832), .o(n_14486) );
oa12f80 g556264 ( .a(n_11671), .b(n_11556), .c(FE_OFN239_n_4162), .o(n_13272) );
oa12f80 g556265 ( .a(FE_OFN9_n_11667), .b(n_11555), .c(n_29683), .o(n_13271) );
oa12f80 g556266 ( .a(n_11665), .b(n_11552), .c(FE_OFN264_n_4280), .o(n_13270) );
oa12f80 g556267 ( .a(n_11663), .b(n_11551), .c(FE_OFN303_n_3069), .o(n_13269) );
oa12f80 g556268 ( .a(n_11669), .b(n_11554), .c(n_28303), .o(n_13268) );
oa12f80 g556269 ( .a(FE_OFN84_n_11673), .b(n_11553), .c(n_23813), .o(n_13267) );
no02f80 g556270 ( .a(n_13712), .b(x_in_63_11), .o(n_14826) );
no02f80 g556271 ( .a(n_13711), .b(x_in_23_11), .o(n_14830) );
no02f80 g556272 ( .a(n_13710), .b(x_in_15_11), .o(n_14828) );
no02f80 g556273 ( .a(n_13709), .b(x_in_55_11), .o(n_14824) );
no02f80 g556274 ( .a(n_12239), .b(n_12238), .o(n_14070) );
no02f80 g556275 ( .a(n_13708), .b(x_in_47_11), .o(n_14822) );
no02f80 g556276 ( .a(n_13707), .b(x_in_31_11), .o(n_14820) );
no02f80 g556277 ( .a(n_12831), .b(x_in_7_11), .o(n_14046) );
na02f80 g556278 ( .a(n_13265), .b(x_in_1_9), .o(n_13266) );
na02f80 g556279 ( .a(n_13498), .b(n_14102), .o(n_15997) );
na02f80 g556280 ( .a(n_13760), .b(n_14102), .o(n_13706) );
na02f80 g556281 ( .a(n_13263), .b(n_13262), .o(n_13264) );
no02f80 g556282 ( .a(n_13704), .b(n_13703), .o(n_13705) );
in01f80 g556283 ( .a(n_13701), .o(n_13702) );
no02f80 g556284 ( .a(n_13261), .b(n_13260), .o(n_13701) );
na02f80 g556285 ( .a(n_13261), .b(n_13260), .o(n_14814) );
oa12f80 g556286 ( .a(n_12868), .b(n_11585), .c(FE_OFN219_n_23315), .o(n_13700) );
in01f80 g556287 ( .a(n_13259), .o(n_14477) );
na02f80 g556288 ( .a(n_12830), .b(n_12829), .o(n_13259) );
no02f80 g556289 ( .a(n_12830), .b(n_12829), .o(n_16297) );
no02f80 g556290 ( .a(n_12828), .b(x_in_27_12), .o(n_14044) );
na02f80 g556291 ( .a(n_13698), .b(n_13697), .o(n_13699) );
no02f80 g556292 ( .a(n_12081), .b(n_13258), .o(n_14503) );
na02f80 g556293 ( .a(n_13695), .b(n_13694), .o(n_13696) );
no02f80 g556294 ( .a(n_13257), .b(n_12508), .o(n_14898) );
na02f80 g556295 ( .a(n_13692), .b(n_13691), .o(n_13693) );
in01f80 g556296 ( .a(n_14100), .o(n_14101) );
no02f80 g556297 ( .a(n_12885), .b(n_5236), .o(n_14100) );
no02f80 g556298 ( .a(n_12884), .b(n_5235), .o(n_14810) );
no02f80 g556299 ( .a(n_13255), .b(n_13254), .o(n_13256) );
no02f80 g556300 ( .a(n_13252), .b(n_13251), .o(n_13253) );
no02f80 g556301 ( .a(n_13249), .b(n_15228), .o(n_13250) );
no02f80 g556302 ( .a(n_13247), .b(n_13246), .o(n_13248) );
no02f80 g556303 ( .a(n_11341), .b(n_12827), .o(n_23674) );
no02f80 g556304 ( .a(n_12826), .b(x_in_43_13), .o(n_14032) );
na02f80 g556305 ( .a(n_13244), .b(n_13243), .o(n_13245) );
in01f80 g556306 ( .a(n_13690), .o(n_15329) );
na02f80 g556307 ( .a(n_13242), .b(n_13241), .o(n_13690) );
ao12f80 g556308 ( .a(n_9799), .b(n_12237), .c(n_9360), .o(n_14488) );
na02f80 g556309 ( .a(n_13239), .b(n_14147), .o(n_13240) );
no02f80 g556310 ( .a(n_13237), .b(n_14147), .o(n_13238) );
no02f80 g556311 ( .a(n_12075), .b(n_13236), .o(n_14514) );
no02f80 g556312 ( .a(n_12823), .b(n_12825), .o(n_25910) );
no02f80 g556313 ( .a(n_12823), .b(n_12822), .o(n_12824) );
na02f80 g556314 ( .a(n_12072), .b(n_13235), .o(n_15577) );
no02f80 g556315 ( .a(n_13688), .b(n_13687), .o(n_13689) );
na02f80 g556316 ( .a(n_14098), .b(n_14097), .o(n_14099) );
na02f80 g556317 ( .a(n_13686), .b(n_13685), .o(n_15027) );
in01f80 g556318 ( .a(n_14095), .o(n_14096) );
no02f80 g556319 ( .a(n_13686), .b(n_13685), .o(n_14095) );
no02f80 g556320 ( .a(n_13233), .b(n_13232), .o(n_13234) );
in01f80 g556321 ( .a(n_13230), .o(n_13231) );
no02f80 g556322 ( .a(n_12821), .b(n_12820), .o(n_13230) );
na02f80 g556323 ( .a(n_12821), .b(n_12820), .o(n_14461) );
in01f80 g556324 ( .a(n_14093), .o(n_14094) );
na02f80 g556325 ( .a(n_12883), .b(n_9111), .o(n_14093) );
na02f80 g556326 ( .a(n_12882), .b(n_9112), .o(n_14806) );
na02f80 g556327 ( .a(n_13683), .b(n_13682), .o(n_13684) );
na02f80 g556328 ( .a(n_12338), .b(n_5187), .o(n_14040) );
na02f80 g556329 ( .a(n_12339), .b(n_5188), .o(n_14460) );
in01f80 g556330 ( .a(n_13680), .o(n_13681) );
no02f80 g556331 ( .a(n_13229), .b(n_13228), .o(n_13680) );
na02f80 g556332 ( .a(n_13229), .b(n_13228), .o(n_14805) );
no02f80 g556333 ( .a(n_14091), .b(n_14090), .o(n_14092) );
no02f80 g556334 ( .a(n_11199), .b(n_12819), .o(n_15233) );
na02f80 g556335 ( .a(n_13798), .b(n_12817), .o(n_12818) );
no02f80 g556336 ( .a(n_13798), .b(n_12815), .o(n_12816) );
na02f80 g556337 ( .a(n_13227), .b(n_13226), .o(n_14801) );
in01f80 g556338 ( .a(n_13678), .o(n_13679) );
no02f80 g556339 ( .a(n_13227), .b(n_13226), .o(n_13678) );
na02f80 g556340 ( .a(n_13677), .b(FE_OFN29_n_13676), .o(n_14624) );
in01f80 g556341 ( .a(n_13224), .o(n_13225) );
na02f80 g556342 ( .a(n_12814), .b(FE_OFN329_n_4860), .o(n_13224) );
na02f80 g556343 ( .a(n_12341), .b(FE_OFN30_n_13676), .o(n_14208) );
na02f80 g556344 ( .a(n_12879), .b(FE_OFN27_n_13676), .o(n_14632) );
na02f80 g556345 ( .a(n_12875), .b(n_13676), .o(n_14628) );
na02f80 g556346 ( .a(n_13675), .b(FE_OFN28_n_13676), .o(n_14630) );
no02f80 g556347 ( .a(n_12483), .b(n_13674), .o(n_27176) );
na02f80 g556348 ( .a(n_12476), .b(n_13673), .o(n_14979) );
oa12f80 g556349 ( .a(n_3855), .b(n_9368), .c(n_32741), .o(n_10324) );
no02f80 g556350 ( .a(n_13211), .b(n_13210), .o(n_14789) );
no02f80 g556351 ( .a(n_12812), .b(n_12811), .o(n_12813) );
in01f80 g556352 ( .a(n_13671), .o(n_13672) );
no02f80 g556353 ( .a(n_13223), .b(n_13222), .o(n_13671) );
na02f80 g556354 ( .a(n_13223), .b(n_13222), .o(n_14791) );
in01f80 g556355 ( .a(n_13220), .o(n_13221) );
na02f80 g556356 ( .a(n_12715), .b(n_12714), .o(n_13220) );
in01f80 g556357 ( .a(n_13218), .o(n_13219) );
no02f80 g556358 ( .a(n_12766), .b(n_12765), .o(n_13218) );
in01f80 g556359 ( .a(n_13216), .o(n_13217) );
na02f80 g556360 ( .a(n_12810), .b(n_12809), .o(n_13216) );
no02f80 g556361 ( .a(n_12810), .b(n_12809), .o(n_14249) );
na02f80 g556362 ( .a(n_13104), .b(n_13103), .o(n_14785) );
in01f80 g556363 ( .a(n_13669), .o(n_13670) );
na02f80 g556364 ( .a(n_13169), .b(n_13168), .o(n_13669) );
in01f80 g556365 ( .a(n_13667), .o(n_13668) );
no02f80 g556366 ( .a(n_13213), .b(n_13212), .o(n_13667) );
in01f80 g556367 ( .a(n_13665), .o(n_13666) );
na02f80 g556368 ( .a(n_13208), .b(n_13207), .o(n_13665) );
in01f80 g556369 ( .a(n_13214), .o(n_13215) );
no02f80 g556370 ( .a(n_11741), .b(n_8258), .o(n_13214) );
na02f80 g556371 ( .a(n_13213), .b(n_13212), .o(n_14787) );
ao12f80 g556372 ( .a(n_11561), .b(n_12506), .c(n_13722), .o(n_15270) );
no02f80 g556373 ( .a(n_11742), .b(n_8259), .o(n_14447) );
in01f80 g556374 ( .a(n_13663), .o(n_13664) );
na02f80 g556375 ( .a(n_13211), .b(n_13210), .o(n_13663) );
na02f80 g556376 ( .a(n_12235), .b(FE_OFN989_n_13374), .o(n_12236) );
na02f80 g556377 ( .a(n_12471), .b(n_13662), .o(n_22872) );
na02f80 g556378 ( .a(n_11805), .b(n_13209), .o(n_15003) );
no02f80 g556379 ( .a(n_12750), .b(n_12749), .o(n_14328) );
oa12f80 g556380 ( .a(n_3863), .b(n_9371), .c(n_32740), .o(n_10323) );
no02f80 g556381 ( .a(n_13661), .b(n_12454), .o(n_19673) );
in01f80 g556382 ( .a(n_17587), .o(n_13660) );
oa12f80 g556383 ( .a(n_12950), .b(n_12306), .c(n_9443), .o(n_17587) );
no02f80 g556384 ( .a(n_12473), .b(n_13659), .o(n_21559) );
in01f80 g556385 ( .a(n_13657), .o(n_13658) );
no02f80 g556386 ( .a(n_12412), .b(n_9706), .o(n_13657) );
no02f80 g556387 ( .a(n_12413), .b(n_9707), .o(n_14795) );
in01f80 g556388 ( .a(n_12808), .o(n_14560) );
oa12f80 g556389 ( .a(n_12137), .b(n_11008), .c(n_13344), .o(n_12808) );
na02f80 g556390 ( .a(n_11043), .b(n_12807), .o(n_14030) );
na02f80 g556391 ( .a(n_12233), .b(n_13376), .o(n_12234) );
no02f80 g556392 ( .a(n_12467), .b(n_13656), .o(n_15973) );
no02f80 g556393 ( .a(n_11726), .b(n_8248), .o(n_14291) );
na02f80 g556394 ( .a(n_12231), .b(n_13375), .o(n_12232) );
no02f80 g556395 ( .a(n_13208), .b(n_13207), .o(n_14788) );
no02f80 g556396 ( .a(n_12805), .b(FE_OFN987_n_12804), .o(n_12806) );
in01f80 g556397 ( .a(n_13654), .o(n_13655) );
na02f80 g556398 ( .a(n_12892), .b(n_7545), .o(n_13654) );
na02f80 g556399 ( .a(n_13206), .b(n_13205), .o(n_14749) );
in01f80 g556400 ( .a(n_13652), .o(n_13653) );
no02f80 g556401 ( .a(n_13206), .b(n_13205), .o(n_13652) );
in01f80 g556402 ( .a(n_12803), .o(n_14553) );
oa12f80 g556403 ( .a(n_12132), .b(n_11002), .c(n_13338), .o(n_12803) );
in01f80 g556404 ( .a(n_13203), .o(n_13204) );
na02f80 g556405 ( .a(n_12799), .b(n_12798), .o(n_13203) );
no02f80 g556406 ( .a(n_12801), .b(FE_OFN572_n_12800), .o(n_12802) );
no02f80 g556407 ( .a(n_12799), .b(n_12798), .o(n_14413) );
na02f80 g556408 ( .a(n_12229), .b(n_13373), .o(n_12230) );
na02f80 g556409 ( .a(n_12797), .b(n_12796), .o(n_14412) );
oa12f80 g556410 ( .a(n_3873), .b(n_9383), .c(n_32738), .o(n_10322) );
in01f80 g556411 ( .a(n_13201), .o(n_13202) );
no02f80 g556412 ( .a(n_12797), .b(n_12796), .o(n_13201) );
in01f80 g556413 ( .a(n_13199), .o(n_13200) );
na02f80 g556414 ( .a(n_12795), .b(n_12794), .o(n_13199) );
no02f80 g556415 ( .a(n_12795), .b(n_12794), .o(n_14405) );
in01f80 g556416 ( .a(n_13650), .o(n_13651) );
na02f80 g556417 ( .a(n_11719), .b(n_8580), .o(n_13650) );
na02f80 g556418 ( .a(n_11718), .b(n_8579), .o(n_14402) );
na02f80 g556419 ( .a(n_11720), .b(n_12793), .o(n_14482) );
in01f80 g556420 ( .a(n_13648), .o(n_13649) );
no02f80 g556421 ( .a(n_11717), .b(n_8571), .o(n_13648) );
no02f80 g556422 ( .a(n_11716), .b(n_8572), .o(n_14399) );
na02f80 g556423 ( .a(n_13386), .b(n_12791), .o(n_12792) );
in01f80 g556424 ( .a(n_13197), .o(n_13198) );
na02f80 g556425 ( .a(n_11714), .b(n_8578), .o(n_13197) );
in01f80 g556426 ( .a(n_12790), .o(n_14558) );
oa12f80 g556427 ( .a(n_12130), .b(n_10998), .c(n_13331), .o(n_12790) );
na02f80 g556428 ( .a(n_11715), .b(n_8577), .o(n_14391) );
in01f80 g556429 ( .a(n_13646), .o(n_13647) );
no02f80 g556430 ( .a(n_11713), .b(n_8574), .o(n_13646) );
no02f80 g556431 ( .a(n_12788), .b(n_12787), .o(n_12789) );
na02f80 g556432 ( .a(n_12227), .b(n_13372), .o(n_12228) );
no02f80 g556433 ( .a(n_11712), .b(n_8575), .o(n_14388) );
na02f80 g556434 ( .a(n_12786), .b(n_12785), .o(n_14387) );
oa12f80 g556435 ( .a(n_3871), .b(n_9380), .c(n_32739), .o(n_10321) );
in01f80 g556436 ( .a(n_13195), .o(n_13196) );
no02f80 g556437 ( .a(n_12786), .b(n_12785), .o(n_13195) );
in01f80 g556438 ( .a(n_13193), .o(n_13194) );
na02f80 g556439 ( .a(n_12784), .b(n_12783), .o(n_13193) );
no02f80 g556440 ( .a(n_12784), .b(n_12783), .o(n_14361) );
in01f80 g556441 ( .a(n_13191), .o(n_13192) );
no02f80 g556442 ( .a(n_12782), .b(n_12781), .o(n_13191) );
na02f80 g556443 ( .a(n_12782), .b(n_12781), .o(n_14363) );
in01f80 g556444 ( .a(n_13189), .o(n_13190) );
na02f80 g556445 ( .a(n_12780), .b(n_12779), .o(n_13189) );
no02f80 g556446 ( .a(n_12780), .b(n_12779), .o(n_14364) );
na02f80 g556447 ( .a(n_13106), .b(n_13105), .o(n_14640) );
in01f80 g556448 ( .a(n_13187), .o(n_13188) );
no02f80 g556449 ( .a(n_12778), .b(n_12777), .o(n_13187) );
in01f80 g556450 ( .a(n_14088), .o(n_14089) );
na02f80 g556451 ( .a(n_12926), .b(n_8818), .o(n_14088) );
na02f80 g556452 ( .a(n_12778), .b(n_12777), .o(n_14365) );
in01f80 g556453 ( .a(n_13185), .o(n_13186) );
na02f80 g556454 ( .a(n_12776), .b(n_12775), .o(n_13185) );
no02f80 g556455 ( .a(n_12776), .b(n_12775), .o(n_14366) );
in01f80 g556456 ( .a(n_13183), .o(n_13184) );
no02f80 g556457 ( .a(n_12774), .b(n_12773), .o(n_13183) );
na02f80 g556458 ( .a(n_12927), .b(n_8819), .o(n_15025) );
na02f80 g556459 ( .a(n_12774), .b(n_12773), .o(n_14367) );
in01f80 g556460 ( .a(n_13181), .o(n_13182) );
na02f80 g556461 ( .a(n_12772), .b(n_12771), .o(n_13181) );
no02f80 g556462 ( .a(n_11938), .b(n_13180), .o(n_26280) );
no02f80 g556463 ( .a(n_12772), .b(n_12771), .o(n_14368) );
in01f80 g556464 ( .a(n_13178), .o(n_13179) );
no02f80 g556465 ( .a(n_12770), .b(n_12769), .o(n_13178) );
na02f80 g556466 ( .a(n_12770), .b(n_12769), .o(n_14369) );
in01f80 g556467 ( .a(n_13176), .o(n_13177) );
na02f80 g556468 ( .a(n_12768), .b(n_12767), .o(n_13176) );
oa12f80 g556469 ( .a(n_11361), .b(n_12851), .c(n_8348), .o(n_14515) );
no02f80 g556470 ( .a(n_12768), .b(n_12767), .o(n_14370) );
in01f80 g556471 ( .a(n_13644), .o(n_13645) );
no02f80 g556472 ( .a(n_13175), .b(n_13174), .o(n_13644) );
na02f80 g556473 ( .a(n_13175), .b(n_13174), .o(n_14728) );
in01f80 g556474 ( .a(n_13642), .o(n_13643) );
no02f80 g556475 ( .a(n_12423), .b(n_11704), .o(n_13642) );
no02f80 g556476 ( .a(n_12424), .b(n_11705), .o(n_14729) );
ao12f80 g556477 ( .a(n_12561), .b(n_13747), .c(n_12098), .o(n_14512) );
no02f80 g556478 ( .a(n_12462), .b(n_13641), .o(n_22877) );
in01f80 g556479 ( .a(n_13172), .o(n_13173) );
na02f80 g556480 ( .a(n_11701), .b(n_8814), .o(n_13172) );
na02f80 g556481 ( .a(n_12766), .b(n_12765), .o(n_14448) );
na02f80 g556482 ( .a(n_11702), .b(n_8815), .o(n_14356) );
na02f80 g556483 ( .a(n_12452), .b(n_13640), .o(n_16871) );
in01f80 g556484 ( .a(n_12764), .o(n_14557) );
oa12f80 g556485 ( .a(n_12126), .b(n_10994), .c(n_13322), .o(n_12764) );
no02f80 g556486 ( .a(n_13170), .b(n_14879), .o(n_13171) );
no02f80 g556487 ( .a(n_12762), .b(FE_OFN1216_n_12761), .o(n_12763) );
na02f80 g556488 ( .a(n_12225), .b(FE_OFN1218_n_13369), .o(n_12226) );
no02f80 g556489 ( .a(n_13170), .b(n_14538), .o(n_14497) );
oa12f80 g556490 ( .a(n_3973), .b(n_9377), .c(n_32737), .o(n_10320) );
no02f80 g556491 ( .a(n_13169), .b(n_13168), .o(n_14786) );
no02f80 g556492 ( .a(n_13380), .b(n_12759), .o(n_12760) );
in01f80 g556493 ( .a(n_12758), .o(n_14537) );
oa12f80 g556494 ( .a(n_12103), .b(n_10959), .c(n_13314), .o(n_12758) );
in01f80 g556495 ( .a(n_12757), .o(n_14556) );
oa12f80 g556496 ( .a(n_12140), .b(n_10990), .c(n_13317), .o(n_12757) );
no02f80 g556497 ( .a(n_12755), .b(FE_OFN1276_n_12754), .o(n_12756) );
na02f80 g556498 ( .a(n_12223), .b(n_13368), .o(n_12224) );
oa12f80 g556499 ( .a(n_3505), .b(n_9374), .c(n_32743), .o(n_10319) );
na02f80 g556500 ( .a(n_13133), .b(n_13132), .o(n_14650) );
oa12f80 g556501 ( .a(n_12945), .b(n_12277), .c(n_14112), .o(n_14900) );
in01f80 g556502 ( .a(n_13638), .o(n_13639) );
no02f80 g556503 ( .a(n_12904), .b(n_12906), .o(n_13638) );
no02f80 g556504 ( .a(n_12905), .b(n_12907), .o(n_14675) );
no02f80 g556505 ( .a(n_12752), .b(n_12751), .o(n_12753) );
in01f80 g556506 ( .a(n_13166), .o(n_13167) );
no02f80 g556507 ( .a(n_12362), .b(n_11471), .o(n_13166) );
no02f80 g556508 ( .a(n_12363), .b(n_12361), .o(n_14329) );
in01f80 g556509 ( .a(n_13636), .o(n_13637) );
na02f80 g556510 ( .a(n_12899), .b(n_11694), .o(n_13636) );
na02f80 g556511 ( .a(n_12900), .b(n_10741), .o(n_14670) );
in01f80 g556512 ( .a(n_13164), .o(n_13165) );
na02f80 g556513 ( .a(n_12750), .b(n_12749), .o(n_13164) );
in01f80 g556514 ( .a(n_13162), .o(n_13163) );
na02f80 g556515 ( .a(n_12359), .b(n_10635), .o(n_13162) );
na02f80 g556516 ( .a(n_12360), .b(n_11693), .o(n_14327) );
in01f80 g556517 ( .a(n_13160), .o(n_13161) );
no02f80 g556518 ( .a(n_12357), .b(n_11692), .o(n_13160) );
no02f80 g556519 ( .a(n_12358), .b(n_10723), .o(n_14326) );
ao12f80 g556520 ( .a(n_11581), .b(n_12530), .c(n_13719), .o(n_14554) );
na02f80 g556521 ( .a(n_13379), .b(n_12747), .o(n_12748) );
in01f80 g556522 ( .a(n_13634), .o(n_13635) );
na02f80 g556523 ( .a(n_12897), .b(n_10724), .o(n_13634) );
na02f80 g556524 ( .a(n_12898), .b(n_11695), .o(n_14669) );
in01f80 g556525 ( .a(n_13632), .o(n_13633) );
na02f80 g556526 ( .a(n_11757), .b(n_12354), .o(n_13632) );
na02f80 g556527 ( .a(n_11756), .b(n_12355), .o(n_14325) );
no02f80 g556528 ( .a(n_11727), .b(n_8249), .o(n_24513) );
na02f80 g556529 ( .a(n_13631), .b(n_13630), .o(n_15023) );
in01f80 g556530 ( .a(n_14086), .o(n_14087) );
no02f80 g556531 ( .a(n_13631), .b(n_13630), .o(n_14086) );
in01f80 g556532 ( .a(n_13158), .o(n_13159) );
na02f80 g556533 ( .a(n_12746), .b(n_12745), .o(n_13158) );
no02f80 g556534 ( .a(n_12746), .b(n_12745), .o(n_14314) );
in01f80 g556535 ( .a(n_13156), .o(n_13157) );
no02f80 g556536 ( .a(n_12744), .b(n_12743), .o(n_13156) );
no02f80 g556537 ( .a(n_12814), .b(n_12045), .o(n_14966) );
na02f80 g556538 ( .a(n_12744), .b(n_12743), .o(n_14315) );
in01f80 g556539 ( .a(n_13154), .o(n_13155) );
na02f80 g556540 ( .a(n_12742), .b(n_12741), .o(n_13154) );
no02f80 g556541 ( .a(n_12742), .b(n_12741), .o(n_14316) );
in01f80 g556542 ( .a(n_13152), .o(n_13153) );
no02f80 g556543 ( .a(n_12740), .b(n_12739), .o(n_13152) );
na02f80 g556544 ( .a(n_12740), .b(n_12739), .o(n_14317) );
in01f80 g556545 ( .a(n_13150), .o(n_13151) );
na02f80 g556546 ( .a(n_12738), .b(n_12737), .o(n_13150) );
no02f80 g556547 ( .a(n_12738), .b(n_12737), .o(n_14318) );
in01f80 g556548 ( .a(n_13148), .o(n_13149) );
no02f80 g556549 ( .a(n_12736), .b(n_12735), .o(n_13148) );
na02f80 g556550 ( .a(n_12736), .b(n_12735), .o(n_14319) );
no02f80 g556551 ( .a(n_12734), .b(n_12733), .o(n_14320) );
in01f80 g556552 ( .a(n_13146), .o(n_13147) );
na02f80 g556553 ( .a(n_12734), .b(n_12733), .o(n_13146) );
in01f80 g556554 ( .a(n_13628), .o(n_13629) );
no02f80 g556555 ( .a(n_13145), .b(n_13144), .o(n_13628) );
na02f80 g556556 ( .a(n_13145), .b(n_13144), .o(n_14662) );
no02f80 g556557 ( .a(n_13627), .b(n_12435), .o(n_17793) );
no02f80 g556558 ( .a(n_11143), .b(n_12732), .o(n_23696) );
oa12f80 g556559 ( .a(n_11768), .b(n_10934), .c(n_13262), .o(n_13143) );
no02f80 g556560 ( .a(n_13141), .b(n_13140), .o(n_13142) );
na02f80 g556561 ( .a(n_12893), .b(n_7546), .o(n_14653) );
in01f80 g556562 ( .a(n_13138), .o(n_13139) );
na02f80 g556563 ( .a(n_12345), .b(n_11688), .o(n_13138) );
na02f80 g556564 ( .a(n_12346), .b(n_11689), .o(n_14295) );
in01f80 g556565 ( .a(n_12731), .o(n_14559) );
oa12f80 g556566 ( .a(n_12129), .b(n_11000), .c(n_13335), .o(n_12731) );
no02f80 g556567 ( .a(n_13136), .b(FE_OFN817_n_13135), .o(n_13137) );
oa12f80 g556568 ( .a(n_12106), .b(n_10964), .c(n_9199), .o(n_14072) );
na02f80 g556569 ( .a(n_11828), .b(n_13134), .o(n_24352) );
no02f80 g556570 ( .a(n_12270), .b(n_13135), .o(n_14565) );
in01f80 g556571 ( .a(n_13625), .o(n_13626) );
no02f80 g556572 ( .a(n_13133), .b(n_13132), .o(n_13625) );
in01f80 g556573 ( .a(n_13130), .o(n_13131) );
na02f80 g556574 ( .a(n_12730), .b(n_12729), .o(n_13130) );
no02f80 g556575 ( .a(n_12730), .b(n_12729), .o(n_14277) );
na02f80 g556576 ( .a(n_12727), .b(n_12726), .o(n_12728) );
na02f80 g556577 ( .a(n_12725), .b(n_12724), .o(n_14276) );
in01f80 g556578 ( .a(n_13128), .o(n_13129) );
no02f80 g556579 ( .a(n_12725), .b(n_12724), .o(n_13128) );
in01f80 g556580 ( .a(n_13126), .o(n_13127) );
na02f80 g556581 ( .a(n_12723), .b(n_12722), .o(n_13126) );
no02f80 g556582 ( .a(n_12723), .b(n_12722), .o(n_14272) );
in01f80 g556583 ( .a(n_13623), .o(n_13624) );
na02f80 g556584 ( .a(n_12337), .b(n_8568), .o(n_13623) );
na02f80 g556585 ( .a(n_12336), .b(n_8567), .o(n_14271) );
ao12f80 g556586 ( .a(n_13301), .b(n_10315), .c(n_10314), .o(n_13488) );
in01f80 g556587 ( .a(n_13124), .o(n_13125) );
na02f80 g556588 ( .a(n_12721), .b(n_12720), .o(n_13124) );
no02f80 g556589 ( .a(n_12721), .b(n_12720), .o(n_14267) );
in01f80 g556590 ( .a(n_13621), .o(n_13622) );
na02f80 g556591 ( .a(n_12328), .b(n_8560), .o(n_13621) );
na02f80 g556592 ( .a(n_12327), .b(n_8559), .o(n_14266) );
in01f80 g556593 ( .a(n_13619), .o(n_13620) );
no02f80 g556594 ( .a(n_12335), .b(n_8554), .o(n_13619) );
no02f80 g556595 ( .a(n_12334), .b(n_8555), .o(n_14265) );
in01f80 g556596 ( .a(n_13122), .o(n_13123) );
na02f80 g556597 ( .a(n_12332), .b(n_8551), .o(n_13122) );
no02f80 g556598 ( .a(n_11817), .b(n_13121), .o(n_25544) );
in01f80 g556599 ( .a(n_13617), .o(n_13618) );
na02f80 g556600 ( .a(n_12880), .b(n_8948), .o(n_13617) );
na02f80 g556601 ( .a(n_12881), .b(n_8949), .o(n_14649) );
no02f80 g556602 ( .a(n_13120), .b(n_11813), .o(n_19667) );
in01f80 g556603 ( .a(n_15102), .o(n_13119) );
no02f80 g556604 ( .a(n_12719), .b(n_13117), .o(n_15102) );
no02f80 g556605 ( .a(n_14146), .b(n_13117), .o(n_13118) );
no02f80 g556606 ( .a(n_13115), .b(n_14876), .o(n_13116) );
na02f80 g556607 ( .a(n_12333), .b(n_8550), .o(n_14281) );
in01f80 g556608 ( .a(n_12718), .o(n_14528) );
ao12f80 g556609 ( .a(n_12066), .b(n_10853), .c(n_13325), .o(n_12718) );
no02f80 g556610 ( .a(n_13115), .b(n_14529), .o(n_14475) );
oa12f80 g556611 ( .a(n_12290), .b(n_12960), .c(n_14097), .o(n_16004) );
no02f80 g556612 ( .a(n_13384), .b(n_12716), .o(n_12717) );
na02f80 g556613 ( .a(n_11796), .b(n_13114), .o(n_24550) );
na02f80 g556614 ( .a(n_11989), .b(n_13113), .o(n_18661) );
no02f80 g556615 ( .a(n_13112), .b(n_12040), .o(n_17790) );
na02f80 g556616 ( .a(n_11811), .b(n_13111), .o(n_16863) );
no02f80 g556617 ( .a(n_11808), .b(n_13110), .o(n_15969) );
no02f80 g556618 ( .a(n_11785), .b(n_13109), .o(n_24198) );
in01f80 g556619 ( .a(n_13615), .o(n_13616) );
na02f80 g556620 ( .a(n_12876), .b(n_8252), .o(n_13615) );
na02f80 g556621 ( .a(n_12877), .b(n_8253), .o(n_14646) );
no02f80 g556622 ( .a(n_12715), .b(n_12714), .o(n_14292) );
no02f80 g556623 ( .a(n_12935), .b(n_14085), .o(n_21557) );
na02f80 g556624 ( .a(n_12468), .b(n_13614), .o(n_18670) );
na02f80 g556625 ( .a(n_13381), .b(n_12712), .o(n_12713) );
no02f80 g556626 ( .a(n_12221), .b(n_14855), .o(n_12222) );
in01f80 g556627 ( .a(n_13612), .o(n_13613) );
na02f80 g556628 ( .a(n_12873), .b(n_6603), .o(n_13612) );
na02f80 g556629 ( .a(n_12874), .b(n_6602), .o(n_14645) );
no02f80 g556630 ( .a(n_12221), .b(n_14526), .o(n_14473) );
no02f80 g556631 ( .a(n_13383), .b(n_12710), .o(n_12711) );
in01f80 g556632 ( .a(n_14083), .o(n_14084) );
na02f80 g556633 ( .a(n_13494), .b(n_8959), .o(n_14083) );
oa12f80 g556634 ( .a(n_11613), .b(n_12540), .c(n_13697), .o(n_16017) );
na02f80 g556635 ( .a(n_13495), .b(n_8960), .o(n_15024) );
ao12f80 g556636 ( .a(n_11621), .b(n_11606), .c(n_12555), .o(n_14063) );
na02f80 g556637 ( .a(n_11778), .b(n_13108), .o(n_24532) );
ao12f80 g556638 ( .a(n_10877), .b(n_12073), .c(n_13279), .o(n_15295) );
no02f80 g556639 ( .a(n_12350), .b(n_13107), .o(n_14463) );
no02f80 g556640 ( .a(n_13382), .b(n_12708), .o(n_12709) );
in01f80 g556641 ( .a(n_13610), .o(n_13611) );
no02f80 g556642 ( .a(n_13106), .b(n_13105), .o(n_13610) );
oa12f80 g556643 ( .a(n_10586), .b(n_12078), .c(n_13347), .o(n_14075) );
in01f80 g556644 ( .a(n_13608), .o(n_13609) );
no02f80 g556645 ( .a(n_13104), .b(n_13103), .o(n_13608) );
oa12f80 g556646 ( .a(n_12139), .b(n_11004), .c(n_13254), .o(n_14531) );
in01f80 g556647 ( .a(n_13606), .o(n_13607) );
no02f80 g556648 ( .a(n_12870), .b(n_8250), .o(n_13606) );
no02f80 g556649 ( .a(n_13101), .b(n_14881), .o(n_13102) );
no02f80 g556650 ( .a(n_13101), .b(n_14071), .o(n_14517) );
no02f80 g556651 ( .a(n_12871), .b(n_8251), .o(n_14798) );
na02f80 g556652 ( .a(n_13385), .b(n_12706), .o(n_12707) );
oa12f80 g556653 ( .a(n_13099), .b(n_994), .c(FE_OFN113_n_27449), .o(n_13100) );
oa12f80 g556654 ( .a(n_13099), .b(n_1594), .c(FE_OFN329_n_4860), .o(n_13098) );
oa12f80 g556655 ( .a(n_12503), .b(n_11545), .c(n_13703), .o(n_14551) );
ao12f80 g556656 ( .a(n_11541), .b(n_12502), .c(n_13691), .o(n_15445) );
na02f80 g556657 ( .a(n_10254), .b(n_13484), .o(n_12220) );
ao12f80 g556658 ( .a(n_12498), .b(n_11534), .c(n_13756), .o(n_14550) );
na02f80 g556659 ( .a(n_12931), .b(n_8390), .o(n_16232) );
ao12f80 g556660 ( .a(n_12450), .b(n_11462), .c(n_13713), .o(n_14042) );
oa12f80 g556661 ( .a(n_10954), .b(n_12101), .c(n_10601), .o(n_14549) );
oa12f80 g556662 ( .a(n_10952), .b(n_12100), .c(n_10600), .o(n_14548) );
na02f80 g556663 ( .a(n_10253), .b(n_13475), .o(n_12219) );
ao12f80 g556664 ( .a(n_12507), .b(n_13738), .c(n_11563), .o(n_14545) );
oa12f80 g556665 ( .a(n_10940), .b(n_12095), .c(n_10604), .o(n_14546) );
na02f80 g556666 ( .a(n_13469), .b(n_10211), .o(n_12218) );
ao12f80 g556667 ( .a(n_12501), .b(n_13682), .c(n_11539), .o(n_14897) );
oa12f80 g556668 ( .a(n_12866), .b(n_12946), .c(n_14103), .o(n_14621) );
ao12f80 g556669 ( .a(n_10710), .b(n_11847), .c(n_14147), .o(n_14069) );
oa22f80 g556670 ( .a(n_12426), .b(n_8963), .c(n_11396), .d(n_12425), .o(n_14462) );
in01f80 g556671 ( .a(n_12704), .o(n_12705) );
na03f80 g556672 ( .a(n_7047), .b(n_12217), .c(n_4948), .o(n_12704) );
ao12f80 g556673 ( .a(n_11326), .b(n_12217), .c(n_9295), .o(n_14021) );
ao22s80 g556674 ( .a(n_11376), .b(n_7846), .c(n_8510), .d(n_8509), .o(n_15944) );
na02f80 g556675 ( .a(n_11261), .b(n_13949), .o(n_12703) );
ao22s80 g556676 ( .a(n_11375), .b(n_7809), .c(n_8452), .d(n_8451), .o(n_15948) );
no02f80 g556677 ( .a(n_11213), .b(n_13906), .o(n_12702) );
na02f80 g556678 ( .a(n_11212), .b(n_13977), .o(n_12701) );
no02f80 g556679 ( .a(n_11205), .b(n_13869), .o(n_12700) );
no02f80 g556680 ( .a(n_11204), .b(n_13889), .o(n_12699) );
ao12f80 g556681 ( .a(n_12136), .b(n_13725), .c(n_12556), .o(n_13097) );
na02f80 g556682 ( .a(n_11200), .b(n_14000), .o(n_12698) );
na02f80 g556683 ( .a(n_10227), .b(n_13432), .o(n_12216) );
no02f80 g556684 ( .a(n_10221), .b(n_13447), .o(n_12215) );
no02f80 g556685 ( .a(n_10217), .b(n_13435), .o(n_12214) );
na02f80 g556686 ( .a(n_10213), .b(n_13417), .o(n_12213) );
in01f80 g556687 ( .a(n_13095), .o(n_13096) );
ao22s80 g556688 ( .a(n_10780), .b(n_9603), .c(n_12627), .d(n_12697), .o(n_13095) );
no02f80 g556689 ( .a(n_10186), .b(n_13462), .o(n_12212) );
no02f80 g556690 ( .a(n_10201), .b(n_13456), .o(n_12211) );
oa22f80 g556691 ( .a(n_10772), .b(n_12601), .c(n_14014), .d(n_12602), .o(n_15209) );
ao22s80 g556692 ( .a(n_12058), .b(n_12696), .c(n_12695), .d(n_12057), .o(n_13994) );
ao22s80 g556693 ( .a(n_13094), .b(n_12692), .c(n_12693), .d(n_13093), .o(n_14397) );
oa22f80 g556694 ( .a(n_12210), .b(n_12149), .c(n_12150), .d(n_12209), .o(n_13401) );
oa12f80 g556695 ( .a(n_14396), .b(n_12693), .c(n_12692), .o(n_12694) );
oa22f80 g556696 ( .a(n_12691), .b(n_12684), .c(n_12685), .d(n_12690), .o(n_14009) );
na02f80 g556697 ( .a(n_12727), .b(n_9087), .o(n_12689) );
oa22f80 g556698 ( .a(n_11196), .b(n_12688), .c(n_12687), .d(n_11195), .o(n_14012) );
ao12f80 g556699 ( .a(n_11337), .b(n_11336), .c(n_11335), .o(n_13919) );
no02f80 g556700 ( .a(n_10182), .b(n_13393), .o(n_12208) );
ao12f80 g556701 ( .a(n_14008), .b(n_12685), .c(n_12684), .o(n_12686) );
na02f80 g556702 ( .a(n_11820), .b(n_14455), .o(n_13092) );
no02f80 g556703 ( .a(n_10210), .b(n_13424), .o(n_12207) );
ao22s80 g556704 ( .a(n_13091), .b(n_6581), .c(n_11404), .d(FE_OFN1190_n_13090), .o(n_14456) );
oa22f80 g556705 ( .a(n_11171), .b(n_12683), .c(n_12682), .d(FE_OFN478_n_11170), .o(n_14004) );
na02f80 g556706 ( .a(n_10197), .b(n_13444), .o(n_12206) );
ao12f80 g556707 ( .a(n_10223), .b(n_12205), .c(n_10222), .o(n_13448) );
oa22f80 g556708 ( .a(n_10208), .b(n_12204), .c(n_12203), .d(n_10207), .o(n_13410) );
in01f80 g556709 ( .a(n_13088), .o(n_13089) );
ao12f80 g556710 ( .a(n_11307), .b(n_11306), .c(n_11305), .o(n_13088) );
oa12f80 g556711 ( .a(n_10206), .b(n_11375), .c(n_10205), .o(n_13413) );
ao22s80 g556712 ( .a(n_12202), .b(n_5843), .c(n_9696), .d(FE_OFN1186_n_12201), .o(n_13445) );
na02f80 g556713 ( .a(n_12440), .b(n_14792), .o(n_13605) );
ao12f80 g556714 ( .a(n_12039), .b(n_12639), .c(FE_OFN484_n_12038), .o(n_14453) );
in01f80 g556715 ( .a(n_13086), .o(n_13087) );
oa12f80 g556716 ( .a(n_11293), .b(n_11292), .c(n_11291), .o(n_13086) );
oa22f80 g556717 ( .a(n_13085), .b(n_13081), .c(n_13082), .d(n_13084), .o(n_14450) );
ao12f80 g556718 ( .a(n_14449), .b(n_13082), .c(n_13081), .o(n_13083) );
no02f80 g556719 ( .a(n_12752), .b(n_8653), .o(n_12681) );
ao12f80 g556720 ( .a(n_11350), .b(n_11349), .c(x_in_43_12), .o(n_12680) );
oa12f80 g556721 ( .a(n_10193), .b(n_12200), .c(n_11148), .o(n_13422) );
oa12f80 g556722 ( .a(n_11374), .b(n_11373), .c(x_in_1_8), .o(n_14061) );
in01f80 g556723 ( .a(n_12678), .o(n_12679) );
oa12f80 g556724 ( .a(n_10272), .b(n_10271), .c(n_10270), .o(n_12678) );
oa12f80 g556725 ( .a(n_10238), .b(n_10237), .c(n_10236), .o(n_13428) );
oa12f80 g556726 ( .a(n_10219), .b(n_12199), .c(n_10218), .o(n_13436) );
in01f80 g556727 ( .a(n_13079), .o(n_13080) );
ao12f80 g556728 ( .a(n_11244), .b(n_11243), .c(n_11682), .o(n_13079) );
ao12f80 g556729 ( .a(n_11360), .b(n_11359), .c(x_in_7_10), .o(n_12677) );
ao12f80 g556730 ( .a(n_10225), .b(n_12198), .c(n_10224), .o(n_13433) );
in01f80 g556731 ( .a(n_12675), .o(n_12676) );
oa12f80 g556732 ( .a(n_10266), .b(n_10265), .c(n_10264), .o(n_12675) );
ao22s80 g556733 ( .a(n_11202), .b(n_12197), .c(n_12196), .d(n_11201), .o(n_13451) );
ao12f80 g556734 ( .a(n_12563), .b(n_12867), .c(n_5904), .o(n_13604) );
in01f80 g556735 ( .a(n_13602), .o(n_13603) );
oa12f80 g556736 ( .a(n_12035), .b(n_12034), .c(n_12033), .o(n_13602) );
oa12f80 g556737 ( .a(n_11165), .b(n_11164), .c(n_11163), .o(n_13944) );
oa12f80 g556738 ( .a(n_12027), .b(n_12026), .c(n_12025), .o(n_14214) );
oa22f80 g556739 ( .a(n_9574), .b(n_23315), .c(n_740), .d(FE_OFN133_n_27449), .o(n_12195) );
in01f80 g556740 ( .a(n_13600), .o(n_13601) );
ao12f80 g556741 ( .a(n_12024), .b(n_12023), .c(n_12022), .o(n_13600) );
oa12f80 g556742 ( .a(n_11865), .b(n_11864), .c(n_11863), .o(n_14212) );
in01f80 g556743 ( .a(n_13598), .o(n_13599) );
oa12f80 g556744 ( .a(n_11975), .b(n_11974), .c(n_11973), .o(n_13598) );
in01f80 g556745 ( .a(n_13596), .o(n_13597) );
ao12f80 g556746 ( .a(n_12021), .b(n_12020), .c(n_12019), .o(n_13596) );
ao12f80 g556747 ( .a(n_10215), .b(n_12194), .c(n_10214), .o(n_13418) );
oa22f80 g556748 ( .a(n_9571), .b(FE_OFN292_n_3069), .c(n_1773), .d(FE_OFN101_n_27449), .o(n_12193) );
oa12f80 g556749 ( .a(n_11162), .b(n_12674), .c(n_12673), .o(n_14065) );
ao12f80 g556750 ( .a(n_11352), .b(n_11351), .c(x_in_27_11), .o(n_12672) );
in01f80 g556751 ( .a(n_13594), .o(n_13595) );
ao12f80 g556752 ( .a(n_11987), .b(n_11986), .c(n_11985), .o(n_13594) );
oa22f80 g556753 ( .a(n_9573), .b(FE_OFN406_n_28303), .c(n_1666), .d(FE_OFN355_n_4860), .o(n_12192) );
oa12f80 g556754 ( .a(n_10204), .b(n_12191), .c(n_11168), .o(n_13442) );
na02f80 g556755 ( .a(n_10203), .b(n_13429), .o(n_12190) );
oa22f80 g556756 ( .a(n_9570), .b(FE_OFN198_n_29637), .c(n_846), .d(FE_OFN94_n_27449), .o(n_12189) );
in01f80 g556757 ( .a(n_13592), .o(n_13593) );
ao12f80 g556758 ( .a(n_12037), .b(n_12036), .c(n_12351), .o(n_13592) );
in01f80 g556759 ( .a(n_13590), .o(n_13591) );
ao12f80 g556760 ( .a(n_12029), .b(n_12028), .c(n_12368), .o(n_13590) );
in01f80 g556761 ( .a(n_13588), .o(n_13589) );
ao12f80 g556762 ( .a(n_11999), .b(n_11998), .c(n_11997), .o(n_13588) );
in01f80 g556763 ( .a(n_13586), .o(n_13587) );
oa12f80 g556764 ( .a(n_11996), .b(n_11995), .c(n_11994), .o(n_13586) );
oa22f80 g556765 ( .a(n_9569), .b(FE_OFN411_n_28303), .c(n_1681), .d(FE_OFN364_n_4860), .o(n_12188) );
oa12f80 g556766 ( .a(n_11099), .b(n_11098), .c(n_11097), .o(n_13863) );
ao12f80 g556767 ( .a(n_12003), .b(n_12002), .c(n_12001), .o(n_14431) );
oa12f80 g556768 ( .a(n_11984), .b(n_11983), .c(n_11982), .o(n_14423) );
in01f80 g556769 ( .a(n_13584), .o(n_13585) );
ao12f80 g556770 ( .a(n_11981), .b(n_11980), .c(n_11979), .o(n_13584) );
oa12f80 g556771 ( .a(n_11978), .b(n_11977), .c(n_11976), .o(n_14358) );
ao12f80 g556772 ( .a(n_11816), .b(n_11815), .c(n_11814), .o(n_14294) );
in01f80 g556773 ( .a(n_13582), .o(n_13583) );
oa12f80 g556774 ( .a(n_12014), .b(n_12013), .c(n_12012), .o(n_13582) );
in01f80 g556775 ( .a(n_13580), .o(n_13581) );
ao12f80 g556776 ( .a(n_11972), .b(n_11971), .c(n_12318), .o(n_13580) );
oa12f80 g556777 ( .a(n_11194), .b(n_11193), .c(n_11192), .o(n_13983) );
oa12f80 g556778 ( .a(n_11970), .b(n_11969), .c(n_11968), .o(n_14236) );
oa12f80 g556779 ( .a(n_12018), .b(n_12017), .c(FE_OFN1196_n_12016), .o(n_14324) );
in01f80 g556780 ( .a(n_13077), .o(n_13078) );
oa12f80 g556781 ( .a(n_11191), .b(n_11190), .c(n_11189), .o(n_13077) );
in01f80 g556782 ( .a(n_13075), .o(n_13076) );
ao12f80 g556783 ( .a(n_11272), .b(n_11271), .c(n_11270), .o(n_13075) );
in01f80 g556784 ( .a(n_13073), .o(n_13074) );
ao12f80 g556785 ( .a(n_11222), .b(n_11221), .c(n_11220), .o(n_13073) );
in01f80 g556786 ( .a(n_13071), .o(n_13072) );
oa12f80 g556787 ( .a(n_11184), .b(n_11183), .c(n_11182), .o(n_13071) );
in01f80 g556788 ( .a(n_13069), .o(n_13070) );
ao12f80 g556789 ( .a(n_11247), .b(n_11246), .c(n_11245), .o(n_13069) );
ao22s80 g556790 ( .a(n_12187), .b(n_3053), .c(n_9681), .d(FE_OFN1254_n_12186), .o(n_13430) );
in01f80 g556791 ( .a(n_13067), .o(n_13068) );
oa12f80 g556792 ( .a(n_11290), .b(n_11289), .c(n_11288), .o(n_13067) );
in01f80 g556793 ( .a(n_13065), .o(n_13066) );
ao12f80 g556794 ( .a(n_11159), .b(n_11158), .c(n_11157), .o(n_13065) );
oa12f80 g556795 ( .a(n_11966), .b(n_11965), .c(n_11964), .o(n_14401) );
in01f80 g556796 ( .a(n_13578), .o(n_13579) );
ao12f80 g556797 ( .a(n_11963), .b(n_11962), .c(n_11961), .o(n_13578) );
oa12f80 g556798 ( .a(n_11960), .b(n_11959), .c(n_11958), .o(n_14393) );
in01f80 g556799 ( .a(n_13063), .o(n_13064) );
ao12f80 g556800 ( .a(n_11208), .b(n_11207), .c(n_11206), .o(n_13063) );
in01f80 g556801 ( .a(n_13576), .o(n_13577) );
ao12f80 g556802 ( .a(n_11957), .b(n_11956), .c(n_11955), .o(n_13576) );
in01f80 g556803 ( .a(n_13574), .o(n_13575) );
oa12f80 g556804 ( .a(n_11954), .b(n_11953), .c(n_11952), .o(n_13574) );
in01f80 g556805 ( .a(n_13572), .o(n_13573) );
ao12f80 g556806 ( .a(n_11951), .b(n_11950), .c(n_11949), .o(n_13572) );
in01f80 g556807 ( .a(n_13570), .o(n_13571) );
ao12f80 g556808 ( .a(n_11948), .b(n_11947), .c(n_11946), .o(n_13570) );
oa12f80 g556809 ( .a(n_11945), .b(n_11944), .c(n_11943), .o(n_14390) );
ao22s80 g556810 ( .a(n_12671), .b(n_2580), .c(n_10485), .d(n_12670), .o(n_13978) );
in01f80 g556811 ( .a(n_13061), .o(n_13062) );
oa12f80 g556812 ( .a(n_11228), .b(n_11227), .c(n_11226), .o(n_13061) );
ao12f80 g556813 ( .a(n_11329), .b(n_11328), .c(n_11327), .o(n_13976) );
in01f80 g556814 ( .a(n_13059), .o(n_13060) );
oa12f80 g556815 ( .a(n_11240), .b(n_11239), .c(n_11238), .o(n_13059) );
in01f80 g556816 ( .a(n_13057), .o(n_13058) );
ao12f80 g556817 ( .a(n_11234), .b(n_11233), .c(n_11232), .o(n_13057) );
in01f80 g556818 ( .a(n_13055), .o(n_13056) );
oa12f80 g556819 ( .a(n_11254), .b(n_11253), .c(n_11252), .o(n_13055) );
in01f80 g556820 ( .a(n_13053), .o(n_13054) );
ao12f80 g556821 ( .a(n_11216), .b(n_11215), .c(n_11214), .o(n_13053) );
in01f80 g556822 ( .a(n_13051), .o(n_13052) );
oa12f80 g556823 ( .a(n_11332), .b(n_11331), .c(n_11330), .o(n_13051) );
in01f80 g556824 ( .a(n_13049), .o(n_13050) );
oa12f80 g556825 ( .a(n_11225), .b(n_11224), .c(n_11223), .o(n_13049) );
in01f80 g556826 ( .a(n_13047), .o(n_13048) );
oa12f80 g556827 ( .a(n_11156), .b(n_11155), .c(n_11154), .o(n_13047) );
in01f80 g556828 ( .a(n_13568), .o(n_13569) );
oa12f80 g556829 ( .a(n_12055), .b(n_12054), .c(n_12053), .o(n_13568) );
oa12f80 g556830 ( .a(n_12006), .b(n_12005), .c(n_12004), .o(n_14435) );
oa22f80 g556831 ( .a(n_12185), .b(n_6519), .c(n_9698), .d(FE_OFN480_n_12184), .o(n_13425) );
oa12f80 g556832 ( .a(n_11862), .b(n_11861), .c(n_11860), .o(n_14467) );
in01f80 g556833 ( .a(n_13045), .o(n_13046) );
ao12f80 g556834 ( .a(n_11260), .b(n_11259), .c(n_11258), .o(n_13045) );
ao12f80 g556835 ( .a(n_10327), .b(n_12183), .c(n_10779), .o(n_13470) );
ao12f80 g556836 ( .a(n_11936), .b(n_11935), .c(n_12367), .o(n_14355) );
in01f80 g556837 ( .a(n_13043), .o(n_13044) );
oa12f80 g556838 ( .a(n_11237), .b(n_11236), .c(n_11235), .o(n_13043) );
oa12f80 g556839 ( .a(n_11934), .b(n_11933), .c(n_12373), .o(n_14349) );
in01f80 g556840 ( .a(n_13041), .o(n_13042) );
ao12f80 g556841 ( .a(n_11287), .b(n_11286), .c(n_11285), .o(n_13041) );
in01f80 g556842 ( .a(n_13566), .o(n_13567) );
ao12f80 g556843 ( .a(n_11929), .b(n_11928), .c(n_11927), .o(n_13566) );
in01f80 g556844 ( .a(n_13564), .o(n_13565) );
oa12f80 g556845 ( .a(n_11932), .b(n_11931), .c(n_11930), .o(n_13564) );
in01f80 g556846 ( .a(n_13039), .o(n_13040) );
oa12f80 g556847 ( .a(n_11257), .b(n_11256), .c(n_11255), .o(n_13039) );
in01f80 g556848 ( .a(n_13562), .o(n_13563) );
ao12f80 g556849 ( .a(n_11926), .b(n_11925), .c(n_11924), .o(n_13562) );
in01f80 g556850 ( .a(n_13560), .o(n_13561) );
ao12f80 g556851 ( .a(n_11923), .b(n_11922), .c(n_11921), .o(n_13560) );
in01f80 g556852 ( .a(n_13037), .o(n_13038) );
ao12f80 g556853 ( .a(n_11319), .b(n_11318), .c(n_11317), .o(n_13037) );
ao12f80 g556854 ( .a(n_11917), .b(n_11916), .c(n_11915), .o(n_14341) );
in01f80 g556855 ( .a(n_13558), .o(n_13559) );
oa12f80 g556856 ( .a(n_11920), .b(n_11919), .c(n_11918), .o(n_13558) );
in01f80 g556857 ( .a(n_13035), .o(n_13036) );
oa12f80 g556858 ( .a(n_11345), .b(n_11344), .c(n_11343), .o(n_13035) );
in01f80 g556859 ( .a(n_13556), .o(n_13557) );
ao12f80 g556860 ( .a(n_11914), .b(n_11913), .c(n_11912), .o(n_13556) );
in01f80 g556861 ( .a(n_13554), .o(n_13555) );
oa12f80 g556862 ( .a(n_11911), .b(n_11910), .c(n_11909), .o(n_13554) );
oa12f80 g556863 ( .a(n_11908), .b(n_11907), .c(n_11906), .o(n_14339) );
in01f80 g556864 ( .a(n_12668), .o(n_12669) );
ao12f80 g556865 ( .a(n_10298), .b(n_10297), .c(n_10296), .o(n_12668) );
in01f80 g556866 ( .a(n_13552), .o(n_13553) );
oa12f80 g556867 ( .a(n_11905), .b(n_11904), .c(n_11903), .o(n_13552) );
oa12f80 g556868 ( .a(n_11152), .b(n_11151), .c(n_11150), .o(n_14880) );
in01f80 g556869 ( .a(n_12666), .o(n_12667) );
ao12f80 g556870 ( .a(n_10246), .b(n_10245), .c(n_10244), .o(n_12666) );
in01f80 g556871 ( .a(n_13550), .o(n_13551) );
ao12f80 g556872 ( .a(n_11902), .b(n_11901), .c(n_11900), .o(n_13550) );
oa22f80 g556873 ( .a(n_10384), .b(n_12665), .c(n_12664), .d(n_9774), .o(n_24557) );
in01f80 g556874 ( .a(n_13548), .o(n_13549) );
oa12f80 g556875 ( .a(n_11898), .b(n_11897), .c(FE_OFN1192_n_11896), .o(n_13548) );
in01f80 g556876 ( .a(n_12662), .o(n_12663) );
oa12f80 g556877 ( .a(n_10290), .b(n_10289), .c(n_10288), .o(n_12662) );
in01f80 g556878 ( .a(n_13546), .o(n_13547) );
ao12f80 g556879 ( .a(n_11895), .b(n_11894), .c(n_11893), .o(n_13546) );
ao12f80 g556880 ( .a(n_12093), .b(n_12092), .c(n_12091), .o(n_14510) );
oa12f80 g556881 ( .a(n_11892), .b(n_11891), .c(FE_OFN1101_n_12369), .o(n_14337) );
in01f80 g556882 ( .a(n_13544), .o(n_13545) );
ao12f80 g556883 ( .a(n_11890), .b(n_11889), .c(n_12372), .o(n_13544) );
oa12f80 g556884 ( .a(n_11888), .b(n_11887), .c(n_12371), .o(n_14335) );
in01f80 g556885 ( .a(n_13542), .o(n_13543) );
ao12f80 g556886 ( .a(n_11886), .b(n_11885), .c(n_12370), .o(n_13542) );
in01f80 g556887 ( .a(n_13540), .o(n_13541) );
oa12f80 g556888 ( .a(n_11884), .b(n_11883), .c(n_11882), .o(n_13540) );
in01f80 g556889 ( .a(n_13538), .o(n_13539) );
ao12f80 g556890 ( .a(n_11881), .b(n_11880), .c(n_11879), .o(n_13538) );
in01f80 g556891 ( .a(n_13536), .o(n_13537) );
oa12f80 g556892 ( .a(n_11878), .b(n_11877), .c(n_11876), .o(n_13536) );
oa12f80 g556893 ( .a(n_11875), .b(n_11874), .c(n_11873), .o(n_14333) );
in01f80 g556894 ( .a(n_13033), .o(n_13034) );
ao12f80 g556895 ( .a(n_11275), .b(n_11274), .c(n_11273), .o(n_13033) );
oa12f80 g556896 ( .a(n_10301), .b(n_10300), .c(n_10299), .o(n_13397) );
in01f80 g556897 ( .a(n_13534), .o(n_13535) );
oa12f80 g556898 ( .a(n_11872), .b(n_11871), .c(n_11870), .o(n_13534) );
in01f80 g556899 ( .a(n_12660), .o(n_12661) );
ao12f80 g556900 ( .a(n_10278), .b(n_10277), .c(n_10276), .o(n_12660) );
in01f80 g556901 ( .a(n_13532), .o(n_13533) );
ao12f80 g556902 ( .a(n_12032), .b(n_12031), .c(n_12030), .o(n_13532) );
in01f80 g556903 ( .a(n_13031), .o(n_13032) );
oa12f80 g556904 ( .a(n_11181), .b(n_11180), .c(n_11179), .o(n_13031) );
in01f80 g556905 ( .a(n_12658), .o(n_12659) );
oa12f80 g556906 ( .a(n_10318), .b(n_10317), .c(n_10316), .o(n_12658) );
in01f80 g556907 ( .a(n_12656), .o(n_12657) );
ao12f80 g556908 ( .a(n_10307), .b(n_10306), .c(n_10305), .o(n_12656) );
na02f80 g556909 ( .a(n_10181), .b(n_13403), .o(n_12182) );
in01f80 g556910 ( .a(n_12654), .o(n_12655) );
oa12f80 g556911 ( .a(n_10313), .b(n_10312), .c(n_10311), .o(n_12654) );
in01f80 g556912 ( .a(n_12652), .o(n_12653) );
ao12f80 g556913 ( .a(n_10233), .b(n_10232), .c(n_10231), .o(n_12652) );
in01f80 g556914 ( .a(n_13530), .o(n_13531) );
oa12f80 g556915 ( .a(n_12113), .b(n_12112), .c(n_12111), .o(n_13530) );
in01f80 g556916 ( .a(n_12650), .o(n_12651) );
ao12f80 g556917 ( .a(n_10230), .b(n_10229), .c(n_10228), .o(n_12650) );
oa22f80 g556918 ( .a(n_13030), .b(n_12979), .c(n_12980), .d(n_13029), .o(n_14238) );
in01f80 g556919 ( .a(n_13027), .o(n_13028) );
oa12f80 g556920 ( .a(n_11369), .b(n_11368), .c(n_11367), .o(n_13027) );
ao12f80 g556921 ( .a(n_10196), .b(n_10195), .c(n_10194), .o(n_14534) );
in01f80 g556922 ( .a(n_12648), .o(n_12649) );
ao12f80 g556923 ( .a(n_10310), .b(n_10309), .c(n_10308), .o(n_12648) );
ao22s80 g556924 ( .a(n_12647), .b(n_2494), .c(n_10416), .d(n_12646), .o(n_13950) );
in01f80 g556925 ( .a(n_12644), .o(n_12645) );
ao12f80 g556926 ( .a(n_10192), .b(n_10191), .c(n_11070), .o(n_12644) );
oa22f80 g556927 ( .a(n_11218), .b(n_12643), .c(n_12642), .d(n_11217), .o(n_13913) );
oa12f80 g556928 ( .a(n_11263), .b(n_11262), .c(x_in_51_12), .o(n_14029) );
in01f80 g556929 ( .a(n_13025), .o(n_13026) );
ao22s80 g556930 ( .a(n_12641), .b(n_9051), .c(FE_OFN1085_n_14427), .d(n_12640), .o(n_13025) );
in01f80 g556931 ( .a(n_32732), .o(n_14048) );
oa12f80 g556933 ( .a(n_11852), .b(n_11851), .c(n_11850), .o(n_14311) );
oa22f80 g556934 ( .a(n_9572), .b(FE_OFN293_n_3069), .c(n_1576), .d(n_29068), .o(n_12181) );
no03m80 g556935 ( .a(n_12449), .b(n_12102), .c(n_9536), .o(n_13529) );
in01f80 g556936 ( .a(n_13527), .o(n_13528) );
oa12f80 g556937 ( .a(n_11868), .b(n_11867), .c(n_11866), .o(n_13527) );
oa22f80 g556938 ( .a(n_12639), .b(n_9467), .c(n_14452), .d(n_5912), .o(n_15803) );
oa22f80 g556939 ( .a(n_12638), .b(n_12613), .c(n_12614), .d(n_12637), .o(n_13865) );
oa22f80 g556940 ( .a(n_12636), .b(x_in_33_12), .c(n_10409), .d(n_12635), .o(n_14038) );
oa22f80 g556941 ( .a(n_12180), .b(n_9017), .c(n_13929), .d(n_12179), .o(n_15513) );
oa12f80 g556942 ( .a(n_11846), .b(n_11845), .c(n_11844), .o(n_14309) );
oa12f80 g556943 ( .a(n_11843), .b(n_11842), .c(n_11841), .o(n_13024) );
ao22s80 g556944 ( .a(n_11241), .b(n_12178), .c(n_12177), .d(x_in_33_11), .o(n_13479) );
ao22s80 g556945 ( .a(n_10403), .b(n_12634), .c(n_12633), .d(x_in_33_10), .o(n_14035) );
in01f80 g556946 ( .a(n_14592), .o(n_14593) );
ao12f80 g556947 ( .a(n_12939), .b(n_12938), .c(n_12937), .o(n_14592) );
in01f80 g556948 ( .a(n_13525), .o(n_13526) );
oa12f80 g556949 ( .a(n_12070), .b(n_12069), .c(FE_OFN1232_n_12068), .o(n_13525) );
ao22s80 g556950 ( .a(n_12176), .b(n_8884), .c(n_9579), .d(x_in_33_9), .o(n_13476) );
oa12f80 g556951 ( .a(n_11840), .b(n_11839), .c(n_11838), .o(n_13023) );
in01f80 g556952 ( .a(n_13021), .o(n_13022) );
ao12f80 g556953 ( .a(n_11142), .b(n_11141), .c(n_11140), .o(n_13021) );
in01f80 g556954 ( .a(n_13019), .o(n_13020) );
oa12f80 g556955 ( .a(n_11304), .b(n_11303), .c(n_11302), .o(n_13019) );
ao22s80 g556956 ( .a(n_11250), .b(n_12175), .c(n_12174), .d(x_in_33_8), .o(n_13473) );
in01f80 g556957 ( .a(n_13017), .o(n_13018) );
ao12f80 g556958 ( .a(n_11139), .b(n_11138), .c(n_11137), .o(n_13017) );
ao22s80 g556959 ( .a(n_12632), .b(n_11111), .c(n_11112), .d(n_12631), .o(n_13940) );
oa12f80 g556960 ( .a(n_11136), .b(n_11135), .c(n_11134), .o(n_13938) );
oa12f80 g556961 ( .a(n_11093), .b(n_11092), .c(n_11091), .o(n_14018) );
ao22s80 g556962 ( .a(n_12173), .b(n_8885), .c(n_9615), .d(x_in_33_7), .o(n_13485) );
ao22s80 g556963 ( .a(n_11248), .b(n_12172), .c(n_12171), .d(x_in_33_6), .o(n_13482) );
oa22f80 g556964 ( .a(n_11298), .b(x_in_33_5), .c(n_12630), .d(n_11297), .o(n_13935) );
oa12f80 g556965 ( .a(n_11231), .b(n_11230), .c(n_11229), .o(n_13933) );
in01f80 g556966 ( .a(n_13015), .o(n_13016) );
ao12f80 g556967 ( .a(n_11133), .b(n_11132), .c(n_11131), .o(n_13015) );
in01f80 g556968 ( .a(n_13013), .o(n_13014) );
ao22s80 g556969 ( .a(n_12629), .b(n_9014), .c(n_14282), .d(n_12628), .o(n_13013) );
in01f80 g556970 ( .a(n_13523), .o(n_13524) );
ao12f80 g556971 ( .a(n_11836), .b(n_11835), .c(n_12344), .o(n_13523) );
oa22f80 g556972 ( .a(n_10402), .b(n_12179), .c(n_12180), .d(n_9016), .o(n_13930) );
oa12f80 g556973 ( .a(n_11834), .b(n_11833), .c(n_11832), .o(n_13012) );
in01f80 g556974 ( .a(n_13010), .o(n_13011) );
oa12f80 g556975 ( .a(n_11130), .b(n_11129), .c(n_12627), .o(n_13010) );
in01f80 g556976 ( .a(n_13008), .o(n_13009) );
oa22f80 g556977 ( .a(n_12626), .b(n_10341), .c(n_14278), .d(n_12625), .o(n_13008) );
oa12f80 g556978 ( .a(n_10690), .b(n_11827), .c(n_10689), .o(n_12170) );
ao22s80 g556979 ( .a(n_11384), .b(n_12628), .c(n_12629), .d(n_9013), .o(n_14283) );
in01f80 g556980 ( .a(n_14896), .o(n_13522) );
ao12f80 g556981 ( .a(n_11824), .b(n_13007), .c(n_11823), .o(n_14896) );
oa12f80 g556982 ( .a(n_10685), .b(n_10701), .c(n_10684), .o(n_12624) );
na02f80 g556983 ( .a(n_11822), .b(n_14268), .o(n_13006) );
oa22f80 g556984 ( .a(n_11391), .b(n_12625), .c(n_12626), .d(FE_OFN1200_n_10340), .o(n_14279) );
oa22f80 g556985 ( .a(n_9599), .b(n_12169), .c(n_12168), .d(n_12167), .o(n_15588) );
no02f80 g556986 ( .a(n_11821), .b(n_14262), .o(n_13005) );
ao22s80 g556987 ( .a(n_13004), .b(n_6553), .c(n_11390), .d(FE_OFN1198_n_13003), .o(n_14269) );
oa22f80 g556988 ( .a(n_13002), .b(n_6542), .c(n_11389), .d(n_13001), .o(n_14263) );
oa12f80 g556989 ( .a(n_11325), .b(n_11324), .c(n_11323), .o(n_13927) );
in01f80 g556990 ( .a(n_12999), .o(n_13000) );
oa12f80 g556991 ( .a(n_11281), .b(n_11280), .c(n_11279), .o(n_12999) );
in01f80 g556992 ( .a(n_12622), .o(n_12623) );
ao12f80 g556993 ( .a(n_10287), .b(n_10286), .c(n_10285), .o(n_12622) );
in01f80 g556994 ( .a(n_12997), .o(n_12998) );
oa12f80 g556995 ( .a(n_11313), .b(n_11312), .c(n_11311), .o(n_12997) );
in01f80 g556996 ( .a(n_12995), .o(n_12996) );
ao12f80 g556997 ( .a(n_11316), .b(n_11315), .c(n_11314), .o(n_12995) );
ao12f80 g556998 ( .a(n_11371), .b(n_10980), .c(n_10094), .o(n_14571) );
ao22s80 g556999 ( .a(n_12166), .b(n_10188), .c(n_10189), .d(n_12165), .o(n_13415) );
in01f80 g557000 ( .a(n_12993), .o(n_12994) );
oa12f80 g557001 ( .a(n_11310), .b(n_11309), .c(n_11308), .o(n_12993) );
in01f80 g557002 ( .a(n_12991), .o(n_12992) );
oa12f80 g557003 ( .a(n_11380), .b(n_11379), .c(n_11378), .o(n_12991) );
oa12f80 g557004 ( .a(n_11117), .b(n_11116), .c(n_11115), .o(n_14877) );
in01f80 g557005 ( .a(n_12620), .o(n_12621) );
oa12f80 g557006 ( .a(n_10295), .b(n_10294), .c(n_10293), .o(n_12620) );
ao12f80 g557007 ( .a(n_12444), .b(n_12443), .c(n_12442), .o(n_14648) );
oa22f80 g557008 ( .a(n_11121), .b(n_12619), .c(n_12618), .d(n_11120), .o(n_13910) );
oa22f80 g557009 ( .a(n_12617), .b(n_2366), .c(n_10373), .d(n_12616), .o(n_13907) );
in01f80 g557010 ( .a(n_12989), .o(n_12990) );
ao12f80 g557011 ( .a(n_11284), .b(n_11283), .c(n_11282), .o(n_12989) );
oa12f80 g557012 ( .a(n_12119), .b(n_12118), .c(n_12117), .o(n_14492) );
ao22s80 g557013 ( .a(n_13521), .b(n_5974), .c(n_12246), .d(FE_OFN482_n_13520), .o(n_14793) );
oa12f80 g557014 ( .a(n_11354), .b(n_11353), .c(x_in_5_12), .o(n_14054) );
ao12f80 g557015 ( .a(n_13864), .b(n_12614), .c(n_12613), .o(n_12615) );
in01f80 g557016 ( .a(n_12611), .o(n_12612) );
oa12f80 g557017 ( .a(n_10249), .b(n_10248), .c(n_10247), .o(n_12611) );
in01f80 g557018 ( .a(n_12609), .o(n_12610) );
ao12f80 g557019 ( .a(n_10263), .b(n_10262), .c(n_10261), .o(n_12609) );
in01f80 g557020 ( .a(n_12607), .o(n_12608) );
oa12f80 g557021 ( .a(n_10241), .b(n_10240), .c(n_10239), .o(n_12607) );
ao22s80 g557022 ( .a(n_12164), .b(n_5833), .c(n_9575), .d(n_12163), .o(n_13404) );
oa22f80 g557023 ( .a(n_11321), .b(n_12606), .c(n_12605), .d(n_11320), .o(n_13896) );
in01f80 g557024 ( .a(n_12987), .o(n_12988) );
oa12f80 g557025 ( .a(n_11296), .b(n_11295), .c(n_11294), .o(n_12987) );
in01f80 g557026 ( .a(n_12985), .o(n_12986) );
ao12f80 g557027 ( .a(n_11269), .b(n_11268), .c(n_11267), .o(n_12985) );
ao22s80 g557028 ( .a(n_12984), .b(n_12579), .c(n_12580), .d(n_12983), .o(n_14274) );
oa12f80 g557029 ( .a(n_11356), .b(n_11355), .c(n_11683), .o(n_14856) );
in01f80 g557030 ( .a(n_12603), .o(n_12604) );
oa12f80 g557031 ( .a(n_10284), .b(n_10283), .c(n_10282), .o(n_12603) );
oa12f80 g557032 ( .a(n_11108), .b(n_11107), .c(n_11106), .o(n_14562) );
na02f80 g557033 ( .a(n_10187), .b(n_13406), .o(n_12162) );
oa22f80 g557034 ( .a(n_10364), .b(n_12602), .c(n_12601), .d(FE_OFN783_n_10771), .o(n_14015) );
ao22s80 g557035 ( .a(n_12161), .b(n_6543), .c(n_9589), .d(n_12160), .o(n_13407) );
oa22f80 g557036 ( .a(n_12159), .b(n_6541), .c(n_9586), .d(FE_OFN779_n_12158), .o(n_13463) );
oa22f80 g557037 ( .a(n_12600), .b(n_2480), .c(n_10361), .d(n_12599), .o(n_13890) );
oa22f80 g557038 ( .a(n_10184), .b(n_12157), .c(n_12156), .d(FE_OFN1226_n_10183), .o(n_13460) );
na02f80 g557039 ( .a(n_11784), .b(n_14240), .o(n_12982) );
oa22f80 g557040 ( .a(n_12155), .b(n_6540), .c(n_9585), .d(n_12154), .o(n_13457) );
ao12f80 g557041 ( .a(n_14237), .b(n_12980), .c(n_12979), .o(n_12981) );
oa22f80 g557042 ( .a(n_11385), .b(n_12978), .c(n_12977), .d(n_6460), .o(n_14241) );
in01f80 g557043 ( .a(n_12975), .o(n_12976) );
oa22f80 g557044 ( .a(n_12598), .b(n_8113), .c(n_9242), .d(n_9241), .o(n_12975) );
in01f80 g557045 ( .a(n_13518), .o(n_13519) );
ao12f80 g557046 ( .a(n_11783), .b(n_12598), .c(n_11782), .o(n_13518) );
ao22s80 g557047 ( .a(n_12153), .b(FE_OFN785_n_10198), .c(n_10199), .d(n_12152), .o(n_13454) );
ao12f80 g557048 ( .a(n_13400), .b(n_12150), .c(n_12149), .o(n_12151) );
ao12f80 g557049 ( .a(n_11105), .b(n_11104), .c(n_11103), .o(n_13887) );
ao22s80 g557050 ( .a(n_12597), .b(n_2379), .c(n_10552), .d(n_12596), .o(n_14001) );
oa12f80 g557051 ( .a(n_10275), .b(n_10274), .c(n_10273), .o(n_13399) );
in01f80 g557052 ( .a(n_12594), .o(n_12595) );
oa12f80 g557053 ( .a(n_10252), .b(n_10251), .c(n_10250), .o(n_12594) );
in01f80 g557054 ( .a(n_12592), .o(n_12593) );
ao12f80 g557055 ( .a(n_10260), .b(n_10259), .c(n_10258), .o(n_12592) );
in01f80 g557056 ( .a(n_12590), .o(n_12591) );
oa12f80 g557057 ( .a(n_10257), .b(n_10256), .c(n_10255), .o(n_12590) );
in01f80 g557058 ( .a(n_12588), .o(n_12589) );
ao12f80 g557059 ( .a(n_10243), .b(n_10242), .c(n_10576), .o(n_12588) );
in01f80 g557060 ( .a(n_12973), .o(n_12974) );
oa12f80 g557061 ( .a(n_11266), .b(n_11265), .c(n_11264), .o(n_12973) );
in01f80 g557062 ( .a(n_12971), .o(n_12972) );
ao12f80 g557063 ( .a(n_11278), .b(n_11277), .c(n_11276), .o(n_12971) );
ao12f80 g557064 ( .a(n_11110), .b(n_11109), .c(FE_OFN1204_n_11679), .o(n_13875) );
ao22s80 g557065 ( .a(n_12587), .b(n_8981), .c(n_14226), .d(n_12586), .o(n_15765) );
in01f80 g557066 ( .a(n_13516), .o(n_13517) );
oa12f80 g557067 ( .a(n_12044), .b(n_12043), .c(n_12042), .o(n_13516) );
in01f80 g557068 ( .a(n_13514), .o(n_13515) );
ao12f80 g557069 ( .a(n_12009), .b(n_12008), .c(n_12007), .o(n_13514) );
in01f80 g557070 ( .a(n_12584), .o(n_12585) );
oa12f80 g557071 ( .a(n_10281), .b(n_10280), .c(n_10279), .o(n_12584) );
oa22f80 g557072 ( .a(n_12641), .b(n_9050), .c(n_11382), .d(n_12640), .o(n_14428) );
ao12f80 g557073 ( .a(n_10202), .b(n_12148), .c(n_11166), .o(n_13439) );
oa12f80 g557074 ( .a(n_11993), .b(n_11992), .c(n_11991), .o(n_14433) );
oa22f80 g557075 ( .a(n_12583), .b(n_2400), .c(n_10353), .d(n_12582), .o(n_13870) );
ao22s80 g557076 ( .a(n_11383), .b(n_12586), .c(n_12587), .d(n_8980), .o(n_14227) );
ao22s80 g557077 ( .a(n_10732), .b(n_8905), .c(n_12365), .d(n_8906), .o(n_13966) );
oa12f80 g557078 ( .a(FE_OFN1081_n_14273), .b(n_12580), .c(n_12579), .o(n_12581) );
no02f80 g557079 ( .a(n_11775), .b(n_14219), .o(n_12970) );
ao12f80 g557080 ( .a(n_11363), .b(n_11366), .c(n_11362), .o(n_12578) );
na02f80 g557081 ( .a(n_11100), .b(n_13859), .o(n_12577) );
oa22f80 g557082 ( .a(n_12969), .b(n_6513), .c(n_11386), .d(n_12968), .o(n_14220) );
in01f80 g557083 ( .a(n_12966), .o(n_12967) );
oa12f80 g557084 ( .a(n_11188), .b(n_11187), .c(n_11186), .o(n_12966) );
ao22s80 g557085 ( .a(n_12576), .b(n_6562), .c(n_10352), .d(n_12575), .o(n_13860) );
in01f80 g557086 ( .a(n_12964), .o(n_12965) );
ao12f80 g557087 ( .a(n_11178), .b(n_11177), .c(n_11176), .o(n_12964) );
in01f80 g557088 ( .a(n_12962), .o(n_12963) );
oa12f80 g557089 ( .a(n_11096), .b(n_11095), .c(n_11094), .o(n_12962) );
in01f80 g557090 ( .a(n_13512), .o(n_13513) );
ao12f80 g557091 ( .a(n_12109), .b(n_12108), .c(n_12107), .o(n_13512) );
ao22s80 g557092 ( .a(n_9578), .b(n_12147), .c(n_12146), .d(n_6582), .o(n_13394) );
in01f80 g557093 ( .a(n_12573), .o(n_12574) );
oa12f80 g557094 ( .a(n_10304), .b(n_10303), .c(n_10302), .o(n_12573) );
oa12f80 g557095 ( .a(n_10269), .b(n_10268), .c(n_10267), .o(n_13392) );
oa12f80 g557096 ( .a(n_10180), .b(n_11376), .c(n_10179), .o(n_13390) );
oa12f80 g557097 ( .a(n_11348), .b(n_11347), .c(n_11346), .o(n_14882) );
ao12f80 g557098 ( .a(n_11211), .b(n_11210), .c(n_11209), .o(n_13946) );
oa22f80 g557099 ( .a(n_9693), .b(n_29046), .c(n_1661), .d(FE_OFN92_n_27449), .o(n_12145) );
oa22f80 g557100 ( .a(FE_OFN680_n_9691), .b(n_29046), .c(n_1135), .d(n_27449), .o(n_12144) );
ao22s80 g557101 ( .a(n_13007), .b(n_12572), .c(n_11147), .d(x_in_24_1), .o(n_14026) );
oa22f80 g557102 ( .a(n_10423), .b(FE_OFN406_n_28303), .c(n_1673), .d(FE_OFN127_n_27449), .o(n_12571) );
oa22f80 g557103 ( .a(n_9688), .b(FE_OFN296_n_3069), .c(n_1006), .d(FE_OFN336_n_4860), .o(n_12143) );
oa22f80 g557104 ( .a(n_10487), .b(n_28682), .c(n_1679), .d(FE_OFN1110_rst), .o(n_12570) );
oa22f80 g557105 ( .a(n_11397), .b(n_22019), .c(n_1481), .d(n_27449), .o(n_12961) );
ao22s80 g557106 ( .a(n_12087), .b(n_11041), .c(n_11670), .d(n_8061), .o(n_12569) );
ao22s80 g557107 ( .a(n_12089), .b(n_11037), .c(n_11666), .d(n_8071), .o(n_12568) );
ao22s80 g557108 ( .a(n_12088), .b(n_11696), .c(n_11668), .d(n_8067), .o(n_12567) );
ao22s80 g557109 ( .a(n_12086), .b(n_11040), .c(n_11672), .d(n_8063), .o(n_12566) );
ao22s80 g557110 ( .a(n_12085), .b(n_11034), .c(n_11664), .d(n_8069), .o(n_12565) );
ao22s80 g557111 ( .a(n_12084), .b(n_11698), .c(n_11662), .d(n_8058), .o(n_12564) );
no02f80 g557138 ( .a(n_12537), .b(x_in_39_10), .o(n_12563) );
no02f80 g557139 ( .a(n_13747), .b(n_12561), .o(n_12562) );
na02f80 g557140 ( .a(n_11373), .b(x_in_1_8), .o(n_11374) );
in01f80 g557141 ( .a(n_12141), .o(n_12142) );
na02f80 g557142 ( .a(n_11372), .b(n_14073), .o(n_12141) );
na02f80 g557143 ( .a(n_10981), .b(n_7852), .o(n_11371) );
no02f80 g557144 ( .a(n_12291), .b(n_12960), .o(n_14098) );
na02f80 g557145 ( .a(n_10991), .b(n_12140), .o(n_13318) );
na02f80 g557146 ( .a(n_11005), .b(n_12139), .o(n_13255) );
na02f80 g557147 ( .a(n_12295), .b(n_12959), .o(n_14487) );
no02f80 g557148 ( .a(n_11011), .b(n_12138), .o(n_13920) );
na02f80 g557149 ( .a(n_11009), .b(n_12137), .o(n_13345) );
na02f80 g557150 ( .a(n_12555), .b(n_12135), .o(n_12136) );
in01f80 g557151 ( .a(n_12559), .o(n_12560) );
na02f80 g557152 ( .a(n_11015), .b(n_12134), .o(n_12559) );
in01f80 g557153 ( .a(n_12557), .o(n_12558) );
na02f80 g557154 ( .a(n_11013), .b(n_12133), .o(n_12557) );
na02f80 g557155 ( .a(n_12556), .b(n_12555), .o(n_13726) );
na02f80 g557156 ( .a(n_11003), .b(n_12132), .o(n_13339) );
na02f80 g557157 ( .a(n_9383), .b(n_32738), .o(n_9384) );
in01f80 g557158 ( .a(n_12553), .o(n_12554) );
na02f80 g557159 ( .a(n_12131), .b(n_10978), .o(n_12553) );
na02f80 g557160 ( .a(n_10999), .b(n_12130), .o(n_13332) );
na02f80 g557161 ( .a(n_9380), .b(n_32739), .o(n_9381) );
na02f80 g557162 ( .a(n_11001), .b(n_12129), .o(n_13336) );
in01f80 g557163 ( .a(n_12551), .o(n_12552) );
no02f80 g557164 ( .a(n_12128), .b(n_12127), .o(n_12551) );
na02f80 g557165 ( .a(n_12128), .b(n_12127), .o(n_13728) );
na02f80 g557166 ( .a(n_10995), .b(n_12126), .o(n_13323) );
na02f80 g557167 ( .a(n_9377), .b(n_32737), .o(n_9378) );
in01f80 g557168 ( .a(n_12549), .o(n_12550) );
na02f80 g557169 ( .a(n_12125), .b(n_10993), .o(n_12549) );
na02f80 g557170 ( .a(n_9374), .b(n_32743), .o(n_9375) );
na02f80 g557171 ( .a(n_11370), .b(x_in_0_6), .o(n_13312) );
in01f80 g557172 ( .a(n_12123), .o(n_12124) );
no02f80 g557173 ( .a(n_11370), .b(x_in_0_6), .o(n_12123) );
in01f80 g557174 ( .a(n_12957), .o(n_12958) );
na02f80 g557175 ( .a(n_12548), .b(n_11618), .o(n_12957) );
in01f80 g557176 ( .a(n_13510), .o(n_13511) );
na02f80 g557177 ( .a(n_12299), .b(n_12956), .o(n_13510) );
na02f80 g557178 ( .a(n_10317), .b(n_10316), .o(n_10318) );
na02f80 g557179 ( .a(n_11368), .b(n_11367), .o(n_11369) );
in01f80 g557180 ( .a(n_13508), .o(n_13509) );
na02f80 g557181 ( .a(n_12297), .b(n_12955), .o(n_13508) );
in01f80 g557182 ( .a(n_13506), .o(n_13507) );
na02f80 g557183 ( .a(n_12305), .b(n_12954), .o(n_13506) );
in01f80 g557184 ( .a(n_13504), .o(n_13505) );
na02f80 g557185 ( .a(n_12303), .b(n_12953), .o(n_13504) );
in01f80 g557186 ( .a(n_13502), .o(n_13503) );
na02f80 g557187 ( .a(n_12301), .b(n_12952), .o(n_13502) );
no02f80 g557188 ( .a(n_11464), .b(n_32733), .o(n_12547) );
na02f80 g557189 ( .a(n_9371), .b(n_32740), .o(n_9372) );
no02f80 g557190 ( .a(n_10315), .b(n_10314), .o(n_13301) );
na02f80 g557191 ( .a(n_9368), .b(n_32741), .o(n_9369) );
in01f80 g557192 ( .a(n_13500), .o(n_13501) );
na02f80 g557193 ( .a(n_12293), .b(n_12951), .o(n_13500) );
in01f80 g557194 ( .a(n_12545), .o(n_12546) );
na02f80 g557195 ( .a(n_11021), .b(n_12122), .o(n_12545) );
in01f80 g557196 ( .a(n_12543), .o(n_12544) );
na02f80 g557197 ( .a(n_11019), .b(n_12121), .o(n_12543) );
in01f80 g557198 ( .a(n_12541), .o(n_12542) );
na02f80 g557199 ( .a(n_11017), .b(n_12120), .o(n_12541) );
na02f80 g557200 ( .a(n_11366), .b(n_11365), .o(n_12840) );
na02f80 g557201 ( .a(n_12118), .b(n_12117), .o(n_12119) );
in01f80 g557202 ( .a(n_12115), .o(n_12116) );
no02f80 g557203 ( .a(n_11364), .b(x_in_4_6), .o(n_12115) );
no02f80 g557204 ( .a(n_11614), .b(n_12540), .o(n_13698) );
na02f80 g557205 ( .a(n_12307), .b(n_12950), .o(n_14091) );
na02f80 g557206 ( .a(n_11364), .b(x_in_4_6), .o(n_13343) );
no02f80 g557207 ( .a(n_11366), .b(n_11362), .o(n_11363) );
na02f80 g557208 ( .a(n_12114), .b(x_in_28_2), .o(n_13746) );
in01f80 g557209 ( .a(n_12538), .o(n_12539) );
no02f80 g557210 ( .a(n_12114), .b(x_in_28_2), .o(n_12538) );
na02f80 g557211 ( .a(n_10312), .b(n_10311), .o(n_10313) );
na02f80 g557212 ( .a(n_12112), .b(n_12111), .o(n_12113) );
no02f80 g557213 ( .a(n_10309), .b(n_10308), .o(n_10310) );
in01f80 g557214 ( .a(n_12110), .o(n_13265) );
na02f80 g557215 ( .a(n_11373), .b(n_1072), .o(n_12110) );
no02f80 g557216 ( .a(n_10306), .b(n_10305), .o(n_10307) );
no02f80 g557217 ( .a(n_12108), .b(n_12107), .o(n_12109) );
in01f80 g557218 ( .a(n_14595), .o(n_14596) );
na02f80 g557219 ( .a(n_12537), .b(n_8851), .o(n_14595) );
no02f80 g557220 ( .a(n_10982), .b(n_10979), .o(n_13286) );
na02f80 g557221 ( .a(n_12106), .b(n_10965), .o(n_13237) );
in01f80 g557222 ( .a(n_12535), .o(n_12536) );
na02f80 g557223 ( .a(n_12105), .b(n_12104), .o(n_12535) );
no02f80 g557224 ( .a(n_12105), .b(n_12104), .o(n_13718) );
na02f80 g557225 ( .a(n_10960), .b(n_12103), .o(n_13315) );
na02f80 g557226 ( .a(n_11361), .b(n_8347), .o(n_12852) );
no02f80 g557227 ( .a(n_11359), .b(x_in_7_10), .o(n_11360) );
no02f80 g557228 ( .a(n_12450), .b(n_13713), .o(n_12102) );
no02f80 g557229 ( .a(n_12101), .b(n_10955), .o(n_13294) );
no02f80 g557230 ( .a(n_12100), .b(n_10953), .o(n_13291) );
na02f80 g557231 ( .a(n_10068), .b(x_in_33_10), .o(n_11358) );
na02f80 g557232 ( .a(n_10067), .b(x_in_33_12), .o(n_11357) );
no02f80 g557233 ( .a(n_12561), .b(n_11593), .o(n_13748) );
na02f80 g557234 ( .a(n_12098), .b(n_12097), .o(n_12099) );
in01f80 g557235 ( .a(n_12948), .o(n_12949) );
na02f80 g557236 ( .a(n_12534), .b(n_11592), .o(n_12948) );
in01f80 g557237 ( .a(n_12532), .o(n_12533) );
na02f80 g557238 ( .a(n_10943), .b(n_12096), .o(n_12532) );
no02f80 g557239 ( .a(n_12095), .b(n_10941), .o(n_13297) );
na02f80 g557240 ( .a(n_11355), .b(n_11683), .o(n_11356) );
na02f80 g557241 ( .a(n_10967), .b(n_12094), .o(n_15239) );
na02f80 g557242 ( .a(n_10935), .b(n_10932), .o(n_13263) );
no02f80 g557243 ( .a(n_12092), .b(n_12091), .o(n_12093) );
na02f80 g557244 ( .a(n_11353), .b(x_in_5_12), .o(n_11354) );
no02f80 g557245 ( .a(n_12531), .b(n_11587), .o(n_14052) );
no02f80 g557246 ( .a(n_11351), .b(x_in_27_11), .o(n_11352) );
no02f80 g557247 ( .a(n_11349), .b(x_in_43_12), .o(n_11350) );
in01f80 g557248 ( .a(n_12831), .o(n_12090) );
na02f80 g557249 ( .a(n_11359), .b(n_8165), .o(n_12831) );
na02f80 g557250 ( .a(n_11347), .b(n_11346), .o(n_11348) );
na02f80 g557251 ( .a(n_12530), .b(n_11582), .o(n_13720) );
in01f80 g557252 ( .a(n_12529), .o(n_13710) );
no02f80 g557253 ( .a(n_12089), .b(x_in_15_10), .o(n_12529) );
in01f80 g557254 ( .a(n_12528), .o(n_13712) );
no02f80 g557255 ( .a(n_12088), .b(x_in_63_10), .o(n_12528) );
in01f80 g557256 ( .a(n_12527), .o(n_13711) );
no02f80 g557257 ( .a(n_12087), .b(x_in_23_10), .o(n_12527) );
in01f80 g557258 ( .a(n_12526), .o(n_13709) );
no02f80 g557259 ( .a(n_12086), .b(x_in_55_10), .o(n_12526) );
in01f80 g557260 ( .a(n_12525), .o(n_13708) );
no02f80 g557261 ( .a(n_12085), .b(x_in_47_10), .o(n_12525) );
in01f80 g557262 ( .a(n_12524), .o(n_13707) );
no02f80 g557263 ( .a(n_12084), .b(x_in_31_10), .o(n_12524) );
in01f80 g557264 ( .a(n_12522), .o(n_12523) );
na02f80 g557265 ( .a(n_10912), .b(n_12083), .o(n_12522) );
na02f80 g557266 ( .a(n_11344), .b(n_11343), .o(n_11345) );
na02f80 g557267 ( .a(n_10303), .b(n_10302), .o(n_10304) );
in01f80 g557268 ( .a(n_12081), .o(n_12082) );
no02f80 g557269 ( .a(n_10374), .b(n_7600), .o(n_12081) );
no02f80 g557270 ( .a(n_10375), .b(n_7601), .o(n_13258) );
no02f80 g557271 ( .a(n_12513), .b(x_in_56_1), .o(n_14200) );
na02f80 g557272 ( .a(n_12947), .b(x_in_24_1), .o(n_14618) );
no02f80 g557273 ( .a(n_12080), .b(n_13694), .o(n_13257) );
no02f80 g557274 ( .a(n_12521), .b(x_in_22_1), .o(n_15472) );
na02f80 g557275 ( .a(n_12515), .b(x_in_12_1), .o(n_15463) );
na02f80 g557276 ( .a(n_12521), .b(x_in_22_1), .o(n_15473) );
na02f80 g557277 ( .a(n_12520), .b(x_in_14_1), .o(n_15475) );
no02f80 g557278 ( .a(n_12520), .b(x_in_14_1), .o(n_15474) );
na02f80 g557279 ( .a(n_12519), .b(x_in_46_1), .o(n_15471) );
no02f80 g557280 ( .a(n_12519), .b(x_in_46_1), .o(n_15470) );
na02f80 g557281 ( .a(n_12518), .b(x_in_30_1), .o(n_15467) );
no02f80 g557282 ( .a(n_12518), .b(x_in_30_1), .o(n_15466) );
no02f80 g557283 ( .a(n_12517), .b(x_in_54_1), .o(n_15468) );
na02f80 g557284 ( .a(n_12517), .b(x_in_54_1), .o(n_15469) );
na02f80 g557285 ( .a(n_12516), .b(x_in_62_1), .o(n_15465) );
no02f80 g557286 ( .a(n_12516), .b(x_in_62_1), .o(n_15464) );
no02f80 g557287 ( .a(n_12515), .b(x_in_12_1), .o(n_15462) );
na02f80 g557288 ( .a(n_12514), .b(x_in_44_1), .o(n_15740) );
no02f80 g557289 ( .a(n_12514), .b(x_in_44_1), .o(n_15739) );
no02f80 g557290 ( .a(n_12947), .b(x_in_24_1), .o(n_14617) );
na02f80 g557291 ( .a(n_12513), .b(x_in_56_1), .o(n_14201) );
na02f80 g557292 ( .a(n_11578), .b(n_12512), .o(n_15198) );
in01f80 g557293 ( .a(n_12828), .o(n_12079) );
na02f80 g557294 ( .a(n_11351), .b(n_8513), .o(n_12828) );
no02f80 g557295 ( .a(n_12078), .b(n_10587), .o(n_13348) );
na02f80 g557296 ( .a(n_12511), .b(n_11576), .o(n_19004) );
in01f80 g557297 ( .a(n_11341), .o(n_11342) );
no02f80 g557298 ( .a(n_9595), .b(n_9449), .o(n_11341) );
no02f80 g557299 ( .a(n_9596), .b(n_8836), .o(n_12827) );
na02f80 g557300 ( .a(n_12510), .b(n_11574), .o(n_17104) );
na02f80 g557301 ( .a(n_10300), .b(n_10299), .o(n_10301) );
in01f80 g557302 ( .a(n_12077), .o(n_13242) );
na02f80 g557303 ( .a(n_11353), .b(n_5888), .o(n_12077) );
in01f80 g557304 ( .a(n_12826), .o(n_12076) );
na02f80 g557305 ( .a(n_11349), .b(n_7263), .o(n_12826) );
na02f80 g557306 ( .a(n_11572), .b(n_12509), .o(n_22911) );
no02f80 g557307 ( .a(n_12080), .b(n_12508), .o(n_13695) );
no02f80 g557308 ( .a(n_11564), .b(n_12507), .o(n_13739) );
in01f80 g557309 ( .a(n_12074), .o(n_12075) );
na02f80 g557310 ( .a(n_11340), .b(n_11339), .o(n_12074) );
no02f80 g557311 ( .a(n_11340), .b(n_11339), .o(n_13236) );
na02f80 g557312 ( .a(n_12506), .b(n_11562), .o(n_13723) );
no02f80 g557313 ( .a(n_12865), .b(n_12946), .o(n_14104) );
no02f80 g557314 ( .a(n_10297), .b(n_10296), .o(n_10298) );
na02f80 g557315 ( .a(n_12073), .b(n_10878), .o(n_13280) );
na02f80 g557316 ( .a(n_12505), .b(n_11560), .o(n_20819) );
na02f80 g557317 ( .a(n_10294), .b(n_10293), .o(n_10295) );
no02f80 g557318 ( .a(n_12504), .b(n_12286), .o(n_16598) );
in01f80 g557319 ( .a(n_11338), .o(n_12823) );
na02f80 g557320 ( .a(n_10292), .b(n_10291), .o(n_11338) );
no02f80 g557321 ( .a(n_11336), .b(n_11335), .o(n_11337) );
no02f80 g557322 ( .a(n_10292), .b(n_10291), .o(n_12825) );
na02f80 g557323 ( .a(n_11334), .b(n_11333), .o(n_13235) );
in01f80 g557324 ( .a(n_12071), .o(n_12072) );
no02f80 g557325 ( .a(n_11334), .b(n_11333), .o(n_12071) );
na02f80 g557326 ( .a(n_11331), .b(n_11330), .o(n_11332) );
no02f80 g557327 ( .a(n_11328), .b(n_11327), .o(n_11329) );
no02f80 g557328 ( .a(n_12217), .b(n_7854), .o(n_11326) );
na02f80 g557329 ( .a(n_11324), .b(n_11323), .o(n_11325) );
na02f80 g557330 ( .a(n_12069), .b(FE_OFN1232_n_12068), .o(n_12070) );
na02f80 g557331 ( .a(n_10289), .b(n_10288), .o(n_10290) );
no02f80 g557332 ( .a(n_11321), .b(n_11320), .o(n_11322) );
no02f80 g557333 ( .a(n_11318), .b(n_11317), .o(n_11319) );
no02f80 g557334 ( .a(n_11315), .b(n_11314), .o(n_11316) );
na02f80 g557335 ( .a(n_10859), .b(n_12067), .o(n_16279) );
na02f80 g557336 ( .a(n_11546), .b(n_12503), .o(n_13704) );
no02f80 g557337 ( .a(n_10286), .b(n_10285), .o(n_10287) );
na02f80 g557338 ( .a(n_11312), .b(n_11311), .o(n_11313) );
na02f80 g557339 ( .a(n_11309), .b(n_11308), .o(n_11310) );
no02f80 g557340 ( .a(n_11306), .b(n_11305), .o(n_11307) );
na02f80 g557341 ( .a(n_10283), .b(n_10282), .o(n_10284) );
na02f80 g557342 ( .a(n_10280), .b(n_10279), .o(n_10281) );
no02f80 g557343 ( .a(n_12066), .b(n_10854), .o(n_13326) );
na02f80 g557344 ( .a(n_11542), .b(n_12502), .o(n_13692) );
no02f80 g557345 ( .a(n_11540), .b(n_12501), .o(n_13683) );
na02f80 g557346 ( .a(n_11303), .b(n_11302), .o(n_11304) );
no02f80 g557347 ( .a(n_10277), .b(n_10276), .o(n_10278) );
in01f80 g557348 ( .a(n_15653), .o(n_12065) );
no02f80 g557349 ( .a(n_11301), .b(n_11300), .o(n_15653) );
no02f80 g557350 ( .a(n_11298), .b(n_11297), .o(n_11299) );
na02f80 g557351 ( .a(n_10274), .b(n_10273), .o(n_10275) );
no02f80 g557352 ( .a(n_10842), .b(n_12064), .o(n_21928) );
no02f80 g557353 ( .a(n_11537), .b(n_12500), .o(n_20024) );
na02f80 g557354 ( .a(n_10271), .b(n_10270), .o(n_10272) );
na02f80 g557355 ( .a(n_11295), .b(n_11294), .o(n_11296) );
na02f80 g557356 ( .a(n_10268), .b(n_10267), .o(n_10269) );
na02f80 g557357 ( .a(n_11292), .b(n_11291), .o(n_11293) );
na02f80 g557358 ( .a(n_11289), .b(n_11288), .o(n_11290) );
no02f80 g557359 ( .a(n_11286), .b(n_11285), .o(n_11287) );
na02f80 g557360 ( .a(n_10265), .b(n_10264), .o(n_10266) );
no02f80 g557361 ( .a(n_11283), .b(n_11282), .o(n_11284) );
no02f80 g557362 ( .a(n_10844), .b(n_12063), .o(n_13302) );
na02f80 g557363 ( .a(n_11280), .b(n_11279), .o(n_11281) );
no02f80 g557364 ( .a(n_11277), .b(n_11276), .o(n_11278) );
no02f80 g557365 ( .a(n_11274), .b(n_11273), .o(n_11275) );
no02f80 g557366 ( .a(n_11271), .b(n_11270), .o(n_11272) );
no02f80 g557367 ( .a(n_12279), .b(n_12499), .o(n_18039) );
no02f80 g557368 ( .a(n_10262), .b(n_10261), .o(n_10263) );
no02f80 g557369 ( .a(n_11268), .b(n_11267), .o(n_11269) );
no02f80 g557370 ( .a(n_10259), .b(n_10258), .o(n_10260) );
na02f80 g557371 ( .a(n_10256), .b(n_10255), .o(n_10257) );
na02f80 g557372 ( .a(n_11265), .b(n_11264), .o(n_11266) );
no02f80 g557373 ( .a(n_11535), .b(n_12498), .o(n_13757) );
na02f80 g557374 ( .a(n_10838), .b(n_12062), .o(n_18037) );
na02f80 g557375 ( .a(n_11262), .b(x_in_51_12), .o(n_11263) );
na02f80 g557376 ( .a(n_12647), .b(n_12646), .o(n_11261) );
no02f80 g557377 ( .a(n_11259), .b(n_11258), .o(n_11260) );
no02f80 g557378 ( .a(n_12497), .b(n_11533), .o(n_21555) );
na02f80 g557379 ( .a(n_11256), .b(n_11255), .o(n_11257) );
na02f80 g557380 ( .a(n_12173), .b(x_in_33_7), .o(n_10254) );
na02f80 g557381 ( .a(n_11253), .b(n_11252), .o(n_11254) );
na02f80 g557382 ( .a(n_10828), .b(n_12061), .o(n_20022) );
na02f80 g557383 ( .a(n_10251), .b(n_10250), .o(n_10252) );
na02f80 g557384 ( .a(n_12176), .b(x_in_33_9), .o(n_10253) );
na02f80 g557385 ( .a(n_11250), .b(x_in_33_8), .o(n_11251) );
na02f80 g557386 ( .a(n_11248), .b(x_in_33_6), .o(n_11249) );
na02f80 g557387 ( .a(n_10248), .b(n_10247), .o(n_10249) );
na02f80 g557388 ( .a(n_10826), .b(n_12060), .o(n_21923) );
no02f80 g557389 ( .a(n_11531), .b(n_12496), .o(n_16284) );
no02f80 g557390 ( .a(n_11246), .b(n_11245), .o(n_11247) );
no02f80 g557391 ( .a(n_11243), .b(n_11682), .o(n_11244) );
na02f80 g557392 ( .a(n_11241), .b(x_in_33_11), .o(n_11242) );
no02f80 g557393 ( .a(n_10245), .b(n_10244), .o(n_10246) );
na02f80 g557394 ( .a(n_11239), .b(n_11238), .o(n_11240) );
na02f80 g557395 ( .a(n_11236), .b(n_11235), .o(n_11237) );
no02f80 g557396 ( .a(n_11233), .b(n_11232), .o(n_11234) );
na02f80 g557397 ( .a(n_11230), .b(n_11229), .o(n_11231) );
na02f80 g557398 ( .a(n_11227), .b(n_11226), .o(n_11228) );
na02f80 g557399 ( .a(n_11224), .b(n_11223), .o(n_11225) );
no02f80 g557400 ( .a(n_11221), .b(n_11220), .o(n_11222) );
no02f80 g557401 ( .a(n_11218), .b(n_11217), .o(n_11219) );
no02f80 g557402 ( .a(n_11215), .b(n_11214), .o(n_11216) );
no02f80 g557403 ( .a(n_12617), .b(n_12616), .o(n_11213) );
na02f80 g557404 ( .a(n_12671), .b(n_12670), .o(n_11212) );
na02f80 g557405 ( .a(n_12058), .b(n_12057), .o(n_12059) );
no02f80 g557406 ( .a(n_10242), .b(n_10576), .o(n_10243) );
na02f80 g557407 ( .a(n_12945), .b(n_12278), .o(n_14113) );
na02f80 g557408 ( .a(n_10648), .b(n_12665), .o(n_12056) );
na02f80 g557409 ( .a(n_12054), .b(n_12053), .o(n_12055) );
no02f80 g557410 ( .a(n_11210), .b(n_11209), .o(n_11211) );
no02f80 g557411 ( .a(n_11207), .b(n_11206), .o(n_11208) );
no02f80 g557412 ( .a(n_12583), .b(n_12582), .o(n_11205) );
na02f80 g557413 ( .a(n_10240), .b(n_10239), .o(n_10241) );
no02f80 g557414 ( .a(n_12600), .b(n_12599), .o(n_11204) );
na02f80 g557415 ( .a(n_10816), .b(n_12052), .o(n_22572) );
na02f80 g557416 ( .a(n_10237), .b(n_10236), .o(n_10238) );
na02f80 g557417 ( .a(n_11202), .b(n_11201), .o(n_11203) );
no02f80 g557418 ( .a(n_12495), .b(n_11519), .o(n_22220) );
na02f80 g557419 ( .a(n_12597), .b(n_12596), .o(n_11200) );
na02f80 g557420 ( .a(n_11517), .b(n_12494), .o(n_14584) );
no02f80 g557421 ( .a(n_10235), .b(n_10234), .o(n_12819) );
in01f80 g557422 ( .a(n_11198), .o(n_11199) );
na02f80 g557423 ( .a(n_10235), .b(n_10234), .o(n_11198) );
no02f80 g557424 ( .a(n_11196), .b(n_11195), .o(n_11197) );
no02f80 g557425 ( .a(n_10808), .b(n_12051), .o(n_15258) );
na02f80 g557426 ( .a(n_10807), .b(n_12050), .o(n_20105) );
na02f80 g557427 ( .a(n_11193), .b(n_11192), .o(n_11194) );
no02f80 g557428 ( .a(n_10232), .b(n_10231), .o(n_10233) );
na02f80 g557429 ( .a(n_11515), .b(n_12493), .o(n_21139) );
na02f80 g557430 ( .a(n_11379), .b(n_11378), .o(n_11380) );
na02f80 g557431 ( .a(n_10802), .b(n_12049), .o(n_14077) );
na02f80 g557432 ( .a(n_11190), .b(n_11189), .o(n_11191) );
na02f80 g557433 ( .a(n_11187), .b(n_11186), .o(n_11188) );
na02f80 g557434 ( .a(n_10800), .b(n_11185), .o(n_21940) );
no02f80 g557435 ( .a(n_10229), .b(n_10228), .o(n_10230) );
na02f80 g557436 ( .a(n_12198), .b(n_10226), .o(n_10227) );
no02f80 g557437 ( .a(n_12198), .b(n_10224), .o(n_10225) );
na02f80 g557438 ( .a(n_11183), .b(n_11182), .o(n_11184) );
no02f80 g557439 ( .a(n_11513), .b(n_12492), .o(n_18679) );
na02f80 g557440 ( .a(n_12275), .b(n_12491), .o(n_19392) );
no02f80 g557441 ( .a(n_10796), .b(n_12048), .o(n_20824) );
na02f80 g557442 ( .a(n_12047), .b(n_11510), .o(n_21567) );
no02f80 g557443 ( .a(n_12205), .b(n_10222), .o(n_10223) );
no02f80 g557444 ( .a(n_12205), .b(n_10220), .o(n_10221) );
na02f80 g557445 ( .a(n_11180), .b(n_11179), .o(n_11181) );
no02f80 g557446 ( .a(n_11177), .b(n_11176), .o(n_11178) );
na02f80 g557447 ( .a(n_12199), .b(n_10218), .o(n_10219) );
no02f80 g557448 ( .a(n_12199), .b(n_10216), .o(n_10217) );
na02f80 g557449 ( .a(n_11507), .b(n_12490), .o(n_16632) );
no02f80 g557450 ( .a(n_12274), .b(n_12944), .o(n_17489) );
no02f80 g557451 ( .a(n_9874), .b(n_11175), .o(n_19386) );
no02f80 g557452 ( .a(n_12194), .b(n_10214), .o(n_10215) );
na02f80 g557453 ( .a(n_12194), .b(n_10212), .o(n_10213) );
na02f80 g557454 ( .a(n_12271), .b(n_12489), .o(n_17446) );
no02f80 g557455 ( .a(n_11505), .b(n_12488), .o(n_20468) );
no02f80 g557456 ( .a(n_10784), .b(n_12046), .o(n_17110) );
no02f80 g557457 ( .a(n_11503), .b(n_12487), .o(n_18348) );
no02f80 g557458 ( .a(n_12183), .b(n_10779), .o(n_10327) );
na02f80 g557459 ( .a(n_12183), .b(n_12697), .o(n_10211) );
no02f80 g557460 ( .a(n_11500), .b(n_12486), .o(n_16882) );
na02f80 g557461 ( .a(n_12045), .b(n_13676), .o(n_13099) );
na02f80 g557462 ( .a(n_11498), .b(n_12485), .o(n_17805) );
in01f80 g557463 ( .a(n_12483), .o(n_12484) );
no02f80 g557464 ( .a(n_11387), .b(n_9823), .o(n_12483) );
no02f80 g557465 ( .a(n_11388), .b(n_9824), .o(n_13674) );
na02f80 g557466 ( .a(n_12043), .b(n_12042), .o(n_12044) );
na02f80 g557467 ( .a(n_11486), .b(n_12482), .o(n_20870) );
no02f80 g557468 ( .a(n_11428), .b(n_12481), .o(n_21974) );
na02f80 g557469 ( .a(n_11439), .b(n_12480), .o(n_22926) );
in01f80 g557470 ( .a(n_12040), .o(n_12041) );
no02f80 g557471 ( .a(n_10380), .b(n_7580), .o(n_12040) );
no02f80 g557472 ( .a(n_11482), .b(n_12479), .o(n_15634) );
oa12f80 g557473 ( .a(n_11145), .b(n_425), .c(FE_OFN355_n_4860), .o(n_11174) );
na02f80 g557474 ( .a(n_9867), .b(n_11173), .o(n_18393) );
no02f80 g557475 ( .a(n_12185), .b(FE_OFN480_n_12184), .o(n_10210) );
no02f80 g557476 ( .a(n_11171), .b(FE_OFN478_n_11170), .o(n_11172) );
no02f80 g557477 ( .a(n_9697), .b(n_11168), .o(n_11169) );
no02f80 g557478 ( .a(n_10208), .b(n_10207), .o(n_10209) );
na02f80 g557479 ( .a(n_11375), .b(n_10205), .o(n_10206) );
na02f80 g557480 ( .a(n_11161), .b(n_11160), .o(n_13113) );
no02f80 g557481 ( .a(n_12639), .b(FE_OFN484_n_12038), .o(n_12039) );
no02f80 g557482 ( .a(n_11426), .b(n_12478), .o(n_19716) );
no02f80 g557483 ( .a(n_12036), .b(n_12351), .o(n_12037) );
no02f80 g557484 ( .a(n_9694), .b(n_11166), .o(n_11167) );
na02f80 g557485 ( .a(n_12191), .b(n_11168), .o(n_10204) );
no02f80 g557486 ( .a(n_11859), .b(n_11858), .o(n_13661) );
in01f80 g557487 ( .a(n_12476), .o(n_12477) );
na02f80 g557488 ( .a(n_11400), .b(n_7584), .o(n_12476) );
na02f80 g557489 ( .a(n_12187), .b(FE_OFN1254_n_12186), .o(n_10203) );
na02f80 g557490 ( .a(n_11401), .b(n_7585), .o(n_13673) );
na02f80 g557491 ( .a(n_11488), .b(n_12475), .o(n_17154) );
in01f80 g557492 ( .a(n_12473), .o(n_12474) );
no02f80 g557493 ( .a(n_11398), .b(n_8940), .o(n_12473) );
no02f80 g557494 ( .a(n_11399), .b(n_8939), .o(n_13659) );
na02f80 g557495 ( .a(n_12034), .b(n_12033), .o(n_12035) );
no02f80 g557496 ( .a(n_12031), .b(n_12030), .o(n_12032) );
no02f80 g557497 ( .a(n_12028), .b(n_12368), .o(n_12029) );
na02f80 g557498 ( .a(n_12026), .b(n_12025), .o(n_12027) );
na02f80 g557499 ( .a(n_11164), .b(n_11163), .o(n_11165) );
no02f80 g557500 ( .a(n_12023), .b(n_12022), .o(n_12024) );
no02f80 g557501 ( .a(n_12148), .b(n_11166), .o(n_10202) );
no02f80 g557502 ( .a(n_12020), .b(n_12019), .o(n_12021) );
na02f80 g557503 ( .a(n_12251), .b(n_12472), .o(n_20856) );
na02f80 g557504 ( .a(n_12674), .b(n_12673), .o(n_11162) );
na02f80 g557505 ( .a(n_12017), .b(FE_OFN1196_n_12016), .o(n_12018) );
na02f80 g557506 ( .a(n_10672), .b(n_12015), .o(n_17122) );
na02f80 g557507 ( .a(n_12013), .b(n_12012), .o(n_12014) );
in01f80 g557508 ( .a(n_12470), .o(n_12471) );
no02f80 g557509 ( .a(n_12011), .b(n_12010), .o(n_12470) );
na02f80 g557510 ( .a(n_12011), .b(n_12010), .o(n_13662) );
no02f80 g557511 ( .a(n_12008), .b(n_12007), .o(n_12009) );
na02f80 g557512 ( .a(n_12005), .b(n_12004), .o(n_12006) );
no02f80 g557513 ( .a(n_12002), .b(n_12001), .o(n_12003) );
no02f80 g557514 ( .a(n_10528), .b(n_10142), .o(n_12000) );
no02f80 g557515 ( .a(n_11998), .b(n_11997), .o(n_11999) );
na02f80 g557516 ( .a(n_11995), .b(n_11994), .o(n_11996) );
na02f80 g557517 ( .a(n_11992), .b(n_11991), .o(n_11993) );
no02f80 g557518 ( .a(n_10560), .b(n_10139), .o(n_11990) );
no02f80 g557519 ( .a(n_11941), .b(n_11940), .o(n_13656) );
no02f80 g557520 ( .a(n_12943), .b(n_12269), .o(n_21188) );
na02f80 g557521 ( .a(n_12135), .b(n_11484), .o(n_14062) );
in01f80 g557522 ( .a(n_11988), .o(n_11989) );
no02f80 g557523 ( .a(n_11161), .b(n_11160), .o(n_11988) );
no02f80 g557524 ( .a(n_12155), .b(n_12154), .o(n_10201) );
no02f80 g557525 ( .a(n_11986), .b(n_11985), .o(n_11987) );
na02f80 g557526 ( .a(n_11983), .b(n_11982), .o(n_11984) );
no02f80 g557527 ( .a(n_11980), .b(n_11979), .o(n_11981) );
na02f80 g557528 ( .a(n_11977), .b(n_11976), .o(n_11978) );
na02f80 g557529 ( .a(n_11974), .b(n_11973), .o(n_11975) );
no02f80 g557530 ( .a(n_11971), .b(n_12318), .o(n_11972) );
na02f80 g557531 ( .a(n_11969), .b(n_11968), .o(n_11970) );
no02f80 g557532 ( .a(n_10509), .b(FE_OFN576_n_10136), .o(n_11967) );
no02f80 g557533 ( .a(n_11158), .b(n_11157), .o(n_11159) );
na02f80 g557534 ( .a(n_11965), .b(n_11964), .o(n_11966) );
no02f80 g557535 ( .a(n_11962), .b(n_11961), .o(n_11963) );
na02f80 g557536 ( .a(n_11959), .b(n_11958), .o(n_11960) );
no02f80 g557537 ( .a(n_11956), .b(n_11955), .o(n_11957) );
na02f80 g557538 ( .a(n_11953), .b(n_11952), .o(n_11954) );
no02f80 g557539 ( .a(n_11950), .b(n_11949), .o(n_11951) );
no02f80 g557540 ( .a(n_11947), .b(n_11946), .o(n_11948) );
na02f80 g557541 ( .a(n_11944), .b(n_11943), .o(n_11945) );
in01f80 g557542 ( .a(n_12468), .o(n_12469) );
na02f80 g557543 ( .a(n_11402), .b(n_8256), .o(n_12468) );
no02f80 g557544 ( .a(n_10484), .b(n_10133), .o(n_11942) );
no02f80 g557545 ( .a(n_12265), .b(n_12942), .o(n_24546) );
in01f80 g557546 ( .a(n_12466), .o(n_12467) );
na02f80 g557547 ( .a(n_11941), .b(n_11940), .o(n_12466) );
in01f80 g557548 ( .a(n_11938), .o(n_11939) );
no02f80 g557549 ( .a(n_10480), .b(n_9446), .o(n_11938) );
no02f80 g557550 ( .a(n_10481), .b(n_9447), .o(n_13180) );
na02f80 g557551 ( .a(n_11155), .b(n_11154), .o(n_11156) );
na02f80 g557552 ( .a(n_12263), .b(n_12465), .o(n_24505) );
na02f80 g557553 ( .a(n_12097), .b(n_12464), .o(n_14511) );
no02f80 g557554 ( .a(n_10749), .b(n_11937), .o(n_19010) );
no02f80 g557555 ( .a(n_11935), .b(n_12367), .o(n_11936) );
in01f80 g557556 ( .a(n_12462), .o(n_12463) );
no02f80 g557557 ( .a(n_11394), .b(n_6596), .o(n_12462) );
no02f80 g557558 ( .a(n_11395), .b(n_6597), .o(n_13641) );
ao22s80 g557559 ( .a(n_11153), .b(n_4784), .c(n_5908), .d(n_5907), .o(n_15222) );
na02f80 g557560 ( .a(n_11933), .b(n_12373), .o(n_11934) );
na02f80 g557561 ( .a(n_11931), .b(n_11930), .o(n_11932) );
no02f80 g557562 ( .a(n_11928), .b(n_11927), .o(n_11929) );
no02f80 g557563 ( .a(n_11925), .b(n_11924), .o(n_11926) );
no02f80 g557564 ( .a(n_11922), .b(n_11921), .o(n_11923) );
na02f80 g557565 ( .a(n_11919), .b(n_11918), .o(n_11920) );
no02f80 g557566 ( .a(n_11916), .b(n_11915), .o(n_11917) );
no02f80 g557567 ( .a(n_11913), .b(n_11912), .o(n_11914) );
na02f80 g557568 ( .a(n_11910), .b(n_11909), .o(n_11911) );
na02f80 g557569 ( .a(n_11907), .b(n_11906), .o(n_11908) );
na02f80 g557570 ( .a(n_11904), .b(n_11903), .o(n_11905) );
na02f80 g557571 ( .a(n_11151), .b(n_11150), .o(n_11152) );
no02f80 g557572 ( .a(n_11901), .b(n_11900), .o(n_11902) );
no02f80 g557573 ( .a(n_10450), .b(n_11031), .o(n_11899) );
na02f80 g557574 ( .a(n_11849), .b(n_11848), .o(n_13640) );
na02f80 g557575 ( .a(n_11897), .b(FE_OFN1192_n_11896), .o(n_11898) );
no02f80 g557576 ( .a(n_11894), .b(n_11893), .o(n_11895) );
na02f80 g557577 ( .a(n_11891), .b(FE_OFN1101_n_12369), .o(n_11892) );
no02f80 g557578 ( .a(n_11889), .b(n_12372), .o(n_11890) );
na02f80 g557579 ( .a(n_11887), .b(n_12371), .o(n_11888) );
no02f80 g557580 ( .a(n_11885), .b(n_12370), .o(n_11886) );
na02f80 g557581 ( .a(n_11883), .b(n_11882), .o(n_11884) );
no02f80 g557582 ( .a(n_10199), .b(FE_OFN785_n_10198), .o(n_10200) );
no02f80 g557583 ( .a(n_11880), .b(n_11879), .o(n_11881) );
na02f80 g557584 ( .a(n_11877), .b(n_11876), .o(n_11878) );
na02f80 g557585 ( .a(n_11874), .b(n_11873), .o(n_11875) );
na02f80 g557586 ( .a(n_11871), .b(n_11870), .o(n_11872) );
no02f80 g557587 ( .a(n_10360), .b(n_11028), .o(n_11869) );
no02f80 g557588 ( .a(n_12461), .b(n_11474), .o(n_14507) );
na02f80 g557589 ( .a(n_11476), .b(n_12460), .o(n_15609) );
na02f80 g557590 ( .a(n_11478), .b(n_12459), .o(n_19341) );
no02f80 g557591 ( .a(n_11480), .b(n_12458), .o(n_20056) );
na02f80 g557592 ( .a(n_11867), .b(n_11866), .o(n_11868) );
na02f80 g557593 ( .a(n_11864), .b(n_11863), .o(n_11865) );
na02f80 g557594 ( .a(n_12202), .b(FE_OFN1186_n_12201), .o(n_10197) );
na02f80 g557595 ( .a(n_11861), .b(n_11860), .o(n_11862) );
no02f80 g557596 ( .a(n_9692), .b(n_11148), .o(n_11149) );
no02f80 g557597 ( .a(n_10195), .b(n_10194), .o(n_10196) );
no02f80 g557598 ( .a(n_11420), .b(n_12457), .o(n_16323) );
na02f80 g557599 ( .a(n_12455), .b(n_14533), .o(n_12456) );
na02f80 g557600 ( .a(n_12455), .b(n_14535), .o(n_14022) );
ao12f80 g557601 ( .a(n_12832), .b(n_10062), .c(n_10061), .o(n_12843) );
no03m80 g557602 ( .a(n_7940), .b(n_11583), .c(FE_OFN1244_n_12940), .o(n_12941) );
na02f80 g557603 ( .a(n_12200), .b(n_11148), .o(n_10193) );
in01f80 g557604 ( .a(n_12453), .o(n_12454) );
na02f80 g557605 ( .a(n_11859), .b(n_11858), .o(n_12453) );
no02f80 g557606 ( .a(n_10191), .b(n_11070), .o(n_10192) );
no02f80 g557607 ( .a(n_11468), .b(n_11857), .o(n_26100) );
in01f80 g557608 ( .a(n_11856), .o(n_13465) );
no02f80 g557609 ( .a(n_11147), .b(n_11823), .o(n_11856) );
na02f80 g557610 ( .a(n_11119), .b(n_11118), .o(n_13111) );
na02f80 g557611 ( .a(n_11467), .b(n_11465), .o(n_23867) );
no02f80 g557612 ( .a(n_11854), .b(n_11853), .o(n_11855) );
oa12f80 g557613 ( .a(n_11145), .b(n_195), .c(FE_OFN1112_rst), .o(n_11146) );
na02f80 g557614 ( .a(n_11851), .b(n_11850), .o(n_11852) );
in01f80 g557615 ( .a(n_12451), .o(n_12452) );
no02f80 g557616 ( .a(n_11849), .b(n_11848), .o(n_12451) );
no02f80 g557617 ( .a(n_12450), .b(n_12449), .o(n_13714) );
na02f80 g557618 ( .a(n_10711), .b(n_11847), .o(n_13239) );
in01f80 g557619 ( .a(n_11143), .o(n_11144) );
no02f80 g557620 ( .a(n_9701), .b(n_9420), .o(n_11143) );
no02f80 g557621 ( .a(n_9702), .b(n_9421), .o(n_12732) );
na02f80 g557622 ( .a(n_11845), .b(n_11844), .o(n_11846) );
na02f80 g557623 ( .a(n_11842), .b(n_11841), .o(n_11843) );
no02f80 g557624 ( .a(n_12938), .b(n_12937), .o(n_12939) );
na02f80 g557625 ( .a(n_11839), .b(n_11838), .o(n_11840) );
no02f80 g557626 ( .a(n_11141), .b(n_11140), .o(n_11142) );
no02f80 g557627 ( .a(n_11138), .b(n_11137), .o(n_11139) );
na02f80 g557628 ( .a(n_11135), .b(n_11134), .o(n_11136) );
no02f80 g557629 ( .a(n_11132), .b(n_11131), .o(n_11133) );
no02f80 g557630 ( .a(n_11777), .b(n_11776), .o(n_13627) );
no02f80 g557631 ( .a(n_11460), .b(n_12448), .o(n_14024) );
na02f80 g557632 ( .a(n_11837), .b(n_10660), .o(n_13467) );
no02f80 g557633 ( .a(n_11835), .b(n_12344), .o(n_11836) );
na02f80 g557634 ( .a(n_11833), .b(n_11832), .o(n_11834) );
na02f80 g557635 ( .a(n_11129), .b(n_12627), .o(n_11130) );
na02f80 g557636 ( .a(n_11831), .b(n_11830), .o(n_19002) );
na02f80 g557637 ( .a(n_11127), .b(n_6029), .o(n_11128) );
no02f80 g557638 ( .a(n_11125), .b(n_10696), .o(n_11126) );
na02f80 g557639 ( .a(n_12447), .b(n_11457), .o(n_14055) );
no02f80 g557640 ( .a(n_11455), .b(n_12446), .o(n_14986) );
in01f80 g557641 ( .a(n_11828), .o(n_11829) );
na02f80 g557642 ( .a(n_10570), .b(n_10331), .o(n_11828) );
no02f80 g557643 ( .a(n_11827), .b(n_11826), .o(n_17162) );
na02f80 g557644 ( .a(n_11127), .b(n_11825), .o(n_16344) );
na02f80 g557645 ( .a(n_12445), .b(n_11453), .o(n_15986) );
na02f80 g557646 ( .a(n_10571), .b(n_10332), .o(n_13134) );
no02f80 g557647 ( .a(n_13007), .b(n_11823), .o(n_11824) );
na02f80 g557648 ( .a(n_13004), .b(FE_OFN1198_n_13003), .o(n_11822) );
no02f80 g557649 ( .a(n_13002), .b(n_13001), .o(n_11821) );
na02f80 g557650 ( .a(n_13091), .b(FE_OFN1190_n_13090), .o(n_11820) );
no02f80 g557651 ( .a(n_10619), .b(n_11819), .o(n_23882) );
in01f80 g557652 ( .a(n_11817), .o(n_11818) );
no02f80 g557653 ( .a(n_10382), .b(n_8552), .o(n_11817) );
no02f80 g557654 ( .a(n_10383), .b(n_8553), .o(n_13121) );
no02f80 g557655 ( .a(n_11815), .b(n_11814), .o(n_11816) );
no02f80 g557656 ( .a(n_10189), .b(n_10188), .o(n_10190) );
no02f80 g557657 ( .a(n_11124), .b(n_11123), .o(n_13120) );
in01f80 g557658 ( .a(n_11812), .o(n_11813) );
na02f80 g557659 ( .a(n_11124), .b(n_11123), .o(n_11812) );
no02f80 g557660 ( .a(n_11121), .b(n_11120), .o(n_11122) );
no02f80 g557661 ( .a(n_10381), .b(n_7579), .o(n_13112) );
in01f80 g557662 ( .a(n_11810), .o(n_11811) );
no02f80 g557663 ( .a(n_11119), .b(n_11118), .o(n_11810) );
na02f80 g557664 ( .a(n_11116), .b(n_11115), .o(n_11117) );
in01f80 g557665 ( .a(n_11808), .o(n_11809) );
no02f80 g557666 ( .a(n_10378), .b(n_8255), .o(n_11808) );
no02f80 g557667 ( .a(n_10674), .b(n_11807), .o(n_16307) );
no02f80 g557668 ( .a(n_10379), .b(n_8254), .o(n_13110) );
in01f80 g557669 ( .a(n_11805), .o(n_11806) );
na02f80 g557670 ( .a(n_10376), .b(n_8820), .o(n_11805) );
no02f80 g557671 ( .a(n_10694), .b(n_11804), .o(n_15252) );
no02f80 g557672 ( .a(n_10770), .b(n_11803), .o(n_18051) );
na02f80 g557673 ( .a(n_11802), .b(n_10676), .o(n_15224) );
no02f80 g557674 ( .a(n_12443), .b(n_12442), .o(n_12444) );
na02f80 g557675 ( .a(n_10670), .b(n_11801), .o(n_19023) );
no02f80 g557676 ( .a(n_10682), .b(n_11800), .o(n_19682) );
na02f80 g557677 ( .a(n_10377), .b(n_8821), .o(n_13209) );
na02f80 g557678 ( .a(n_10664), .b(n_11799), .o(n_20836) );
no02f80 g557679 ( .a(n_10662), .b(n_11798), .o(n_21938) );
oa12f80 g557680 ( .a(n_12118), .b(n_14491), .c(n_12117), .o(n_14502) );
na02f80 g557681 ( .a(n_11447), .b(n_12441), .o(n_22891) );
in01f80 g557682 ( .a(n_11796), .o(n_11797) );
na02f80 g557683 ( .a(n_10371), .b(n_8938), .o(n_11796) );
na02f80 g557684 ( .a(n_10372), .b(n_8937), .o(n_13114) );
na02f80 g557685 ( .a(n_13521), .b(FE_OFN482_n_13520), .o(n_12440) );
no02f80 g557686 ( .a(n_10422), .b(n_10145), .o(n_11795) );
in01f80 g557687 ( .a(n_17357), .o(n_11114) );
oa12f80 g557688 ( .a(n_8418), .b(n_11521), .c(n_9566), .o(n_17357) );
in01f80 g557689 ( .a(n_12935), .o(n_12936) );
no02f80 g557690 ( .a(n_12243), .b(n_8947), .o(n_12935) );
no02f80 g557691 ( .a(n_12244), .b(n_8946), .o(n_14085) );
no02f80 g557692 ( .a(n_10728), .b(n_11794), .o(n_14984) );
na02f80 g557693 ( .a(n_10658), .b(n_11793), .o(n_15984) );
no02f80 g557694 ( .a(n_10760), .b(n_11792), .o(n_16880) );
na02f80 g557695 ( .a(n_10656), .b(n_11791), .o(n_17803) );
no02f80 g557696 ( .a(n_11491), .b(n_11790), .o(n_18677) );
no02f80 g557697 ( .a(n_11112), .b(n_11111), .o(n_11113) );
na02f80 g557698 ( .a(n_11445), .b(n_11789), .o(n_19390) );
no02f80 g557699 ( .a(n_10653), .b(n_11788), .o(n_20466) );
na02f80 g557700 ( .a(n_10651), .b(n_11787), .o(n_21565) );
no02f80 g557701 ( .a(n_11443), .b(n_12439), .o(n_22580) );
in01f80 g557702 ( .a(n_11785), .o(n_11786) );
no02f80 g557703 ( .a(n_10365), .b(n_8935), .o(n_11785) );
no02f80 g557704 ( .a(n_11109), .b(FE_OFN1204_n_11679), .o(n_11110) );
na02f80 g557705 ( .a(n_11107), .b(n_11106), .o(n_11108) );
na02f80 g557706 ( .a(n_12161), .b(n_12160), .o(n_10187) );
no02f80 g557707 ( .a(n_12159), .b(FE_OFN779_n_12158), .o(n_10186) );
no02f80 g557708 ( .a(n_10184), .b(FE_OFN1226_n_10183), .o(n_10185) );
na02f80 g557709 ( .a(n_12977), .b(n_12978), .o(n_11784) );
no02f80 g557710 ( .a(n_12598), .b(n_11782), .o(n_11783) );
no02f80 g557711 ( .a(n_11104), .b(n_11103), .o(n_11105) );
oa12f80 g557712 ( .a(n_11102), .b(n_10778), .c(n_10777), .o(n_12850) );
na02f80 g557713 ( .a(n_12258), .b(n_12934), .o(n_15237) );
no02f80 g557714 ( .a(n_12256), .b(n_12933), .o(n_16327) );
na02f80 g557715 ( .a(n_11433), .b(n_12438), .o(n_17142) );
no02f80 g557716 ( .a(n_10366), .b(n_8934), .o(n_13109) );
no02f80 g557717 ( .a(n_12261), .b(n_12437), .o(n_18069) );
na02f80 g557718 ( .a(n_12253), .b(n_12436), .o(n_19045) );
no02f80 g557719 ( .a(n_10642), .b(n_11781), .o(n_19702) );
no02f80 g557720 ( .a(n_12249), .b(n_12932), .o(n_21960) );
no02f80 g557721 ( .a(n_10638), .b(n_11780), .o(n_23847) );
in01f80 g557722 ( .a(n_11778), .o(n_11779) );
na02f80 g557723 ( .a(n_10356), .b(n_9394), .o(n_11778) );
na02f80 g557724 ( .a(n_10357), .b(n_9395), .o(n_13108) );
in01f80 g557725 ( .a(n_12434), .o(n_12435) );
na02f80 g557726 ( .a(n_11777), .b(n_11776), .o(n_12434) );
no02f80 g557727 ( .a(n_12431), .b(FE_OFN642_n_12432), .o(n_12433) );
oa12f80 g557728 ( .a(n_11101), .b(n_10848), .c(n_10847), .o(n_12848) );
no02f80 g557729 ( .a(n_12969), .b(n_12968), .o(n_11775) );
na02f80 g557730 ( .a(n_12576), .b(n_12575), .o(n_11100) );
na02f80 g557731 ( .a(n_11098), .b(n_11097), .o(n_11099) );
na02f80 g557732 ( .a(n_11403), .b(n_8257), .o(n_13614) );
no02f80 g557733 ( .a(n_12146), .b(n_12147), .o(n_10182) );
na02f80 g557734 ( .a(n_11095), .b(n_11094), .o(n_11096) );
na02f80 g557735 ( .a(n_12164), .b(n_12163), .o(n_10181) );
na02f80 g557736 ( .a(n_11092), .b(n_11091), .o(n_11093) );
na02f80 g557737 ( .a(n_11376), .b(n_10179), .o(n_10180) );
no02f80 g557738 ( .a(n_12431), .b(n_14524), .o(n_14050) );
no02f80 g557739 ( .a(n_11422), .b(n_12430), .o(n_18083) );
na02f80 g557740 ( .a(n_11424), .b(n_12429), .o(n_19041) );
oa12f80 g557741 ( .a(n_10177), .b(n_11090), .c(n_10178), .o(n_12845) );
in01f80 g557742 ( .a(n_11088), .o(n_11089) );
no03m80 g557743 ( .a(n_10178), .b(n_11090), .c(n_10177), .o(n_11088) );
in01f80 g557744 ( .a(n_11086), .o(n_11087) );
no03m80 g557745 ( .a(n_10176), .b(n_14432), .c(n_10175), .o(n_11086) );
in01f80 g557746 ( .a(n_10174), .o(n_12856) );
oa12f80 g557747 ( .a(n_2755), .b(n_9366), .c(n_2186), .o(n_10174) );
in01f80 g557748 ( .a(n_10173), .o(n_12858) );
oa12f80 g557749 ( .a(n_3065), .b(n_9361), .c(n_2192), .o(n_10173) );
in01f80 g557750 ( .a(n_11084), .o(n_11085) );
no03m80 g557751 ( .a(n_10172), .b(n_14323), .c(n_10171), .o(n_11084) );
oa12f80 g557752 ( .a(n_11082), .b(n_14389), .c(n_11083), .o(n_13334) );
in01f80 g557753 ( .a(n_11773), .o(n_11774) );
no03m80 g557754 ( .a(n_11083), .b(n_14389), .c(n_11082), .o(n_11773) );
in01f80 g557755 ( .a(n_11080), .o(n_11081) );
no03m80 g557756 ( .a(n_10170), .b(n_14332), .c(n_10169), .o(n_11080) );
oa12f80 g557757 ( .a(n_10169), .b(n_14332), .c(n_10170), .o(n_12844) );
in01f80 g557758 ( .a(n_11079), .o(n_13366) );
oa12f80 g557759 ( .a(n_9563), .b(n_10168), .c(n_8402), .o(n_11079) );
ao12f80 g557760 ( .a(n_11078), .b(n_7878), .c(n_7877), .o(n_12835) );
oa12f80 g557761 ( .a(n_10175), .b(n_14432), .c(n_10176), .o(n_12841) );
in01f80 g557762 ( .a(n_11077), .o(n_13370) );
oa12f80 g557763 ( .a(n_9200), .b(n_10167), .c(n_7956), .o(n_11077) );
oa12f80 g557764 ( .a(n_10171), .b(n_14323), .c(n_10172), .o(n_12846) );
oa12f80 g557765 ( .a(n_11075), .b(n_103), .c(FE_OFN355_n_4860), .o(n_11076) );
oa12f80 g557766 ( .a(n_11075), .b(n_1375), .c(FE_OFN127_n_27449), .o(n_11074) );
oa12f80 g557767 ( .a(n_11770), .b(n_498), .c(FE_OFN330_n_4860), .o(n_11772) );
oa12f80 g557768 ( .a(n_11770), .b(n_1189), .c(FE_OFN330_n_4860), .o(n_11771) );
ao12f80 g557769 ( .a(n_9042), .b(n_8809), .c(n_6032), .o(n_11377) );
oa12f80 g557770 ( .a(n_9209), .b(n_9208), .c(n_9207), .o(n_23956) );
in01f80 g557771 ( .a(n_11073), .o(n_13377) );
ao12f80 g557772 ( .a(n_5269), .b(n_10166), .c(n_5268), .o(n_11073) );
oa12f80 g557773 ( .a(n_12245), .b(n_9428), .c(n_9429), .o(n_12931) );
ao12f80 g557774 ( .a(n_11769), .b(n_8317), .c(n_8316), .o(n_13278) );
ao12f80 g557775 ( .a(n_9785), .b(n_10559), .c(n_10558), .o(n_11072) );
ao12f80 g557776 ( .a(n_10933), .b(n_10708), .c(n_10707), .o(n_11768) );
in01f80 g557777 ( .a(n_12427), .o(n_12428) );
oa12f80 g557778 ( .a(n_10597), .b(n_10530), .c(n_10529), .o(n_12427) );
in01f80 g557779 ( .a(n_11766), .o(n_11767) );
oa22f80 g557780 ( .a(n_9165), .b(n_11991), .c(n_10420), .d(n_10421), .o(n_11766) );
in01f80 g557781 ( .a(n_11764), .o(n_11765) );
oa22f80 g557782 ( .a(n_9169), .b(n_11943), .c(n_10488), .d(n_10489), .o(n_11764) );
in01f80 g557783 ( .a(n_11762), .o(n_11763) );
oa22f80 g557784 ( .a(n_9159), .b(n_11906), .c(n_10454), .d(n_10455), .o(n_11762) );
in01f80 g557785 ( .a(n_11760), .o(n_11761) );
oa22f80 g557786 ( .a(n_9162), .b(n_11873), .c(n_10433), .d(n_10434), .o(n_11760) );
ao12f80 g557787 ( .a(n_10596), .b(n_10388), .c(n_10385), .o(n_14235) );
oa12f80 g557788 ( .a(n_10855), .b(n_9976), .c(n_9975), .o(n_12830) );
oa12f80 g557789 ( .a(n_11861), .b(n_14466), .c(n_11860), .o(n_14807) );
no02f80 g557790 ( .a(n_10834), .b(n_9933), .o(n_22181) );
oa22f80 g557791 ( .a(n_11071), .b(n_3994), .c(n_5282), .d(x_in_33_4), .o(n_15515) );
in01f80 g557792 ( .a(n_12929), .o(n_12930) );
na03f80 g557793 ( .a(n_6558), .b(n_12426), .c(n_12425), .o(n_12929) );
ao12f80 g557794 ( .a(n_10165), .b(n_9983), .c(n_9982), .o(n_12239) );
in01f80 g557795 ( .a(n_11758), .o(n_11759) );
ao12f80 g557796 ( .a(n_9777), .b(n_9614), .c(n_9612), .o(n_11758) );
in01f80 g557797 ( .a(n_12242), .o(n_10164) );
oa12f80 g557798 ( .a(n_5688), .b(n_9365), .c(n_4770), .o(n_12242) );
in01f80 g557799 ( .a(n_11756), .o(n_11757) );
ao22s80 g557800 ( .a(n_9119), .b(n_9244), .c(n_11070), .d(x_in_49_14), .o(n_11756) );
in01f80 g557801 ( .a(n_10162), .o(n_10163) );
oa22f80 g557802 ( .a(n_8172), .b(n_9279), .c(n_9278), .d(n_10264), .o(n_10162) );
in01f80 g557803 ( .a(n_11068), .o(n_11069) );
oa22f80 g557804 ( .a(n_8716), .b(n_9687), .c(n_9686), .d(n_11291), .o(n_11068) );
in01f80 g557805 ( .a(n_10160), .o(n_10161) );
oa22f80 g557806 ( .a(n_8170), .b(n_9216), .c(n_9215), .d(n_10270), .o(n_10160) );
in01f80 g557807 ( .a(n_11754), .o(n_11755) );
ao12f80 g557808 ( .a(n_9771), .b(n_9607), .c(n_9608), .o(n_11754) );
in01f80 g557809 ( .a(n_11752), .o(n_11753) );
ao12f80 g557810 ( .a(n_9720), .b(n_9648), .c(n_9646), .o(n_11752) );
in01f80 g557811 ( .a(n_11066), .o(n_11067) );
ao22s80 g557812 ( .a(n_10159), .b(n_7805), .c(n_12811), .d(x_in_23_10), .o(n_11066) );
in01f80 g557813 ( .a(n_11064), .o(n_11065) );
ao22s80 g557814 ( .a(n_10158), .b(n_7806), .c(FE_OFN987_n_12804), .d(x_in_55_10), .o(n_11064) );
in01f80 g557815 ( .a(n_11062), .o(n_11063) );
ao22s80 g557816 ( .a(n_10157), .b(n_8343), .c(FE_OFN572_n_12800), .d(x_in_15_10), .o(n_11062) );
in01f80 g557817 ( .a(n_11060), .o(n_11061) );
ao22s80 g557818 ( .a(n_10156), .b(n_7801), .c(n_12787), .d(x_in_47_10), .o(n_11060) );
in01f80 g557819 ( .a(n_11058), .o(n_11059) );
ao22s80 g557820 ( .a(n_10155), .b(n_7804), .c(FE_OFN1216_n_12761), .d(x_in_31_10), .o(n_11058) );
in01f80 g557821 ( .a(n_11056), .o(n_11057) );
ao22s80 g557822 ( .a(n_10154), .b(n_7798), .c(FE_OFN1276_n_12754), .d(x_in_63_10), .o(n_11056) );
oa22f80 g557823 ( .a(n_14112), .b(n_7943), .c(n_9206), .d(n_9205), .o(n_16000) );
in01f80 g557824 ( .a(n_15708), .o(n_11751) );
oa12f80 g557825 ( .a(n_8945), .b(n_11055), .c(n_8944), .o(n_15708) );
in01f80 g557826 ( .a(n_15711), .o(n_11750) );
oa12f80 g557827 ( .a(n_11054), .b(n_11053), .c(n_12313), .o(n_15711) );
in01f80 g557828 ( .a(n_14802), .o(n_11749) );
oa12f80 g557829 ( .a(n_6657), .b(n_11052), .c(n_6659), .o(n_14802) );
in01f80 g557830 ( .a(n_12423), .o(n_12424) );
ao12f80 g557831 ( .a(n_10577), .b(n_10479), .c(x_in_17_13), .o(n_12423) );
in01f80 g557832 ( .a(n_11747), .o(n_11748) );
oa12f80 g557833 ( .a(n_9715), .b(n_9655), .c(x_in_17_10), .o(n_11747) );
in01f80 g557834 ( .a(n_11745), .o(n_11746) );
oa12f80 g557835 ( .a(n_9711), .b(n_9652), .c(x_in_17_8), .o(n_11745) );
in01f80 g557836 ( .a(n_11050), .o(n_11051) );
oa22f80 g557837 ( .a(n_8689), .b(n_9588), .c(n_9587), .d(n_11378), .o(n_11050) );
in01f80 g557838 ( .a(n_11743), .o(n_11744) );
oa12f80 g557839 ( .a(n_9710), .b(n_9649), .c(x_in_17_6), .o(n_11743) );
oa12f80 g557840 ( .a(n_9712), .b(n_9656), .c(x_in_17_11), .o(n_13975) );
oa22f80 g557841 ( .a(n_9363), .b(n_5806), .c(n_7211), .d(n_7212), .o(n_9364) );
ao22s80 g557842 ( .a(n_10153), .b(n_6037), .c(n_10152), .d(n_10151), .o(n_14470) );
ao12f80 g557843 ( .a(n_10040), .b(n_10039), .c(n_13246), .o(n_11049) );
in01f80 g557844 ( .a(n_15377), .o(n_12928) );
oa12f80 g557845 ( .a(n_11567), .b(n_11566), .c(n_11565), .o(n_15377) );
in01f80 g557846 ( .a(n_12421), .o(n_12422) );
ao12f80 g557847 ( .a(n_10748), .b(n_10747), .c(n_10746), .o(n_12421) );
oa12f80 g557848 ( .a(n_10019), .b(n_10018), .c(n_10017), .o(n_12810) );
in01f80 g557849 ( .a(n_12221), .o(n_11048) );
no03m80 g557850 ( .a(n_10150), .b(n_14855), .c(n_6594), .o(n_12221) );
ao12f80 g557851 ( .a(n_9843), .b(n_11047), .c(FE_OFN1244_n_12940), .o(n_14059) );
ao12f80 g557852 ( .a(n_10904), .b(n_10903), .c(n_10902), .o(n_13213) );
in01f80 g557853 ( .a(n_11741), .o(n_11742) );
ao12f80 g557854 ( .a(n_9865), .b(n_9864), .c(n_9863), .o(n_11741) );
oa12f80 g557855 ( .a(n_10767), .b(n_10766), .c(n_10765), .o(n_13211) );
in01f80 g557856 ( .a(n_12419), .o(n_12420) );
ao12f80 g557857 ( .a(n_10533), .b(n_10542), .c(n_10541), .o(n_12419) );
ao12f80 g557858 ( .a(n_9912), .b(n_9911), .c(n_9910), .o(n_12752) );
in01f80 g557859 ( .a(n_11739), .o(n_11740) );
oa22f80 g557860 ( .a(n_9056), .b(n_11863), .c(n_10429), .d(n_10430), .o(n_11739) );
in01f80 g557861 ( .a(n_11737), .o(n_11738) );
oa12f80 g557862 ( .a(n_10058), .b(n_10057), .c(n_10056), .o(n_11737) );
ao12f80 g557863 ( .a(n_9782), .b(n_10553), .c(n_5961), .o(n_11046) );
in01f80 g557864 ( .a(n_12417), .o(n_12418) );
ao22s80 g557865 ( .a(n_9511), .b(n_12025), .c(n_10536), .d(n_10535), .o(n_12417) );
in01f80 g557866 ( .a(n_11044), .o(n_11045) );
ao12f80 g557867 ( .a(n_9358), .b(n_10130), .c(n_9357), .o(n_11044) );
oa22f80 g557868 ( .a(n_9026), .b(n_12042), .c(n_10417), .d(n_10418), .o(n_14211) );
in01f80 g557869 ( .a(n_11735), .o(n_11736) );
oa12f80 g557870 ( .a(n_9776), .b(n_9583), .c(n_11273), .o(n_11735) );
ao12f80 g557871 ( .a(n_9909), .b(n_9908), .c(n_9907), .o(n_13382) );
in01f80 g557872 ( .a(n_15689), .o(n_12416) );
oa12f80 g557873 ( .a(n_10958), .b(n_10957), .c(n_10956), .o(n_15689) );
oa12f80 g557874 ( .a(n_11602), .b(n_11657), .c(n_12288), .o(n_13759) );
in01f80 g557875 ( .a(n_11733), .o(n_11734) );
oa12f80 g557876 ( .a(n_9775), .b(n_9580), .c(n_11282), .o(n_11733) );
ao22s80 g557877 ( .a(n_11055), .b(n_8847), .c(n_9441), .d(x_in_38_1), .o(n_13252) );
in01f80 g557878 ( .a(n_11731), .o(n_11732) );
oa12f80 g557879 ( .a(n_9780), .b(n_9685), .c(n_11163), .o(n_11731) );
ao12f80 g557880 ( .a(n_10908), .b(n_10907), .c(n_13251), .o(n_11730) );
ao22s80 g557881 ( .a(n_9508), .b(n_12022), .c(n_10397), .d(n_10398), .o(n_14213) );
in01f80 g557882 ( .a(n_12414), .o(n_12415) );
ao12f80 g557883 ( .a(n_10534), .b(n_10504), .c(FE_OFN656_n_10503), .o(n_12414) );
in01f80 g557884 ( .a(n_12412), .o(n_12413) );
ao12f80 g557885 ( .a(n_10762), .b(n_11153), .c(n_10761), .o(n_12412) );
oa12f80 g557886 ( .a(n_10148), .b(n_13943), .c(n_10149), .o(n_12807) );
in01f80 g557887 ( .a(n_11042), .o(n_11043) );
no03m80 g557888 ( .a(n_10149), .b(n_13943), .c(n_10148), .o(n_11042) );
in01f80 g557889 ( .a(n_11728), .o(n_11729) );
oa12f80 g557890 ( .a(n_10044), .b(n_10043), .c(n_10042), .o(n_11728) );
in01f80 g557891 ( .a(n_12410), .o(n_12411) );
ao12f80 g557892 ( .a(n_10545), .b(n_10401), .c(n_10400), .o(n_12410) );
ao22s80 g557893 ( .a(n_8850), .b(x_in_23_10), .c(n_10159), .d(n_11041), .o(n_12812) );
oa12f80 g557894 ( .a(n_10000), .b(n_9999), .c(n_9998), .o(n_12715) );
ao12f80 g557895 ( .a(n_10399), .b(n_10391), .c(n_10390), .o(n_13141) );
in01f80 g557896 ( .a(n_12408), .o(n_12409) );
ao12f80 g557897 ( .a(n_10439), .b(n_10436), .c(n_10435), .o(n_12408) );
oa22f80 g557898 ( .a(n_8586), .b(n_10147), .c(n_10146), .d(n_10145), .o(n_12233) );
ao22s80 g557899 ( .a(n_9361), .b(n_4047), .c(n_8141), .d(n_4046), .o(n_9362) );
in01f80 g557900 ( .a(n_11726), .o(n_11727) );
oa12f80 g557901 ( .a(n_9890), .b(n_9889), .c(n_9888), .o(n_11726) );
in01f80 g557902 ( .a(n_12406), .o(n_12407) );
ao22s80 g557903 ( .a(n_9516), .b(n_11968), .c(n_10551), .d(n_10550), .o(n_12406) );
in01f80 g557904 ( .a(n_12404), .o(n_12405) );
ao22s80 g557905 ( .a(n_9453), .b(n_12004), .c(n_10527), .d(n_10526), .o(n_12404) );
oa22f80 g557906 ( .a(n_8549), .b(n_10144), .c(n_10143), .d(n_10142), .o(n_12231) );
in01f80 g557907 ( .a(n_12402), .o(n_12403) );
ao12f80 g557908 ( .a(n_10523), .b(n_10521), .c(FE_OFN1256_n_10520), .o(n_12402) );
in01f80 g557909 ( .a(n_12400), .o(n_12401) );
ao12f80 g557910 ( .a(n_10519), .b(n_10540), .c(n_10539), .o(n_12400) );
ao22s80 g557911 ( .a(n_8930), .b(x_in_55_10), .c(n_10158), .d(n_11040), .o(n_12805) );
oa12f80 g557912 ( .a(n_10865), .b(n_10968), .c(n_10864), .o(n_13283) );
oa22f80 g557913 ( .a(n_8587), .b(n_10141), .c(n_10140), .d(n_10139), .o(n_12235) );
oa12f80 g557914 ( .a(n_10871), .b(n_10870), .c(n_10869), .o(n_13208) );
oa12f80 g557915 ( .a(n_9675), .b(n_10538), .c(n_10537), .o(n_14357) );
ao12f80 g557916 ( .a(n_10896), .b(n_10895), .c(n_10894), .o(n_13104) );
in01f80 g557917 ( .a(n_11724), .o(n_11725) );
oa22f80 g557918 ( .a(n_9065), .b(n_11976), .c(n_10554), .d(n_10555), .o(n_11724) );
oa12f80 g557919 ( .a(n_10756), .b(n_10755), .c(n_10754), .o(n_13206) );
in01f80 g557920 ( .a(n_11038), .o(n_11039) );
ao12f80 g557921 ( .a(n_9349), .b(n_9363), .c(n_9348), .o(n_11038) );
in01f80 g557922 ( .a(n_12398), .o(n_12399) );
ao12f80 g557923 ( .a(n_10512), .b(n_10556), .c(n_10557), .o(n_12398) );
ao22s80 g557924 ( .a(n_8923), .b(x_in_15_10), .c(n_10157), .d(n_11037), .o(n_12801) );
oa12f80 g557925 ( .a(n_10047), .b(n_10046), .c(n_10045), .o(n_12799) );
oa22f80 g557926 ( .a(n_8592), .b(n_10138), .c(FE_OFN574_n_10137), .d(FE_OFN576_n_10136), .o(n_12229) );
in01f80 g557927 ( .a(n_11722), .o(n_11723) );
oa12f80 g557928 ( .a(n_9664), .b(n_9663), .c(n_9662), .o(n_11722) );
oa12f80 g557929 ( .a(n_10015), .b(n_10014), .c(n_10013), .o(n_12797) );
oa22f80 g557930 ( .a(n_8993), .b(n_11979), .c(n_10514), .d(n_10513), .o(n_14422) );
in01f80 g557931 ( .a(n_11720), .o(n_11721) );
na03f80 g557932 ( .a(n_9061), .b(n_11036), .c(n_6599), .o(n_11720) );
oa12f80 g557933 ( .a(n_6598), .b(n_11035), .c(n_9062), .o(n_12793) );
oa12f80 g557934 ( .a(n_10038), .b(n_10037), .c(n_10036), .o(n_12795) );
ao22s80 g557935 ( .a(n_9501), .b(n_11961), .c(n_10505), .d(FE_OFN869_n_10506), .o(n_14400) );
in01f80 g557936 ( .a(n_11718), .o(n_11719) );
ao12f80 g557937 ( .a(n_10029), .b(n_10028), .c(n_10027), .o(n_11718) );
in01f80 g557938 ( .a(n_12396), .o(n_12397) );
ao22s80 g557939 ( .a(n_9498), .b(n_11958), .c(n_10502), .d(FE_OFN865_n_10501), .o(n_12396) );
ao22s80 g557940 ( .a(n_9495), .b(n_11955), .c(n_10498), .d(FE_OFN1240_n_10499), .o(n_14392) );
in01f80 g557941 ( .a(n_11716), .o(n_11717) );
oa12f80 g557942 ( .a(n_10035), .b(n_10034), .c(n_10033), .o(n_11716) );
in01f80 g557943 ( .a(n_12394), .o(n_12395) );
ao12f80 g557944 ( .a(n_10500), .b(n_10496), .c(FE_OFN863_n_10495), .o(n_12394) );
in01f80 g557945 ( .a(n_12392), .o(n_12393) );
oa12f80 g557946 ( .a(n_10497), .b(n_10493), .c(FE_OFN861_n_10492), .o(n_12392) );
in01f80 g557947 ( .a(n_12390), .o(n_12391) );
ao12f80 g557948 ( .a(n_10494), .b(n_10490), .c(FE_OFN1238_n_10491), .o(n_12390) );
oa12f80 g557949 ( .a(n_9885), .b(n_9884), .c(n_9883), .o(n_13386) );
in01f80 g557950 ( .a(n_11714), .o(n_11715) );
oa12f80 g557951 ( .a(n_10026), .b(n_10025), .c(n_10024), .o(n_11714) );
in01f80 g557952 ( .a(n_11712), .o(n_11713) );
oa12f80 g557953 ( .a(n_10032), .b(n_10031), .c(n_10030), .o(n_11712) );
in01f80 g557954 ( .a(n_12388), .o(n_12389) );
ao22s80 g557955 ( .a(n_9489), .b(n_11964), .c(n_10508), .d(n_10507), .o(n_12388) );
ao22s80 g557956 ( .a(n_8922), .b(x_in_47_10), .c(n_10156), .d(n_11034), .o(n_12788) );
oa12f80 g557957 ( .a(n_10078), .b(n_10077), .c(n_10076), .o(n_14951) );
oa22f80 g557958 ( .a(n_8591), .b(n_10135), .c(n_10134), .d(n_10133), .o(n_12227) );
in01f80 g557959 ( .a(n_12386), .o(n_12387) );
ao22s80 g557960 ( .a(n_9519), .b(n_12001), .c(n_10546), .d(n_10547), .o(n_12386) );
oa12f80 g557961 ( .a(n_9951), .b(n_9950), .c(n_9949), .o(n_12786) );
ao12f80 g557962 ( .a(n_9870), .b(n_9869), .c(n_9868), .o(n_13353) );
oa12f80 g557963 ( .a(n_9928), .b(n_9927), .c(n_9926), .o(n_12784) );
oa12f80 g557964 ( .a(n_9925), .b(n_9924), .c(n_9923), .o(n_12782) );
in01f80 g557965 ( .a(n_15121), .o(n_12385) );
oa12f80 g557966 ( .a(n_10946), .b(n_10945), .c(n_10944), .o(n_15121) );
oa12f80 g557967 ( .a(n_9986), .b(n_9985), .c(n_9984), .o(n_12780) );
ao12f80 g557968 ( .a(n_9942), .b(n_9941), .c(n_9940), .o(n_12778) );
in01f80 g557969 ( .a(n_12926), .o(n_12927) );
oa12f80 g557970 ( .a(n_11529), .b(n_11528), .c(x_in_53_13), .o(n_12926) );
oa12f80 g557971 ( .a(n_9960), .b(n_9959), .c(n_9958), .o(n_12776) );
in01f80 g557972 ( .a(n_11710), .o(n_11711) );
ao22s80 g557973 ( .a(n_9110), .b(n_11252), .c(n_9653), .d(n_9654), .o(n_11710) );
ao12f80 g557974 ( .a(n_9948), .b(n_9947), .c(n_9946), .o(n_12774) );
in01f80 g557975 ( .a(n_11708), .o(n_11709) );
ao22s80 g557976 ( .a(n_9115), .b(n_11330), .c(n_9650), .d(n_9651), .o(n_11708) );
oa12f80 g557977 ( .a(n_9898), .b(n_9897), .c(n_9896), .o(n_12772) );
oa12f80 g557978 ( .a(n_9971), .b(n_9970), .c(n_9969), .o(n_12770) );
oa12f80 g557979 ( .a(n_9963), .b(n_9962), .c(n_9961), .o(n_12768) );
oa12f80 g557980 ( .a(n_10753), .b(n_10752), .c(n_10751), .o(n_13175) );
in01f80 g557981 ( .a(n_11706), .o(n_11707) );
oa12f80 g557982 ( .a(n_9768), .b(n_9657), .c(x_in_17_12), .o(n_11706) );
in01f80 g557983 ( .a(n_11704), .o(n_11705) );
ao12f80 g557984 ( .a(n_9857), .b(n_9856), .c(n_9855), .o(n_11704) );
ao12f80 g557985 ( .a(n_12283), .b(n_12282), .c(n_12281), .o(n_14116) );
oa22f80 g557986 ( .a(n_9483), .b(n_11930), .c(n_10474), .d(n_4603), .o(n_14354) );
in01f80 g557987 ( .a(n_15694), .o(n_11703) );
oa12f80 g557988 ( .a(n_9966), .b(n_9965), .c(n_9964), .o(n_15694) );
in01f80 g557989 ( .a(n_11701), .o(n_11702) );
oa12f80 g557990 ( .a(n_9893), .b(n_9892), .c(n_9891), .o(n_11701) );
in01f80 g557991 ( .a(n_12383), .o(n_12384) );
oa22f80 g557992 ( .a(n_9481), .b(n_11915), .c(n_10461), .d(n_11700), .o(n_12383) );
ao22s80 g557993 ( .a(n_9479), .b(n_11927), .c(n_10471), .d(n_10472), .o(n_14348) );
in01f80 g557994 ( .a(n_12381), .o(n_12382) );
ao12f80 g557995 ( .a(n_10473), .b(n_10468), .c(FE_OFN1214_n_10469), .o(n_12381) );
in01f80 g557996 ( .a(n_12379), .o(n_12380) );
oa12f80 g557997 ( .a(n_10470), .b(n_10466), .c(FE_OFN1212_n_10465), .o(n_12379) );
in01f80 g557998 ( .a(n_12377), .o(n_12378) );
ao12f80 g557999 ( .a(n_10467), .b(n_10463), .c(FE_OFN704_n_10462), .o(n_12377) );
in01f80 g558000 ( .a(n_12375), .o(n_12376) );
oa12f80 g558001 ( .a(n_10464), .b(n_10459), .c(FE_OFN1210_n_10458), .o(n_12375) );
in01f80 g558002 ( .a(n_12924), .o(n_12925) );
ao12f80 g558003 ( .a(n_10460), .b(n_10457), .c(FE_OFN1208_n_10456), .o(n_12924) );
ao12f80 g558004 ( .a(n_6591), .b(n_11699), .c(n_9041), .o(n_14538) );
in01f80 g558005 ( .a(n_12374), .o(n_13170) );
na02f80 g558006 ( .a(n_9854), .b(n_11699), .o(n_12374) );
in01f80 g558007 ( .a(n_12922), .o(n_12923) );
ao12f80 g558008 ( .a(n_10451), .b(n_10447), .c(n_9038), .o(n_12922) );
in01f80 g558009 ( .a(n_12920), .o(n_12921) );
ao22s80 g558010 ( .a(n_9486), .b(n_12373), .c(n_10476), .d(n_10475), .o(n_12920) );
ao22s80 g558011 ( .a(n_8912), .b(x_in_31_10), .c(n_10155), .d(n_11698), .o(n_12762) );
ao12f80 g558012 ( .a(n_11431), .b(n_11430), .c(n_11429), .o(n_24439) );
oa22f80 g558013 ( .a(n_8585), .b(n_11033), .c(n_11032), .d(n_11031), .o(n_12225) );
in01f80 g558014 ( .a(n_12918), .o(n_12919) );
oa12f80 g558015 ( .a(n_10448), .b(n_10446), .c(n_9034), .o(n_12918) );
oa12f80 g558016 ( .a(n_9906), .b(n_9905), .c(x_in_53_3), .o(n_12821) );
ao12f80 g558017 ( .a(n_9939), .b(n_9938), .c(n_9937), .o(n_13380) );
oa12f80 g558018 ( .a(n_10884), .b(n_10883), .c(n_10882), .o(n_13169) );
ao12f80 g558019 ( .a(n_10006), .b(n_10005), .c(n_10004), .o(n_12766) );
ao22s80 g558020 ( .a(n_9475), .b(n_12372), .c(n_10354), .d(n_10355), .o(n_14336) );
in01f80 g558021 ( .a(n_12916), .o(n_12917) );
ao22s80 g558022 ( .a(n_9472), .b(n_12371), .c(n_10443), .d(n_10442), .o(n_12916) );
oa12f80 g558023 ( .a(n_10049), .b(n_11697), .c(n_10048), .o(n_13798) );
ao22s80 g558024 ( .a(n_9525), .b(n_12370), .c(n_10369), .d(n_10370), .o(n_14334) );
in01f80 g558025 ( .a(n_12914), .o(n_12915) );
ao12f80 g558026 ( .a(n_10441), .b(n_10368), .c(n_10367), .o(n_12914) );
in01f80 g558027 ( .a(n_12912), .o(n_12913) );
oa12f80 g558028 ( .a(n_10440), .b(n_10438), .c(n_10437), .o(n_12912) );
ao12f80 g558029 ( .a(n_10051), .b(n_11697), .c(n_10050), .o(n_25530) );
oa12f80 g558030 ( .a(n_10868), .b(n_10867), .c(n_10866), .o(n_13261) );
ao12f80 g558031 ( .a(n_10832), .b(n_10831), .c(x_in_19_12), .o(n_13229) );
in01f80 g558032 ( .a(n_12910), .o(n_12911) );
ao22s80 g558033 ( .a(n_9492), .b(FE_OFN1101_n_12369), .c(n_10445), .d(n_10444), .o(n_12910) );
ao22s80 g558034 ( .a(n_8852), .b(x_in_63_10), .c(n_10154), .d(n_11696), .o(n_12755) );
oa22f80 g558035 ( .a(n_8590), .b(n_11030), .c(n_11029), .d(n_11028), .o(n_12223) );
ao22s80 g558036 ( .a(n_9463), .b(n_12368), .c(n_10543), .d(n_10544), .o(n_14430) );
in01f80 g558037 ( .a(FE_OFN1194_n_12908), .o(n_12909) );
oa22f80 g558038 ( .a(n_9469), .b(n_12367), .c(n_10478), .d(n_12366), .o(n_12908) );
oa12f80 g558039 ( .a(n_9356), .b(n_9355), .c(n_9354), .o(n_14574) );
in01f80 g558040 ( .a(n_12906), .o(n_12907) );
ao12f80 g558041 ( .a(n_10428), .b(n_10432), .c(n_10431), .o(n_12906) );
in01f80 g558042 ( .a(n_12904), .o(n_12905) );
ao12f80 g558043 ( .a(n_10764), .b(n_10763), .c(n_12365), .o(n_12904) );
oa12f80 g558044 ( .a(n_10923), .b(n_10922), .c(x_in_1_7), .o(n_13313) );
ao22s80 g558045 ( .a(n_9565), .b(n_10167), .c(n_8635), .d(n_9564), .o(n_12364) );
ao22s80 g558046 ( .a(n_10349), .b(n_10168), .c(n_10348), .d(n_8654), .o(n_12903) );
ao12f80 g558047 ( .a(n_10731), .b(n_10730), .c(n_10729), .o(n_13965) );
in01f80 g558048 ( .a(n_15696), .o(n_13499) );
oa12f80 g558049 ( .a(n_11605), .b(n_11604), .c(n_11603), .o(n_15696) );
in01f80 g558050 ( .a(n_12901), .o(n_12902) );
oa12f80 g558051 ( .a(n_10453), .b(n_10449), .c(n_9042), .o(n_12901) );
oa12f80 g558052 ( .a(n_9974), .b(n_9973), .c(n_9972), .o(n_12727) );
ao12f80 g558053 ( .a(n_10863), .b(n_10862), .c(n_10861), .o(n_13106) );
in01f80 g558054 ( .a(n_11027), .o(n_12854) );
oa12f80 g558055 ( .a(n_8808), .b(n_8809), .c(n_8807), .o(n_11027) );
in01f80 g558056 ( .a(n_12362), .o(n_12363) );
ao12f80 g558057 ( .a(n_11695), .b(n_9847), .c(n_9846), .o(n_12362) );
in01f80 g558058 ( .a(n_12899), .o(n_12900) );
oa12f80 g558059 ( .a(n_12361), .b(n_10726), .c(n_10725), .o(n_12899) );
oa12f80 g558060 ( .a(n_11694), .b(n_9849), .c(n_9848), .o(n_12750) );
in01f80 g558061 ( .a(n_12359), .o(n_12360) );
oa12f80 g558062 ( .a(n_12749), .b(n_9859), .c(n_9858), .o(n_12359) );
in01f80 g558063 ( .a(n_12357), .o(n_12358) );
ao12f80 g558064 ( .a(n_11693), .b(n_9804), .c(n_9803), .o(n_12357) );
ao12f80 g558065 ( .a(n_11692), .b(n_9845), .c(n_9844), .o(n_12833) );
ao12f80 g558066 ( .a(n_10891), .b(n_10890), .c(n_10889), .o(n_13223) );
oa12f80 g558067 ( .a(n_9880), .b(n_9879), .c(n_9878), .o(n_13379) );
in01f80 g558068 ( .a(n_12897), .o(n_12898) );
oa12f80 g558069 ( .a(n_12356), .b(n_10722), .c(n_10721), .o(n_12897) );
in01f80 g558070 ( .a(n_12354), .o(n_12355) );
oa12f80 g558071 ( .a(n_9842), .b(n_9841), .c(n_9840), .o(n_12354) );
in01f80 g558072 ( .a(n_15698), .o(n_14590) );
oa12f80 g558073 ( .a(n_12864), .b(n_12863), .c(n_12862), .o(n_15698) );
oa12f80 g558074 ( .a(n_10090), .b(n_10089), .c(n_10088), .o(n_14926) );
in01f80 g558075 ( .a(n_12352), .o(n_12353) );
oa12f80 g558076 ( .a(n_9839), .b(n_9838), .c(n_9837), .o(n_12352) );
oa12f80 g558077 ( .a(n_10985), .b(n_10984), .c(n_10983), .o(n_13233) );
oa12f80 g558078 ( .a(n_11527), .b(n_11526), .c(x_in_51_11), .o(n_13631) );
oa12f80 g558079 ( .a(n_9920), .b(n_9919), .c(x_in_51_10), .o(n_12837) );
oa12f80 g558080 ( .a(n_9902), .b(n_9901), .c(x_in_51_9), .o(n_12746) );
in01f80 g558081 ( .a(n_15358), .o(n_13730) );
oa12f80 g558082 ( .a(n_10624), .b(n_10623), .c(n_10622), .o(n_15358) );
ao12f80 g558083 ( .a(n_9918), .b(n_9917), .c(x_in_51_8), .o(n_12744) );
ao22s80 g558084 ( .a(n_9504), .b(n_12351), .c(n_10524), .d(n_10525), .o(n_14434) );
oa12f80 g558085 ( .a(n_9900), .b(n_9899), .c(x_in_51_7), .o(n_12742) );
ao12f80 g558086 ( .a(n_10822), .b(n_10821), .c(n_10820), .o(n_13309) );
ao12f80 g558087 ( .a(n_9916), .b(n_9915), .c(x_in_51_6), .o(n_12740) );
ao12f80 g558088 ( .a(n_9914), .b(n_9913), .c(x_in_51_5), .o(n_12738) );
ao12f80 g558089 ( .a(n_9895), .b(n_9894), .c(x_in_51_4), .o(n_12736) );
ao22s80 g558090 ( .a(n_11052), .b(n_8438), .c(n_9393), .d(x_in_28_1), .o(n_13247) );
ao22s80 g558091 ( .a(n_9366), .b(n_3718), .c(n_8150), .d(n_3717), .o(n_10132) );
ao12f80 g558092 ( .a(n_9836), .b(n_9835), .c(n_9834), .o(n_12734) );
ao12f80 g558093 ( .a(n_10716), .b(n_10715), .c(n_10714), .o(n_13145) );
oa12f80 g558094 ( .a(n_10819), .b(n_10818), .c(n_10817), .o(n_13307) );
in01f80 g558095 ( .a(n_13760), .o(n_13498) );
oa12f80 g558096 ( .a(n_11629), .b(n_11628), .c(n_11627), .o(n_13760) );
oa12f80 g558097 ( .a(n_11558), .b(n_12237), .c(n_11557), .o(n_13732) );
in01f80 g558098 ( .a(n_13830), .o(n_12896) );
ao12f80 g558099 ( .a(n_10919), .b(n_12313), .c(n_11579), .o(n_13830) );
oa12f80 g558100 ( .a(n_10415), .b(n_10411), .c(FE_OFN843_n_10412), .o(n_14310) );
oa12f80 g558101 ( .a(n_10874), .b(n_10873), .c(n_10872), .o(n_13244) );
in01f80 g558102 ( .a(n_12894), .o(n_12895) );
ao12f80 g558103 ( .a(n_10410), .b(n_10407), .c(n_10406), .o(n_12894) );
oa12f80 g558104 ( .a(n_10408), .b(n_10404), .c(n_10405), .o(n_14308) );
in01f80 g558105 ( .a(n_12349), .o(n_12350) );
na03f80 g558106 ( .a(n_11691), .b(n_13874), .c(n_11690), .o(n_12349) );
in01f80 g558107 ( .a(n_13675), .o(n_13497) );
oa12f80 g558108 ( .a(n_11596), .b(n_11595), .c(n_11594), .o(n_13675) );
in01f80 g558109 ( .a(n_12892), .o(n_12893) );
oa12f80 g558110 ( .a(n_10706), .b(n_11071), .c(n_10705), .o(n_12892) );
in01f80 g558111 ( .a(n_12347), .o(n_12348) );
oa12f80 g558112 ( .a(n_9680), .b(n_10549), .c(n_10548), .o(n_12347) );
ao12f80 g558113 ( .a(n_10704), .b(n_10703), .c(n_10702), .o(n_13140) );
in01f80 g558114 ( .a(n_12345), .o(n_12346) );
oa12f80 g558115 ( .a(n_9605), .b(n_9606), .c(n_6760), .o(n_12345) );
in01f80 g558116 ( .a(n_11688), .o(n_11689) );
oa12f80 g558117 ( .a(n_9347), .b(n_9708), .c(x_in_41_14), .o(n_11688) );
in01f80 g558118 ( .a(n_12890), .o(n_12891) );
ao22s80 g558119 ( .a(n_9460), .b(n_12344), .c(n_10350), .d(n_10351), .o(n_12890) );
in01f80 g558120 ( .a(n_12888), .o(n_12889) );
ao12f80 g558121 ( .a(n_10394), .b(n_10414), .c(n_10413), .o(n_12888) );
oa12f80 g558122 ( .a(n_10947), .b(n_12343), .c(n_12342), .o(n_22420) );
in01f80 g558123 ( .a(n_15124), .o(n_12341) );
ao12f80 g558124 ( .a(n_10123), .b(n_10122), .c(n_10121), .o(n_15124) );
in01f80 g558125 ( .a(n_12886), .o(n_12887) );
oa12f80 g558126 ( .a(n_10522), .b(n_10425), .c(FE_OFN658_n_10424), .o(n_12886) );
ao12f80 g558127 ( .a(n_11125), .b(n_11687), .c(n_9813), .o(n_17164) );
na02f80 g558128 ( .a(n_12340), .b(n_10686), .o(n_20335) );
in01f80 g558129 ( .a(n_12338), .o(n_12339) );
oa12f80 g558130 ( .a(n_9955), .b(n_9954), .c(x_in_25_3), .o(n_12338) );
ao12f80 g558131 ( .a(n_10681), .b(n_10680), .c(n_10679), .o(n_13133) );
in01f80 g558132 ( .a(n_12884), .o(n_12885) );
oa22f80 g558133 ( .a(n_9410), .b(n_12635), .c(n_9411), .d(x_in_33_12), .o(n_12884) );
oa12f80 g558134 ( .a(n_10055), .b(n_10054), .c(n_10053), .o(n_12730) );
oa12f80 g558135 ( .a(n_10022), .b(n_10021), .c(n_10020), .o(n_12725) );
in01f80 g558136 ( .a(n_12882), .o(n_12883) );
ao12f80 g558137 ( .a(n_10899), .b(n_10898), .c(n_10897), .o(n_12882) );
oa12f80 g558138 ( .a(n_10012), .b(n_10011), .c(n_10010), .o(n_12723) );
in01f80 g558139 ( .a(n_12336), .o(n_12337) );
ao12f80 g558140 ( .a(n_10009), .b(n_10008), .c(n_10007), .o(n_12336) );
ao12f80 g558141 ( .a(n_10087), .b(n_10086), .c(n_10085), .o(n_24195) );
oa12f80 g558142 ( .a(n_10003), .b(n_10002), .c(n_10001), .o(n_12721) );
in01f80 g558143 ( .a(n_12334), .o(n_12335) );
oa12f80 g558144 ( .a(n_9991), .b(n_9990), .c(n_9989), .o(n_12334) );
in01f80 g558145 ( .a(n_12332), .o(n_12333) );
ao12f80 g558146 ( .a(n_9994), .b(n_9993), .c(n_9992), .o(n_12332) );
in01f80 g558147 ( .a(n_15428), .o(n_13496) );
oa12f80 g558148 ( .a(n_11570), .b(n_11569), .c(n_11568), .o(n_15428) );
in01f80 g558149 ( .a(n_12880), .o(n_12881) );
oa12f80 g558150 ( .a(n_10836), .b(n_10835), .c(x_in_25_13), .o(n_12880) );
in01f80 g558151 ( .a(n_12330), .o(n_12331) );
ao12f80 g558152 ( .a(n_9695), .b(n_9593), .c(n_9592), .o(n_12330) );
ao12f80 g558153 ( .a(n_6593), .b(n_11684), .c(n_9006), .o(n_14529) );
in01f80 g558154 ( .a(n_11685), .o(n_11686) );
ao12f80 g558155 ( .a(n_9353), .b(n_10126), .c(n_9352), .o(n_11685) );
in01f80 g558156 ( .a(n_12329), .o(n_13115) );
na02f80 g558157 ( .a(n_9862), .b(n_11684), .o(n_12329) );
in01f80 g558158 ( .a(n_15100), .o(n_12879) );
ao12f80 g558159 ( .a(n_10988), .b(n_10987), .c(n_10986), .o(n_15100) );
ao12f80 g558160 ( .a(n_11451), .b(n_11450), .c(n_11449), .o(n_13686) );
ao12f80 g558161 ( .a(n_11459), .b(FE_OFN815_n_12310), .c(n_11458), .o(n_12878) );
ao12f80 g558162 ( .a(n_9979), .b(n_9978), .c(n_9977), .o(n_13384) );
oa12f80 g558163 ( .a(n_10795), .b(n_10794), .c(n_10793), .o(n_13289) );
ao12f80 g558164 ( .a(n_9877), .b(n_9876), .c(n_9875), .o(n_13381) );
oa22f80 g558165 ( .a(n_10130), .b(n_5815), .c(n_6583), .d(n_6584), .o(n_10131) );
in01f80 g558166 ( .a(n_12327), .o(n_12328) );
ao12f80 g558167 ( .a(n_9997), .b(n_9996), .c(n_9995), .o(n_12327) );
in01f80 g558168 ( .a(n_12876), .o(n_12877) );
oa12f80 g558169 ( .a(n_10881), .b(n_10880), .c(n_10879), .o(n_12876) );
in01f80 g558170 ( .a(n_14081), .o(n_12875) );
ao12f80 g558171 ( .a(n_10939), .b(n_10938), .c(n_10937), .o(n_14081) );
in01f80 g558172 ( .a(n_12325), .o(n_12326) );
ao22s80 g558173 ( .a(n_9003), .b(n_11683), .c(n_9590), .d(n_9591), .o(n_12325) );
no02f80 g558174 ( .a(n_10650), .b(n_6595), .o(n_14526) );
in01f80 g558175 ( .a(n_12873), .o(n_12874) );
oa12f80 g558176 ( .a(n_10792), .b(n_10791), .c(n_10790), .o(n_12873) );
in01f80 g558177 ( .a(n_12323), .o(n_12324) );
oa12f80 g558178 ( .a(n_9745), .b(n_9689), .c(n_11682), .o(n_12323) );
ao12f80 g558179 ( .a(n_11611), .b(n_11610), .c(n_11609), .o(n_13688) );
ao12f80 g558180 ( .a(n_9945), .b(n_9944), .c(n_9943), .o(n_13383) );
in01f80 g558181 ( .a(n_11680), .o(n_11681) );
ao12f80 g558182 ( .a(n_9351), .b(n_10128), .c(n_9350), .o(n_11680) );
in01f80 g558183 ( .a(n_12321), .o(n_12322) );
oa22f80 g558184 ( .a(n_9081), .b(n_11982), .c(n_10515), .d(n_10516), .o(n_12321) );
oa22f80 g558185 ( .a(n_10128), .b(n_5809), .c(n_6507), .d(n_6508), .o(n_10129) );
in01f80 g558186 ( .a(n_13494), .o(n_13495) );
oa12f80 g558187 ( .a(n_11442), .b(n_11441), .c(n_11440), .o(n_13494) );
oa12f80 g558188 ( .a(n_10668), .b(n_10667), .c(n_10666), .o(n_13886) );
in01f80 g558189 ( .a(n_15421), .o(n_13493) );
oa12f80 g558190 ( .a(n_11550), .b(n_11549), .c(n_11548), .o(n_15421) );
ao12f80 g558191 ( .a(n_11523), .b(n_11522), .c(n_11521), .o(n_12872) );
oa12f80 g558192 ( .a(n_10972), .b(n_10971), .c(n_10970), .o(n_13227) );
in01f80 g558193 ( .a(n_12319), .o(n_12320) );
ao22s80 g558194 ( .a(n_8990), .b(FE_OFN1204_n_11679), .c(n_9597), .d(n_9598), .o(n_12319) );
ao12f80 g558195 ( .a(n_11690), .b(n_13874), .c(n_11691), .o(n_13107) );
ao22s80 g558196 ( .a(n_9456), .b(n_12318), .c(n_10395), .d(n_10396), .o(n_14293) );
oa22f80 g558197 ( .a(n_10126), .b(n_5812), .c(n_6457), .d(n_6458), .o(n_10127) );
ao12f80 g558198 ( .a(n_10974), .b(n_11676), .c(n_10973), .o(n_12317) );
oa12f80 g558199 ( .a(n_10084), .b(n_10166), .c(n_10083), .o(n_12814) );
na02f80 g558200 ( .a(n_12316), .b(n_10691), .o(n_18092) );
in01f80 g558201 ( .a(n_13677), .o(n_13492) );
oa12f80 g558202 ( .a(n_11599), .b(n_11598), .c(n_11597), .o(n_13677) );
ao12f80 g558203 ( .a(n_6607), .b(n_11678), .c(n_8970), .o(n_14071) );
in01f80 g558204 ( .a(n_12315), .o(n_13101) );
na02f80 g558205 ( .a(n_9814), .b(n_11678), .o(n_12315) );
in01f80 g558206 ( .a(n_12870), .o(n_12871) );
ao12f80 g558207 ( .a(n_10617), .b(n_10616), .c(n_10615), .o(n_12870) );
oa12f80 g558208 ( .a(n_10649), .b(n_12314), .c(FE_OFN642_n_12432), .o(n_15235) );
oa12f80 g558209 ( .a(n_9931), .b(n_9930), .c(n_9929), .o(n_13385) );
ao22s80 g558210 ( .a(n_12313), .b(n_12312), .c(n_11580), .d(x_in_8_1), .o(n_13249) );
oa22f80 g558211 ( .a(FE_OFN829_n_8424), .b(n_23291), .c(n_721), .d(FE_OFN1118_rst), .o(n_11026) );
oa22f80 g558212 ( .a(n_8423), .b(n_21988), .c(n_1730), .d(FE_OFN105_n_27449), .o(n_11025) );
oa22f80 g558213 ( .a(FE_OFN815_n_12310), .b(FE_OFN405_n_28303), .c(n_337), .d(n_29104), .o(n_12311) );
oa22f80 g558214 ( .a(n_8481), .b(FE_OFN406_n_28303), .c(n_905), .d(FE_OFN127_n_27449), .o(n_11024) );
oa22f80 g558215 ( .a(n_8422), .b(FE_OFN149_n_25677), .c(n_1828), .d(FE_OFN63_n_27012), .o(n_11023) );
oa22f80 g558216 ( .a(n_11676), .b(FE_OFN411_n_28303), .c(n_987), .d(FE_OFN335_n_4860), .o(n_11677) );
oa22f80 g558217 ( .a(n_11365), .b(FE_OFN265_n_4280), .c(n_1284), .d(FE_OFN1181_rst), .o(n_11675) );
oa22f80 g558218 ( .a(n_8006), .b(FE_OFN267_n_4280), .c(n_1318), .d(FE_OFN1110_rst), .o(n_10125) );
oa22f80 g558219 ( .a(n_8008), .b(FE_OFN260_n_4280), .c(n_1433), .d(FE_OFN127_n_27449), .o(n_10124) );
oa22f80 g558220 ( .a(n_8890), .b(n_29046), .c(n_439), .d(FE_OFN326_n_4860), .o(n_11674) );
oa22f80 g558221 ( .a(n_8447), .b(FE_OFN208_n_29661), .c(n_308), .d(FE_OFN326_n_4860), .o(n_11022) );
oa22f80 g558222 ( .a(FE_OFN538_n_10328), .b(n_23291), .c(n_1025), .d(FE_OFN63_n_27012), .o(n_12869) );
oa22f80 g558223 ( .a(n_9392), .b(FE_OFN303_n_3069), .c(n_1005), .d(FE_OFN63_n_27012), .o(n_12309) );
ao22s80 g558224 ( .a(n_11672), .b(n_4300), .c(x_out_59_25), .d(FE_OFN280_n_16656), .o(n_11673) );
ao22s80 g558225 ( .a(n_12867), .b(n_4350), .c(x_out_57_25), .d(FE_OFN279_n_16656), .o(n_12868) );
ao22s80 g558226 ( .a(n_11670), .b(n_2777), .c(x_out_58_25), .d(FE_OFN276_n_16893), .o(n_11671) );
ao22s80 g558227 ( .a(n_11668), .b(n_4298), .c(x_out_63_25), .d(FE_OFN271_n_16028), .o(n_11669) );
ao22s80 g558228 ( .a(n_11666), .b(n_2822), .c(x_out_60_25), .d(n_27400), .o(n_11667) );
ao22s80 g558229 ( .a(n_11664), .b(n_2824), .c(x_out_61_25), .d(n_16656), .o(n_11665) );
ao22s80 g558230 ( .a(n_11662), .b(n_4302), .c(x_out_62_25), .d(FE_OFN274_n_16893), .o(n_11663) );
in01f80 g558231 ( .a(n_12719), .o(n_14146) );
oa22f80 g558232 ( .a(n_8962), .b(n_7977), .c(n_8961), .d(n_8794), .o(n_12719) );
ao22s80 g558233 ( .a(n_9142), .b(x_in_43_11), .c(n_10016), .d(n_8443), .o(n_11661) );
oa22f80 g558234 ( .a(n_10023), .b(n_5754), .c(n_9144), .d(x_in_5_11), .o(n_12839) );
ao22s80 g558235 ( .a(n_9145), .b(x_in_27_10), .c(n_10041), .d(n_7417), .o(n_11660) );
ao22s80 g558236 ( .a(n_9170), .b(x_in_7_9), .c(n_10052), .d(n_7320), .o(n_11659) );
in01f80 g558237 ( .a(FE_OFN817_n_13135), .o(n_11658) );
oa22f80 g558238 ( .a(n_9365), .b(n_6324), .c(n_8604), .d(n_6323), .o(n_13135) );
ao12f80 g558239 ( .a(n_10709), .b(n_8860), .c(n_8861), .o(n_12308) );
in01f80 g558251 ( .a(n_17657), .o(n_12520) );
na02f80 g558252 ( .a(n_15285), .b(x_in_14_0), .o(n_17657) );
in01f80 g558253 ( .a(n_12306), .o(n_12307) );
no02f80 g558254 ( .a(n_11657), .b(x_in_38_2), .o(n_12306) );
in01f80 g558255 ( .a(n_17663), .o(n_12521) );
na02f80 g558256 ( .a(n_15340), .b(x_in_22_0), .o(n_17663) );
na02f80 g558257 ( .a(n_9505), .b(n_1511), .o(n_11656) );
na02f80 g558258 ( .a(n_11654), .b(n_11653), .o(n_11655) );
in01f80 g558259 ( .a(n_12519), .o(n_17654) );
no02f80 g558260 ( .a(n_11654), .b(n_11653), .o(n_12519) );
in01f80 g558261 ( .a(n_17660), .o(n_12517) );
na02f80 g558262 ( .a(n_15647), .b(x_in_54_0), .o(n_17660) );
na02f80 g558263 ( .a(n_11657), .b(x_in_38_2), .o(n_12950) );
na02f80 g558264 ( .a(n_11651), .b(n_11650), .o(n_11652) );
in01f80 g558265 ( .a(n_12515), .o(n_17642) );
no02f80 g558266 ( .a(n_11651), .b(n_11650), .o(n_12515) );
na02f80 g558267 ( .a(n_11648), .b(n_11647), .o(n_11649) );
in01f80 g558268 ( .a(n_12518), .o(n_17651) );
no02f80 g558269 ( .a(n_11648), .b(n_11647), .o(n_12518) );
na02f80 g558270 ( .a(n_11645), .b(n_11644), .o(n_11646) );
in01f80 g558271 ( .a(n_12516), .o(n_17648) );
no02f80 g558272 ( .a(n_11645), .b(n_11644), .o(n_12516) );
na02f80 g558273 ( .a(n_9513), .b(n_738), .o(n_11643) );
na02f80 g558274 ( .a(n_11641), .b(n_11640), .o(n_11642) );
in01f80 g558275 ( .a(n_12514), .o(n_17639) );
no02f80 g558276 ( .a(n_11641), .b(n_11640), .o(n_12514) );
in01f80 g558277 ( .a(n_12304), .o(n_12305) );
no02f80 g558278 ( .a(n_11639), .b(n_11638), .o(n_12304) );
na02f80 g558279 ( .a(n_11639), .b(n_11638), .o(n_12954) );
in01f80 g558280 ( .a(n_12302), .o(n_12303) );
no02f80 g558281 ( .a(n_11637), .b(n_11636), .o(n_12302) );
na02f80 g558282 ( .a(n_11637), .b(n_11636), .o(n_12953) );
in01f80 g558283 ( .a(n_12300), .o(n_12301) );
no02f80 g558284 ( .a(n_11635), .b(n_11634), .o(n_12300) );
na02f80 g558285 ( .a(n_11635), .b(n_11634), .o(n_12952) );
in01f80 g558286 ( .a(n_12298), .o(n_12299) );
no02f80 g558287 ( .a(n_11633), .b(n_11632), .o(n_12298) );
na02f80 g558288 ( .a(n_11633), .b(n_11632), .o(n_12956) );
in01f80 g558289 ( .a(n_12296), .o(n_12297) );
no02f80 g558290 ( .a(n_11631), .b(n_11630), .o(n_12296) );
na02f80 g558291 ( .a(n_11631), .b(n_11630), .o(n_12955) );
in01f80 g558292 ( .a(n_12294), .o(n_12295) );
no02f80 g558293 ( .a(n_11626), .b(n_11625), .o(n_12294) );
na02f80 g558294 ( .a(n_11628), .b(n_11627), .o(n_11629) );
na02f80 g558295 ( .a(n_11626), .b(n_11625), .o(n_12959) );
na02f80 g558296 ( .a(n_9512), .b(n_900), .o(n_11624) );
no02f80 g558297 ( .a(n_10122), .b(n_10121), .o(n_10123) );
in01f80 g558298 ( .a(n_12292), .o(n_12293) );
no02f80 g558299 ( .a(n_11623), .b(n_11622), .o(n_12292) );
na02f80 g558300 ( .a(n_11623), .b(n_11622), .o(n_12951) );
in01f80 g558301 ( .a(n_11020), .o(n_11021) );
no02f80 g558302 ( .a(n_10120), .b(n_10119), .o(n_11020) );
na02f80 g558303 ( .a(n_10120), .b(n_10119), .o(n_12122) );
in01f80 g558304 ( .a(n_11018), .o(n_11019) );
no02f80 g558305 ( .a(n_10118), .b(n_10117), .o(n_11018) );
na02f80 g558306 ( .a(n_10118), .b(n_10117), .o(n_12121) );
in01f80 g558307 ( .a(n_11016), .o(n_11017) );
no02f80 g558308 ( .a(n_10116), .b(n_10115), .o(n_11016) );
na02f80 g558309 ( .a(n_10116), .b(n_10115), .o(n_12120) );
in01f80 g558310 ( .a(n_11014), .o(n_11015) );
no02f80 g558311 ( .a(n_10114), .b(n_10113), .o(n_11014) );
na02f80 g558312 ( .a(n_10114), .b(n_10113), .o(n_12134) );
in01f80 g558313 ( .a(n_11012), .o(n_11013) );
no02f80 g558314 ( .a(n_10112), .b(n_10111), .o(n_11012) );
na02f80 g558315 ( .a(n_10112), .b(n_10111), .o(n_12133) );
in01f80 g558316 ( .a(n_11010), .o(n_11011) );
na02f80 g558317 ( .a(n_10110), .b(n_10109), .o(n_11010) );
no02f80 g558318 ( .a(n_10110), .b(n_10109), .o(n_12138) );
in01f80 g558319 ( .a(n_11008), .o(n_11009) );
no02f80 g558320 ( .a(n_10108), .b(n_10107), .o(n_11008) );
in01f80 g558321 ( .a(n_11621), .o(n_12556) );
no02f80 g558322 ( .a(n_11007), .b(n_11006), .o(n_11621) );
na02f80 g558323 ( .a(n_10989), .b(x_in_0_5), .o(n_12548) );
in01f80 g558324 ( .a(n_15868), .o(n_12947) );
na02f80 g558325 ( .a(n_11823), .b(x_in_24_0), .o(n_15868) );
na02f80 g558326 ( .a(n_10108), .b(n_10107), .o(n_12137) );
na02f80 g558327 ( .a(n_10104), .b(n_10103), .o(n_12129) );
na02f80 g558328 ( .a(n_11007), .b(n_11006), .o(n_12555) );
in01f80 g558329 ( .a(n_11004), .o(n_11005) );
no02f80 g558330 ( .a(n_10092), .b(n_10091), .o(n_11004) );
na02f80 g558331 ( .a(n_10106), .b(n_10105), .o(n_12132) );
in01f80 g558332 ( .a(n_11002), .o(n_11003) );
no02f80 g558333 ( .a(n_10106), .b(n_10105), .o(n_11002) );
na02f80 g558334 ( .a(n_10102), .b(n_10101), .o(n_12130) );
in01f80 g558335 ( .a(n_11000), .o(n_11001) );
no02f80 g558336 ( .a(n_10104), .b(n_10103), .o(n_11000) );
in01f80 g558337 ( .a(n_10998), .o(n_10999) );
no02f80 g558338 ( .a(n_10102), .b(n_10101), .o(n_10998) );
na02f80 g558339 ( .a(n_9204), .b(n_4097), .o(n_10997) );
na02f80 g558340 ( .a(n_10334), .b(n_8387), .o(n_13747) );
in01f80 g558341 ( .a(n_11619), .o(n_11620) );
na02f80 g558342 ( .a(n_10996), .b(n_9198), .o(n_11619) );
na02f80 g558343 ( .a(n_9386), .b(n_9385), .o(n_12126) );
in01f80 g558344 ( .a(n_10994), .o(n_10995) );
no02f80 g558345 ( .a(n_9386), .b(n_9385), .o(n_10994) );
na02f80 g558346 ( .a(n_10100), .b(n_10099), .o(n_12125) );
in01f80 g558347 ( .a(n_10992), .o(n_10993) );
no02f80 g558348 ( .a(n_10100), .b(n_10099), .o(n_10992) );
na02f80 g558349 ( .a(n_10098), .b(n_10097), .o(n_12140) );
in01f80 g558350 ( .a(n_10990), .o(n_10991) );
no02f80 g558351 ( .a(n_10098), .b(n_10097), .o(n_10990) );
in01f80 g558352 ( .a(n_11617), .o(n_11618) );
no02f80 g558353 ( .a(n_10989), .b(x_in_0_5), .o(n_11617) );
no02f80 g558354 ( .a(n_10987), .b(n_10986), .o(n_10988) );
na02f80 g558355 ( .a(n_8809), .b(n_8807), .o(n_8808) );
na02f80 g558356 ( .a(n_10984), .b(n_10983), .o(n_10985) );
no02f80 g558357 ( .a(n_8897), .b(n_7169), .o(n_11078) );
na03f80 g558358 ( .a(n_15228), .b(n_7984), .c(FE_OFN419_n_16909), .o(n_11145) );
na02f80 g558359 ( .a(n_9359), .b(n_6517), .o(n_9360) );
in01f80 g558360 ( .a(n_12290), .o(n_12291) );
na02f80 g558361 ( .a(n_11616), .b(n_11615), .o(n_12290) );
no02f80 g558362 ( .a(n_11616), .b(n_11615), .o(n_12960) );
in01f80 g558363 ( .a(n_11613), .o(n_11614) );
na02f80 g558364 ( .a(n_10976), .b(n_10975), .o(n_11613) );
na02f80 g558365 ( .a(n_10333), .b(n_1300), .o(n_12289) );
in01f80 g558366 ( .a(n_16510), .o(n_12513) );
na02f80 g558367 ( .a(n_13117), .b(x_in_56_0), .o(n_16510) );
na02f80 g558368 ( .a(n_9414), .b(n_20), .o(n_11612) );
in01f80 g558369 ( .a(n_10981), .o(n_10982) );
na02f80 g558370 ( .a(n_10096), .b(n_10095), .o(n_10981) );
in01f80 g558371 ( .a(n_10979), .o(n_10980) );
no02f80 g558372 ( .a(n_10096), .b(n_10095), .o(n_10979) );
no02f80 g558373 ( .a(n_10094), .b(n_8589), .o(n_13285) );
no02f80 g558374 ( .a(n_10130), .b(n_9357), .o(n_9358) );
no02f80 g558375 ( .a(n_8902), .b(n_10973), .o(n_11366) );
na02f80 g558376 ( .a(n_10093), .b(x_in_4_5), .o(n_12131) );
in01f80 g558377 ( .a(n_10977), .o(n_10978) );
no02f80 g558378 ( .a(n_10093), .b(x_in_4_5), .o(n_10977) );
no02f80 g558379 ( .a(n_11610), .b(n_11609), .o(n_11611) );
no02f80 g558380 ( .a(n_10976), .b(n_10975), .o(n_12540) );
no02f80 g558381 ( .a(n_11676), .b(n_10973), .o(n_10974) );
na02f80 g558382 ( .a(n_10971), .b(n_10970), .o(n_10972) );
in01f80 g558383 ( .a(n_11607), .o(n_11608) );
na02f80 g558384 ( .a(n_10969), .b(n_9202), .o(n_11607) );
no02f80 g558385 ( .a(n_9196), .b(n_9203), .o(n_23562) );
na02f80 g558386 ( .a(n_10092), .b(n_10091), .o(n_12139) );
na02f80 g558387 ( .a(n_9355), .b(n_9354), .o(n_9356) );
na02f80 g558388 ( .a(n_10089), .b(n_10088), .o(n_10090) );
in01f80 g558389 ( .a(n_11606), .o(n_13725) );
na02f80 g558390 ( .a(n_10968), .b(n_8385), .o(n_11606) );
no02f80 g558391 ( .a(n_9194), .b(x_in_1_7), .o(n_11373) );
na02f80 g558392 ( .a(n_11604), .b(n_11603), .o(n_11605) );
na02f80 g558393 ( .a(n_11657), .b(n_12288), .o(n_11602) );
no02f80 g558394 ( .a(n_10086), .b(n_10085), .o(n_10087) );
na02f80 g558395 ( .a(n_10166), .b(n_10083), .o(n_10084) );
na02f80 g558396 ( .a(n_8082), .b(n_5432), .o(n_13484) );
in01f80 g558397 ( .a(n_10966), .o(n_10967) );
no02f80 g558398 ( .a(n_10082), .b(n_10081), .o(n_10966) );
na02f80 g558399 ( .a(n_10082), .b(n_10081), .o(n_12094) );
no02f80 g558400 ( .a(n_10126), .b(n_9352), .o(n_9353) );
no02f80 g558401 ( .a(n_11584), .b(x_in_39_9), .o(n_12537) );
na02f80 g558402 ( .a(n_10080), .b(n_10079), .o(n_12106) );
in01f80 g558403 ( .a(n_10964), .o(n_10965) );
no02f80 g558404 ( .a(n_10080), .b(n_10079), .o(n_10964) );
no02f80 g558405 ( .a(n_10128), .b(n_9350), .o(n_9351) );
na02f80 g558406 ( .a(n_10077), .b(n_10076), .o(n_10078) );
no02f80 g558407 ( .a(n_10963), .b(n_10962), .o(n_25654) );
na02f80 g558408 ( .a(n_10075), .b(FE_OFN28_n_13676), .o(n_11075) );
in01f80 g558409 ( .a(n_11600), .o(n_11601) );
na02f80 g558410 ( .a(n_10961), .b(n_9184), .o(n_11600) );
na02f80 g558411 ( .a(n_10074), .b(n_10073), .o(n_12103) );
in01f80 g558412 ( .a(n_10959), .o(n_10960) );
no02f80 g558413 ( .a(n_10074), .b(n_10073), .o(n_10959) );
na02f80 g558414 ( .a(n_11598), .b(n_11597), .o(n_11599) );
na02f80 g558415 ( .a(n_11595), .b(n_11594), .o(n_11596) );
no02f80 g558416 ( .a(n_9404), .b(n_7929), .o(n_11769) );
na02f80 g558417 ( .a(n_8077), .b(n_5427), .o(n_13481) );
na02f80 g558418 ( .a(n_10957), .b(n_10956), .o(n_10958) );
in01f80 g558419 ( .a(n_10954), .o(n_10955) );
na02f80 g558420 ( .a(n_10072), .b(n_10071), .o(n_10954) );
no02f80 g558421 ( .a(n_10072), .b(n_10071), .o(n_12101) );
in01f80 g558422 ( .a(n_10952), .o(n_10953) );
na02f80 g558423 ( .a(n_10070), .b(n_10069), .o(n_10952) );
no02f80 g558424 ( .a(n_10070), .b(n_10069), .o(n_12100) );
na02f80 g558425 ( .a(n_8967), .b(n_6636), .o(n_13478) );
in01f80 g558426 ( .a(n_14034), .o(n_10068) );
na02f80 g558427 ( .a(n_8080), .b(n_5064), .o(n_14034) );
na02f80 g558428 ( .a(n_8079), .b(n_5422), .o(n_13475) );
na02f80 g558429 ( .a(n_8081), .b(n_5424), .o(n_13472) );
in01f80 g558430 ( .a(n_14037), .o(n_10067) );
na02f80 g558431 ( .a(n_8078), .b(n_5423), .o(n_14037) );
no02f80 g558432 ( .a(n_10951), .b(n_10950), .o(n_12561) );
in01f80 g558433 ( .a(n_12098), .o(n_11593) );
na02f80 g558434 ( .a(n_10951), .b(n_10950), .o(n_12098) );
na02f80 g558435 ( .a(n_10949), .b(n_10948), .o(n_12534) );
in01f80 g558436 ( .a(n_11591), .o(n_11592) );
no02f80 g558437 ( .a(n_10949), .b(n_10948), .o(n_11591) );
na02f80 g558438 ( .a(n_12343), .b(n_12342), .o(n_10947) );
na02f80 g558439 ( .a(n_11590), .b(n_9556), .o(n_22568) );
na02f80 g558440 ( .a(n_10945), .b(n_10944), .o(n_10946) );
in01f80 g558441 ( .a(n_10942), .o(n_10943) );
no02f80 g558442 ( .a(n_10066), .b(n_10065), .o(n_10942) );
na02f80 g558443 ( .a(n_10066), .b(n_10065), .o(n_12096) );
in01f80 g558444 ( .a(n_10940), .o(n_10941) );
na02f80 g558445 ( .a(n_10064), .b(n_10063), .o(n_10940) );
no02f80 g558446 ( .a(n_10064), .b(n_10063), .o(n_12095) );
no02f80 g558447 ( .a(n_10938), .b(n_10937), .o(n_10939) );
na02f80 g558448 ( .a(n_8606), .b(n_5759), .o(n_13469) );
in01f80 g558449 ( .a(n_11588), .o(n_11589) );
na02f80 g558450 ( .a(n_10936), .b(n_9176), .o(n_11588) );
no02f80 g558451 ( .a(n_10062), .b(n_10061), .o(n_12832) );
in01f80 g558452 ( .a(n_10934), .o(n_10935) );
no02f80 g558453 ( .a(n_10060), .b(n_10059), .o(n_10934) );
in01f80 g558454 ( .a(n_10932), .o(n_10933) );
na02f80 g558455 ( .a(n_10060), .b(n_10059), .o(n_10932) );
no02f80 g558456 ( .a(n_9363), .b(n_9348), .o(n_9349) );
na02f80 g558457 ( .a(n_10057), .b(n_10056), .o(n_10058) );
in01f80 g558458 ( .a(n_11586), .o(n_11587) );
na02f80 g558459 ( .a(n_10931), .b(n_10930), .o(n_11586) );
no02f80 g558460 ( .a(n_10931), .b(n_10930), .o(n_12531) );
oa12f80 g558461 ( .a(n_8433), .b(n_8355), .c(FE_OFN236_n_4162), .o(n_10929) );
oa12f80 g558462 ( .a(n_8435), .b(n_8352), .c(FE_OFN240_n_4162), .o(n_10928) );
oa12f80 g558463 ( .a(n_8431), .b(n_8350), .c(FE_OFN306_n_3069), .o(n_10927) );
oa12f80 g558464 ( .a(n_8429), .b(n_8351), .c(FE_OFN303_n_3069), .o(n_10926) );
oa12f80 g558465 ( .a(n_8437), .b(n_8353), .c(FE_OFN258_n_4280), .o(n_10925) );
oa12f80 g558466 ( .a(n_8427), .b(n_8354), .c(FE_OFN293_n_3069), .o(n_10924) );
na02f80 g558467 ( .a(n_11584), .b(n_4514), .o(n_11585) );
na02f80 g558468 ( .a(n_10054), .b(n_10053), .o(n_10055) );
no02f80 g558469 ( .a(n_10052), .b(x_in_7_9), .o(n_11359) );
na02f80 g558470 ( .a(n_10339), .b(n_12288), .o(n_16131) );
na02f80 g558471 ( .a(n_10922), .b(x_in_1_7), .o(n_10923) );
in01f80 g558472 ( .a(n_12530), .o(n_11583) );
na02f80 g558473 ( .a(n_10921), .b(n_10920), .o(n_12530) );
in01f80 g558474 ( .a(n_11581), .o(n_11582) );
no02f80 g558475 ( .a(n_10921), .b(n_10920), .o(n_11581) );
no02f80 g558476 ( .a(n_11580), .b(n_11579), .o(n_14102) );
no02f80 g558477 ( .a(n_12313), .b(n_11579), .o(n_10919) );
na02f80 g558478 ( .a(n_11670), .b(n_10918), .o(n_12087) );
na02f80 g558479 ( .a(n_11666), .b(n_10917), .o(n_12089) );
na02f80 g558480 ( .a(n_11668), .b(n_10916), .o(n_12088) );
na02f80 g558481 ( .a(n_11672), .b(n_10915), .o(n_12086) );
na02f80 g558482 ( .a(n_11662), .b(n_10914), .o(n_12084) );
na02f80 g558483 ( .a(n_11664), .b(n_10913), .o(n_12085) );
in01f80 g558484 ( .a(n_10911), .o(n_10912) );
no02f80 g558485 ( .a(n_9388), .b(n_9387), .o(n_10911) );
na02f80 g558486 ( .a(n_9388), .b(n_9387), .o(n_12083) );
no02f80 g558487 ( .a(n_11697), .b(n_10050), .o(n_10051) );
na02f80 g558488 ( .a(n_11697), .b(n_10048), .o(n_10049) );
na02f80 g558489 ( .a(n_10046), .b(n_10045), .o(n_10047) );
na02f80 g558490 ( .a(n_15247), .b(FE_OFN290_n_27194), .o(n_11770) );
na02f80 g558491 ( .a(n_10043), .b(n_10042), .o(n_10044) );
in01f80 g558492 ( .a(n_11577), .o(n_11578) );
no02f80 g558493 ( .a(n_10910), .b(n_10909), .o(n_11577) );
na02f80 g558494 ( .a(n_10910), .b(n_10909), .o(n_12512) );
no02f80 g558495 ( .a(n_10041), .b(x_in_27_10), .o(n_11351) );
no02f80 g558496 ( .a(n_10039), .b(n_13246), .o(n_10040) );
no02f80 g558497 ( .a(n_10907), .b(n_13251), .o(n_10908) );
in01f80 g558498 ( .a(n_11575), .o(n_11576) );
no02f80 g558499 ( .a(n_10906), .b(n_10905), .o(n_11575) );
na02f80 g558500 ( .a(n_10906), .b(n_10905), .o(n_12511) );
na02f80 g558501 ( .a(n_10037), .b(n_10036), .o(n_10038) );
na02f80 g558502 ( .a(n_10034), .b(n_10033), .o(n_10035) );
no02f80 g558503 ( .a(n_10903), .b(n_10902), .o(n_10904) );
na02f80 g558504 ( .a(n_10031), .b(n_10030), .o(n_10032) );
in01f80 g558505 ( .a(n_11573), .o(n_11574) );
no02f80 g558506 ( .a(n_10901), .b(n_10900), .o(n_11573) );
na02f80 g558507 ( .a(n_10901), .b(n_10900), .o(n_12510) );
no02f80 g558508 ( .a(n_10028), .b(n_10027), .o(n_10029) );
no02f80 g558509 ( .a(n_10898), .b(n_10897), .o(n_10899) );
na02f80 g558510 ( .a(n_10025), .b(n_10024), .o(n_10026) );
no02f80 g558511 ( .a(n_10023), .b(x_in_5_11), .o(n_11353) );
na02f80 g558512 ( .a(n_10021), .b(n_10020), .o(n_10022) );
na02f80 g558513 ( .a(n_10018), .b(n_10017), .o(n_10019) );
no02f80 g558514 ( .a(n_10016), .b(x_in_43_11), .o(n_11349) );
no02f80 g558515 ( .a(n_10895), .b(n_10894), .o(n_10896) );
na02f80 g558516 ( .a(n_10014), .b(n_10013), .o(n_10015) );
na02f80 g558517 ( .a(n_10011), .b(n_10010), .o(n_10012) );
na02f80 g558518 ( .a(n_10893), .b(n_10892), .o(n_12509) );
in01f80 g558519 ( .a(n_11571), .o(n_11572) );
no02f80 g558520 ( .a(n_10893), .b(n_10892), .o(n_11571) );
na02f80 g558521 ( .a(n_11569), .b(n_11568), .o(n_11570) );
na02f80 g558522 ( .a(n_11566), .b(n_11565), .o(n_11567) );
no02f80 g558523 ( .a(n_10008), .b(n_10007), .o(n_10009) );
no02f80 g558524 ( .a(n_9417), .b(n_5804), .o(n_12080) );
no02f80 g558525 ( .a(n_9418), .b(n_5803), .o(n_12508) );
no02f80 g558526 ( .a(n_10005), .b(n_10004), .o(n_10006) );
no02f80 g558527 ( .a(n_10890), .b(n_10889), .o(n_10891) );
no02f80 g558528 ( .a(n_10888), .b(n_10887), .o(n_12507) );
in01f80 g558529 ( .a(n_11563), .o(n_11564) );
na02f80 g558530 ( .a(n_10888), .b(n_10887), .o(n_11563) );
na02f80 g558531 ( .a(n_10886), .b(n_10885), .o(n_12506) );
in01f80 g558532 ( .a(n_11561), .o(n_11562) );
no02f80 g558533 ( .a(n_10886), .b(n_10885), .o(n_11561) );
in01f80 g558534 ( .a(n_12865), .o(n_12866) );
no02f80 g558535 ( .a(n_10336), .b(n_4577), .o(n_12865) );
no02f80 g558536 ( .a(n_10335), .b(n_4578), .o(n_12946) );
na02f80 g558537 ( .a(n_10002), .b(n_10001), .o(n_10003) );
na02f80 g558538 ( .a(n_9999), .b(n_9998), .o(n_10000) );
na02f80 g558539 ( .a(n_10883), .b(n_10882), .o(n_10884) );
no02f80 g558540 ( .a(n_9996), .b(n_9995), .o(n_9997) );
na02f80 g558541 ( .a(n_10880), .b(n_10879), .o(n_10881) );
no02f80 g558542 ( .a(n_9993), .b(n_9992), .o(n_9994) );
na02f80 g558543 ( .a(n_9990), .b(n_9989), .o(n_9991) );
in01f80 g558544 ( .a(n_10877), .o(n_10878) );
no02f80 g558545 ( .a(n_9988), .b(n_9987), .o(n_10877) );
na02f80 g558546 ( .a(n_10876), .b(n_10875), .o(n_12505) );
in01f80 g558547 ( .a(n_11559), .o(n_11560) );
no02f80 g558548 ( .a(n_10876), .b(n_10875), .o(n_11559) );
na02f80 g558549 ( .a(n_9988), .b(n_9987), .o(n_12073) );
na02f80 g558550 ( .a(n_10873), .b(n_10872), .o(n_10874) );
na02f80 g558551 ( .a(n_10870), .b(n_10869), .o(n_10871) );
in01f80 g558552 ( .a(n_12286), .o(n_12287) );
no02f80 g558553 ( .a(n_9431), .b(n_4544), .o(n_12286) );
no02f80 g558554 ( .a(n_9430), .b(n_4545), .o(n_12504) );
na02f80 g558555 ( .a(n_12237), .b(n_11557), .o(n_11558) );
na02f80 g558556 ( .a(n_9551), .b(n_10918), .o(n_11556) );
na02f80 g558557 ( .a(n_9549), .b(n_10917), .o(n_11555) );
na02f80 g558558 ( .a(n_9550), .b(n_10916), .o(n_11554) );
na02f80 g558559 ( .a(n_9548), .b(n_10915), .o(n_11553) );
na02f80 g558560 ( .a(n_10867), .b(n_10866), .o(n_10868) );
na02f80 g558561 ( .a(n_9547), .b(n_10913), .o(n_11552) );
na02f80 g558562 ( .a(n_9546), .b(n_10914), .o(n_11551) );
na02f80 g558563 ( .a(n_11549), .b(n_11548), .o(n_11550) );
na02f80 g558564 ( .a(n_9985), .b(n_9984), .o(n_9986) );
na02f80 g558565 ( .a(n_10968), .b(n_10864), .o(n_10865) );
no02f80 g558566 ( .a(n_10862), .b(n_10861), .o(n_10863) );
in01f80 g558567 ( .a(n_12238), .o(n_10860) );
no02f80 g558568 ( .a(n_9983), .b(n_9982), .o(n_12238) );
in01f80 g558569 ( .a(n_12284), .o(n_12285) );
na02f80 g558570 ( .a(n_11547), .b(n_9561), .o(n_12284) );
in01f80 g558571 ( .a(n_10858), .o(n_10859) );
no02f80 g558572 ( .a(n_9981), .b(n_9980), .o(n_10858) );
na02f80 g558573 ( .a(n_9981), .b(n_9980), .o(n_12067) );
na02f80 g558574 ( .a(n_10857), .b(n_10856), .o(n_12503) );
in01f80 g558575 ( .a(n_11545), .o(n_11546) );
no02f80 g558576 ( .a(n_10857), .b(n_10856), .o(n_11545) );
no02f80 g558577 ( .a(n_9978), .b(n_9977), .o(n_9979) );
in01f80 g558578 ( .a(n_10855), .o(n_12842) );
na02f80 g558579 ( .a(n_9976), .b(n_9975), .o(n_10855) );
no02f80 g558580 ( .a(n_11543), .b(n_4167), .o(n_11544) );
na02f80 g558581 ( .a(n_9973), .b(n_9972), .o(n_9974) );
na02f80 g558582 ( .a(n_9970), .b(n_9969), .o(n_9971) );
na02f80 g558583 ( .a(n_10852), .b(n_10851), .o(n_12502) );
no02f80 g558584 ( .a(n_9968), .b(n_9967), .o(n_12066) );
in01f80 g558585 ( .a(n_10853), .o(n_10854) );
na02f80 g558586 ( .a(n_9968), .b(n_9967), .o(n_10853) );
in01f80 g558587 ( .a(n_11541), .o(n_11542) );
no02f80 g558588 ( .a(n_10852), .b(n_10851), .o(n_11541) );
no02f80 g558589 ( .a(n_10850), .b(n_10849), .o(n_12501) );
in01f80 g558590 ( .a(n_11539), .o(n_11540) );
na02f80 g558591 ( .a(n_10850), .b(n_10849), .o(n_11539) );
na02f80 g558592 ( .a(n_9965), .b(n_9964), .o(n_9966) );
na02f80 g558593 ( .a(n_9962), .b(n_9961), .o(n_9963) );
in01f80 g558594 ( .a(n_12847), .o(n_11538) );
na02f80 g558595 ( .a(n_10848), .b(n_10847), .o(n_12847) );
no02f80 g558596 ( .a(n_8033), .b(n_4633), .o(n_9347) );
no02f80 g558597 ( .a(n_12282), .b(n_12281), .o(n_12283) );
no02f80 g558598 ( .a(n_10846), .b(n_10845), .o(n_12500) );
no02f80 g558599 ( .a(n_9953), .b(n_9952), .o(n_12064) );
in01f80 g558600 ( .a(n_11536), .o(n_11537) );
na02f80 g558601 ( .a(n_10846), .b(n_10845), .o(n_11536) );
na02f80 g558602 ( .a(n_9959), .b(n_9958), .o(n_9960) );
no02f80 g558603 ( .a(n_9957), .b(n_9956), .o(n_12063) );
in01f80 g558604 ( .a(n_10843), .o(n_10844) );
na02f80 g558605 ( .a(n_9957), .b(n_9956), .o(n_10843) );
na02f80 g558606 ( .a(n_9954), .b(x_in_25_3), .o(n_9955) );
in01f80 g558607 ( .a(n_10841), .o(n_10842) );
na02f80 g558608 ( .a(n_9953), .b(n_9952), .o(n_10841) );
na02f80 g558609 ( .a(n_9950), .b(n_9949), .o(n_9951) );
no02f80 g558610 ( .a(n_10840), .b(n_10839), .o(n_12498) );
no02f80 g558611 ( .a(n_9947), .b(n_9946), .o(n_9948) );
in01f80 g558612 ( .a(n_11534), .o(n_11535) );
na02f80 g558613 ( .a(n_10840), .b(n_10839), .o(n_11534) );
no02f80 g558614 ( .a(n_9944), .b(n_9943), .o(n_9945) );
in01f80 g558615 ( .a(n_12279), .o(n_12280) );
no02f80 g558616 ( .a(n_9439), .b(n_5999), .o(n_12279) );
no02f80 g558617 ( .a(n_9438), .b(n_5998), .o(n_12499) );
no02f80 g558618 ( .a(n_9941), .b(n_9940), .o(n_9942) );
no02f80 g558619 ( .a(n_9938), .b(n_9937), .o(n_9939) );
in01f80 g558620 ( .a(n_10837), .o(n_10838) );
no02f80 g558621 ( .a(n_9936), .b(n_9935), .o(n_10837) );
na02f80 g558622 ( .a(n_9936), .b(n_9935), .o(n_12062) );
na02f80 g558623 ( .a(n_10835), .b(x_in_25_13), .o(n_10836) );
in01f80 g558624 ( .a(n_10833), .o(n_10834) );
na02f80 g558625 ( .a(n_9934), .b(n_9932), .o(n_10833) );
no02f80 g558626 ( .a(n_9934), .b(n_9932), .o(n_9933) );
na02f80 g558627 ( .a(n_9930), .b(n_9929), .o(n_9931) );
no02f80 g558628 ( .a(n_10831), .b(x_in_19_12), .o(n_10832) );
no02f80 g558629 ( .a(n_10830), .b(n_10829), .o(n_12497) );
in01f80 g558630 ( .a(n_11532), .o(n_11533) );
na02f80 g558631 ( .a(n_10830), .b(n_10829), .o(n_11532) );
na02f80 g558632 ( .a(n_9537), .b(n_9538), .o(n_14041) );
na02f80 g558633 ( .a(n_9927), .b(n_9926), .o(n_9928) );
na02f80 g558634 ( .a(n_9924), .b(n_9923), .o(n_9925) );
in01f80 g558635 ( .a(n_10827), .o(n_10828) );
no02f80 g558636 ( .a(n_9922), .b(n_9921), .o(n_10827) );
na02f80 g558637 ( .a(n_9922), .b(n_9921), .o(n_12061) );
na02f80 g558638 ( .a(n_9919), .b(x_in_51_10), .o(n_9920) );
no02f80 g558639 ( .a(n_9917), .b(x_in_51_8), .o(n_9918) );
no02f80 g558640 ( .a(n_9915), .b(x_in_51_6), .o(n_9916) );
no02f80 g558641 ( .a(n_9913), .b(x_in_51_5), .o(n_9914) );
no02f80 g558642 ( .a(n_9911), .b(n_9910), .o(n_9912) );
no02f80 g558643 ( .a(n_9908), .b(n_9907), .o(n_9909) );
na02f80 g558644 ( .a(n_9905), .b(x_in_53_3), .o(n_9906) );
in01f80 g558645 ( .a(n_10825), .o(n_10826) );
no02f80 g558646 ( .a(n_9904), .b(n_9903), .o(n_10825) );
na02f80 g558647 ( .a(n_9904), .b(n_9903), .o(n_12060) );
oa12f80 g558648 ( .a(n_5421), .b(n_7132), .c(n_8476), .o(n_12836) );
na02f80 g558649 ( .a(n_9901), .b(x_in_51_9), .o(n_9902) );
na02f80 g558650 ( .a(n_9899), .b(x_in_51_7), .o(n_9900) );
no02f80 g558651 ( .a(n_10824), .b(n_10823), .o(n_12496) );
in01f80 g558652 ( .a(n_11530), .o(n_11531) );
na02f80 g558653 ( .a(n_10824), .b(n_10823), .o(n_11530) );
no02f80 g558654 ( .a(n_10821), .b(n_10820), .o(n_10822) );
na02f80 g558655 ( .a(n_11528), .b(x_in_53_13), .o(n_11529) );
na02f80 g558656 ( .a(n_9897), .b(n_9896), .o(n_9898) );
no02f80 g558657 ( .a(n_9894), .b(x_in_51_4), .o(n_9895) );
oa12f80 g558658 ( .a(n_6628), .b(n_8364), .c(n_9440), .o(n_14028) );
na02f80 g558659 ( .a(n_11526), .b(x_in_51_11), .o(n_11527) );
na02f80 g558660 ( .a(n_9892), .b(n_9891), .o(n_9893) );
na02f80 g558661 ( .a(n_9889), .b(n_9888), .o(n_9890) );
na02f80 g558662 ( .a(n_11525), .b(n_11524), .o(n_12945) );
in01f80 g558663 ( .a(n_12277), .o(n_12278) );
no02f80 g558664 ( .a(n_11525), .b(n_11524), .o(n_12277) );
na02f80 g558665 ( .a(n_12863), .b(n_12862), .o(n_12864) );
no02f80 g558666 ( .a(n_11522), .b(n_11521), .o(n_11523) );
na02f80 g558667 ( .a(n_10818), .b(n_10817), .o(n_10819) );
na02f80 g558668 ( .a(n_9532), .b(n_11520), .o(n_22271) );
na02f80 g558669 ( .a(n_9887), .b(n_9886), .o(n_12052) );
in01f80 g558670 ( .a(n_10815), .o(n_10816) );
no02f80 g558671 ( .a(n_9887), .b(n_9886), .o(n_10815) );
na02f80 g558672 ( .a(n_9529), .b(n_10814), .o(n_18396) );
na02f80 g558673 ( .a(n_9884), .b(n_9883), .o(n_9885) );
no02f80 g558674 ( .a(n_10813), .b(n_10812), .o(n_12495) );
in01f80 g558675 ( .a(n_11518), .o(n_11519) );
na02f80 g558676 ( .a(n_10813), .b(n_10812), .o(n_11518) );
in01f80 g558677 ( .a(n_11516), .o(n_11517) );
no02f80 g558678 ( .a(n_10811), .b(n_10810), .o(n_11516) );
na02f80 g558679 ( .a(n_10811), .b(n_10810), .o(n_12494) );
in01f80 g558680 ( .a(n_10808), .o(n_10809) );
no02f80 g558681 ( .a(n_8917), .b(n_7414), .o(n_10808) );
no02f80 g558682 ( .a(n_8918), .b(n_7415), .o(n_12051) );
na02f80 g558683 ( .a(n_9882), .b(n_9881), .o(n_12050) );
in01f80 g558684 ( .a(n_10806), .o(n_10807) );
no02f80 g558685 ( .a(n_9882), .b(n_9881), .o(n_10806) );
na02f80 g558686 ( .a(n_10805), .b(n_10804), .o(n_12493) );
in01f80 g558687 ( .a(n_11514), .o(n_11515) );
no02f80 g558688 ( .a(n_10805), .b(n_10804), .o(n_11514) );
in01f80 g558689 ( .a(n_10802), .o(n_10803) );
na02f80 g558690 ( .a(n_8887), .b(n_5394), .o(n_10802) );
na02f80 g558691 ( .a(n_8888), .b(n_5393), .o(n_12049) );
in01f80 g558692 ( .a(n_10800), .o(n_10801) );
na02f80 g558693 ( .a(n_8473), .b(n_4267), .o(n_10800) );
na02f80 g558694 ( .a(n_8472), .b(n_4266), .o(n_11185) );
na02f80 g558695 ( .a(n_9879), .b(n_9878), .o(n_9880) );
no02f80 g558696 ( .a(n_9876), .b(n_9875), .o(n_9877) );
no02f80 g558697 ( .a(n_10799), .b(n_10798), .o(n_12492) );
in01f80 g558698 ( .a(n_12275), .o(n_12276) );
na02f80 g558699 ( .a(n_9413), .b(n_5818), .o(n_12275) );
na02f80 g558700 ( .a(n_9412), .b(n_5819), .o(n_12491) );
in01f80 g558701 ( .a(n_11512), .o(n_11513) );
na02f80 g558702 ( .a(n_10799), .b(n_10798), .o(n_11512) );
in01f80 g558703 ( .a(n_10796), .o(n_10797) );
no02f80 g558704 ( .a(n_8913), .b(n_5404), .o(n_10796) );
no02f80 g558705 ( .a(n_8914), .b(n_5405), .o(n_12048) );
na02f80 g558706 ( .a(n_10794), .b(n_10793), .o(n_10795) );
in01f80 g558707 ( .a(n_11510), .o(n_11511) );
na02f80 g558708 ( .a(n_8883), .b(n_5816), .o(n_11510) );
na02f80 g558709 ( .a(n_8882), .b(n_5817), .o(n_12047) );
na02f80 g558710 ( .a(n_10791), .b(n_10790), .o(n_10792) );
no02f80 g558711 ( .a(n_10789), .b(n_9105), .o(n_24650) );
na02f80 g558712 ( .a(n_10788), .b(n_10787), .o(n_12490) );
in01f80 g558713 ( .a(n_12273), .o(n_12274) );
na02f80 g558714 ( .a(n_11509), .b(n_11508), .o(n_12273) );
no02f80 g558715 ( .a(n_11509), .b(n_11508), .o(n_12944) );
no02f80 g558716 ( .a(n_9346), .b(n_9345), .o(n_11175) );
in01f80 g558717 ( .a(n_11506), .o(n_11507) );
no02f80 g558718 ( .a(n_10788), .b(n_10787), .o(n_11506) );
in01f80 g558719 ( .a(n_9873), .o(n_9874) );
na02f80 g558720 ( .a(n_9346), .b(n_9345), .o(n_9873) );
in01f80 g558721 ( .a(n_12271), .o(n_12272) );
na02f80 g558722 ( .a(n_9433), .b(n_4526), .o(n_12271) );
na02f80 g558723 ( .a(n_9432), .b(n_4525), .o(n_12489) );
in01f80 g558724 ( .a(n_11504), .o(n_11505) );
na02f80 g558725 ( .a(n_10786), .b(n_10785), .o(n_11504) );
no02f80 g558726 ( .a(n_10786), .b(n_10785), .o(n_12488) );
in01f80 g558727 ( .a(n_10783), .o(n_10784) );
na02f80 g558728 ( .a(n_9872), .b(n_9871), .o(n_10783) );
no02f80 g558729 ( .a(n_9872), .b(n_9871), .o(n_12046) );
in01f80 g558730 ( .a(n_11502), .o(n_11503) );
na02f80 g558731 ( .a(n_10782), .b(n_10781), .o(n_11502) );
no02f80 g558732 ( .a(n_10782), .b(n_10781), .o(n_12487) );
na02f80 g558733 ( .a(n_8889), .b(n_10779), .o(n_10780) );
in01f80 g558734 ( .a(n_12849), .o(n_11501) );
na02f80 g558735 ( .a(n_10778), .b(n_10777), .o(n_12849) );
no02f80 g558736 ( .a(n_9869), .b(n_9868), .o(n_9870) );
no02f80 g558737 ( .a(n_10776), .b(n_10775), .o(n_12486) );
in01f80 g558738 ( .a(n_11499), .o(n_11500) );
na02f80 g558739 ( .a(n_10776), .b(n_10775), .o(n_11499) );
in01f80 g558740 ( .a(n_11497), .o(n_11498) );
no02f80 g558741 ( .a(n_10774), .b(n_10773), .o(n_11497) );
na02f80 g558742 ( .a(n_10774), .b(n_10773), .o(n_12485) );
no02f80 g558743 ( .a(n_9000), .b(FE_OFN783_n_10771), .o(n_10772) );
in01f80 g558744 ( .a(n_10769), .o(n_10770) );
na02f80 g558745 ( .a(n_9851), .b(n_9850), .o(n_10769) );
na02f80 g558746 ( .a(n_8995), .b(n_10768), .o(n_25972) );
in01f80 g558747 ( .a(n_12270), .o(n_13136) );
na02f80 g558748 ( .a(FE_OFN815_n_12310), .b(n_8275), .o(n_12270) );
na02f80 g558749 ( .a(n_9344), .b(n_9343), .o(n_11173) );
no02f80 g558750 ( .a(n_11496), .b(n_11495), .o(n_12943) );
in01f80 g558751 ( .a(n_12268), .o(n_12269) );
na02f80 g558752 ( .a(n_11496), .b(n_11495), .o(n_12268) );
oa12f80 g558753 ( .a(n_11493), .b(n_137), .c(FE_OFN69_n_27012), .o(n_11494) );
in01f80 g558754 ( .a(n_9866), .o(n_9867) );
no02f80 g558755 ( .a(n_9344), .b(n_9343), .o(n_9866) );
no02f80 g558756 ( .a(n_9864), .b(n_9863), .o(n_9865) );
na02f80 g558757 ( .a(n_10766), .b(n_10765), .o(n_10767) );
no02f80 g558758 ( .a(n_10763), .b(n_12365), .o(n_10764) );
no02f80 g558759 ( .a(n_12267), .b(n_11543), .o(n_23565) );
in01f80 g558760 ( .a(n_11491), .o(n_11492) );
no02f80 g558761 ( .a(n_8869), .b(n_6615), .o(n_11491) );
oa12f80 g558762 ( .a(FE_OFN25_n_11489), .b(n_1115), .c(FE_OFN364_n_4860), .o(n_11490) );
in01f80 g558763 ( .a(n_11487), .o(n_11488) );
no02f80 g558764 ( .a(n_10628), .b(n_10627), .o(n_11487) );
no02f80 g558765 ( .a(n_11153), .b(n_10761), .o(n_10762) );
ao12f80 g558766 ( .a(n_7912), .b(n_9166), .c(n_10956), .o(n_13756) );
no02f80 g558767 ( .a(n_10621), .b(n_10620), .o(n_14524) );
no02f80 g558768 ( .a(n_9861), .b(n_9860), .o(n_11792) );
no02f80 g558769 ( .a(n_9005), .b(n_6592), .o(n_9862) );
ao12f80 g558770 ( .a(n_9543), .b(n_8291), .c(n_11627), .o(n_13731) );
in01f80 g558771 ( .a(n_11485), .o(n_11486) );
no02f80 g558772 ( .a(n_10637), .b(n_10636), .o(n_11485) );
in01f80 g558773 ( .a(n_11483), .o(n_11484) );
no02f80 g558774 ( .a(n_10758), .b(n_10757), .o(n_11483) );
in01f80 g558775 ( .a(n_10759), .o(n_10760) );
na02f80 g558776 ( .a(n_9861), .b(n_9860), .o(n_10759) );
na02f80 g558777 ( .a(n_10758), .b(n_10757), .o(n_12135) );
na02f80 g558778 ( .a(n_9859), .b(n_9858), .o(n_12749) );
na02f80 g558779 ( .a(n_10755), .b(n_10754), .o(n_10756) );
na02f80 g558780 ( .a(n_9808), .b(n_9807), .o(n_11793) );
no02f80 g558781 ( .a(n_9820), .b(n_9819), .o(n_11807) );
no02f80 g558782 ( .a(n_10743), .b(n_10742), .o(n_12479) );
in01f80 g558783 ( .a(n_12265), .o(n_12266) );
no02f80 g558784 ( .a(n_10337), .b(n_8543), .o(n_12265) );
no02f80 g558785 ( .a(n_10338), .b(n_8544), .o(n_12942) );
oa12f80 g558786 ( .a(n_7922), .b(n_9174), .c(n_10944), .o(n_12851) );
na02f80 g558787 ( .a(n_10752), .b(n_10751), .o(n_10753) );
no02f80 g558788 ( .a(n_9856), .b(n_9855), .o(n_9857) );
in01f80 g558789 ( .a(n_12263), .o(n_12264) );
na02f80 g558790 ( .a(n_9445), .b(n_6761), .o(n_12263) );
na02f80 g558791 ( .a(n_9444), .b(n_6762), .o(n_12465) );
na02f80 g558792 ( .a(n_9434), .b(n_7578), .o(n_12097) );
na02f80 g558793 ( .a(n_9435), .b(n_7577), .o(n_12464) );
in01f80 g558794 ( .a(n_10749), .o(n_10750) );
no02f80 g558795 ( .a(n_8915), .b(n_5402), .o(n_10749) );
no02f80 g558796 ( .a(n_8916), .b(n_5403), .o(n_11937) );
no02f80 g558797 ( .a(n_9040), .b(n_6590), .o(n_9854) );
in01f80 g558798 ( .a(n_12261), .o(n_12262) );
no02f80 g558799 ( .a(n_9402), .b(n_6608), .o(n_12261) );
no02f80 g558800 ( .a(n_10747), .b(n_10746), .o(n_10748) );
in01f80 g558801 ( .a(n_10744), .o(n_10745) );
ao22s80 g558802 ( .a(n_9853), .b(n_6672), .c(n_12091), .d(n_9852), .o(n_10744) );
no02f80 g558803 ( .a(n_9851), .b(n_9850), .o(n_11803) );
in01f80 g558804 ( .a(n_11481), .o(n_11482) );
na02f80 g558805 ( .a(n_10743), .b(n_10742), .o(n_11481) );
in01f80 g558806 ( .a(n_11694), .o(n_10741) );
na02f80 g558807 ( .a(n_9849), .b(n_9848), .o(n_11694) );
in01f80 g558808 ( .a(n_11479), .o(n_11480) );
na02f80 g558809 ( .a(n_10740), .b(n_10739), .o(n_11479) );
no02f80 g558810 ( .a(n_10740), .b(n_10739), .o(n_12458) );
in01f80 g558811 ( .a(n_11477), .o(n_11478) );
no02f80 g558812 ( .a(n_10738), .b(n_10737), .o(n_11477) );
na02f80 g558813 ( .a(n_10738), .b(n_10737), .o(n_12459) );
in01f80 g558814 ( .a(n_11475), .o(n_11476) );
no02f80 g558815 ( .a(n_10736), .b(n_10735), .o(n_11475) );
na02f80 g558816 ( .a(n_10736), .b(n_10735), .o(n_12460) );
in01f80 g558817 ( .a(n_11473), .o(n_11474) );
na02f80 g558818 ( .a(n_10734), .b(n_10733), .o(n_11473) );
no02f80 g558819 ( .a(n_10734), .b(n_10733), .o(n_12461) );
na02f80 g558820 ( .a(n_8931), .b(n_8904), .o(n_10732) );
no02f80 g558821 ( .a(n_10730), .b(n_10729), .o(n_10731) );
in01f80 g558822 ( .a(n_10727), .o(n_10728) );
na02f80 g558823 ( .a(n_9810), .b(n_9809), .o(n_10727) );
oa12f80 g558824 ( .a(FE_OFN25_n_11489), .b(n_1260), .c(FE_OFN128_n_27449), .o(n_11472) );
ao12f80 g558825 ( .a(n_8374), .b(n_9552), .c(n_11603), .o(n_13738) );
in01f80 g558826 ( .a(n_12361), .o(n_11471) );
na02f80 g558827 ( .a(n_10726), .b(n_10725), .o(n_12361) );
in01f80 g558828 ( .a(n_11695), .o(n_10724) );
no02f80 g558829 ( .a(n_9847), .b(n_9846), .o(n_11695) );
in01f80 g558830 ( .a(n_11692), .o(n_10723) );
no02f80 g558831 ( .a(n_9845), .b(n_9844), .o(n_11692) );
no02f80 g558832 ( .a(n_11047), .b(FE_OFN1244_n_12940), .o(n_9843) );
in01f80 g558833 ( .a(n_12356), .o(n_11470) );
na02f80 g558834 ( .a(n_10722), .b(n_10721), .o(n_12356) );
na02f80 g558835 ( .a(n_9841), .b(n_9840), .o(n_9842) );
in01f80 g558836 ( .a(n_11468), .o(n_11469) );
no02f80 g558837 ( .a(n_8942), .b(n_5919), .o(n_11468) );
no02f80 g558838 ( .a(n_8941), .b(n_5920), .o(n_11857) );
na02f80 g558839 ( .a(n_9838), .b(n_9837), .o(n_9839) );
oa12f80 g558840 ( .a(n_10719), .b(n_780), .c(FE_OFN352_n_4860), .o(n_10720) );
in01f80 g558841 ( .a(n_11854), .o(n_11467) );
no02f80 g558842 ( .a(n_10718), .b(n_10717), .o(n_11854) );
in01f80 g558843 ( .a(n_11465), .o(n_11466) );
na02f80 g558844 ( .a(n_10718), .b(n_10717), .o(n_11465) );
no02f80 g558845 ( .a(n_9835), .b(n_9834), .o(n_9836) );
no02f80 g558846 ( .a(n_10715), .b(n_10714), .o(n_10716) );
in01f80 g558848 ( .a(n_11463), .o(n_11464) );
na03f80 g558849 ( .a(n_9797), .b(n_9796), .c(n_9798), .o(n_11463) );
no02f80 g558850 ( .a(n_10713), .b(n_10712), .o(n_12450) );
in01f80 g558851 ( .a(n_11462), .o(n_12449) );
na02f80 g558852 ( .a(n_10713), .b(n_10712), .o(n_11462) );
in01f80 g558853 ( .a(n_10710), .o(n_10711) );
no02f80 g558854 ( .a(n_9832), .b(n_9831), .o(n_10710) );
na02f80 g558855 ( .a(n_9832), .b(n_9831), .o(n_11847) );
no02f80 g558856 ( .a(n_10708), .b(n_10707), .o(n_10709) );
na02f80 g558857 ( .a(n_12260), .b(n_12259), .o(n_14981) );
na02f80 g558858 ( .a(n_11071), .b(n_10705), .o(n_10706) );
in01f80 g558859 ( .a(n_11460), .o(n_11461) );
no02f80 g558860 ( .a(n_9415), .b(n_7582), .o(n_11460) );
no02f80 g558861 ( .a(n_9416), .b(n_7583), .o(n_12448) );
no02f80 g558862 ( .a(n_10703), .b(n_10702), .o(n_10704) );
no02f80 g558863 ( .a(FE_OFN815_n_12310), .b(n_11458), .o(n_11459) );
in01f80 g558864 ( .a(n_11831), .o(n_10701) );
na02f80 g558865 ( .a(n_9830), .b(n_9829), .o(n_11831) );
in01f80 g558866 ( .a(n_10700), .o(n_11830) );
no02f80 g558867 ( .a(n_9830), .b(n_9829), .o(n_10700) );
in01f80 g558868 ( .a(n_11827), .o(n_10699) );
no02f80 g558869 ( .a(n_9828), .b(n_9827), .o(n_11827) );
in01f80 g558870 ( .a(n_10698), .o(n_11826) );
na02f80 g558871 ( .a(n_9828), .b(n_9827), .o(n_10698) );
na02f80 g558872 ( .a(n_8895), .b(n_6423), .o(n_12316) );
in01f80 g558873 ( .a(n_11127), .o(n_10697) );
na02f80 g558874 ( .a(n_9826), .b(n_9825), .o(n_11127) );
in01f80 g558875 ( .a(n_10696), .o(n_11825) );
no02f80 g558876 ( .a(n_9826), .b(n_9825), .o(n_10696) );
in01f80 g558877 ( .a(n_10694), .o(n_10695) );
no02f80 g558878 ( .a(n_8899), .b(n_6034), .o(n_10694) );
na02f80 g558879 ( .a(n_10693), .b(n_10692), .o(n_12447) );
no02f80 g558880 ( .a(n_8900), .b(n_6033), .o(n_11804) );
in01f80 g558881 ( .a(n_11456), .o(n_11457) );
no02f80 g558882 ( .a(n_10693), .b(n_10692), .o(n_11456) );
ao12f80 g558883 ( .a(n_5701), .b(n_9342), .c(n_5700), .o(n_10315) );
in01f80 g558884 ( .a(n_11454), .o(n_11455) );
na02f80 g558885 ( .a(n_10678), .b(n_10677), .o(n_11454) );
na02f80 g558886 ( .a(n_10690), .b(n_10689), .o(n_10691) );
na02f80 g558887 ( .a(n_10688), .b(n_10687), .o(n_12445) );
in01f80 g558888 ( .a(n_11452), .o(n_11453) );
no02f80 g558889 ( .a(n_10688), .b(n_10687), .o(n_11452) );
na02f80 g558890 ( .a(n_10685), .b(n_10684), .o(n_10686) );
na02f80 g558891 ( .a(n_8886), .b(n_6422), .o(n_12340) );
in01f80 g558892 ( .a(n_10682), .o(n_10683) );
no02f80 g558893 ( .a(n_8874), .b(n_6612), .o(n_10682) );
na02f80 g558894 ( .a(n_10632), .b(n_10631), .o(n_12429) );
no02f80 g558895 ( .a(n_10680), .b(n_10679), .o(n_10681) );
no02f80 g558896 ( .a(n_10678), .b(n_10677), .o(n_12446) );
no02f80 g558897 ( .a(n_10630), .b(n_10629), .o(n_12430) );
in01f80 g558898 ( .a(n_9823), .o(n_9824) );
ao22s80 g558899 ( .a(n_7200), .b(n_8811), .c(n_8810), .d(x_in_25_13), .o(n_9823) );
ao12f80 g558900 ( .a(n_7935), .b(n_9190), .c(n_10986), .o(n_13325) );
in01f80 g558901 ( .a(n_10675), .o(n_10676) );
no02f80 g558902 ( .a(n_9822), .b(n_9821), .o(n_10675) );
na02f80 g558903 ( .a(n_9822), .b(n_9821), .o(n_11802) );
in01f80 g558904 ( .a(n_10673), .o(n_10674) );
na02f80 g558905 ( .a(n_9820), .b(n_9819), .o(n_10673) );
in01f80 g558906 ( .a(n_10671), .o(n_10672) );
no02f80 g558907 ( .a(n_9818), .b(n_9817), .o(n_10671) );
na02f80 g558908 ( .a(n_9818), .b(n_9817), .o(n_12015) );
in01f80 g558909 ( .a(n_10669), .o(n_10670) );
no02f80 g558910 ( .a(n_9816), .b(n_9815), .o(n_10669) );
na02f80 g558911 ( .a(n_9816), .b(n_9815), .o(n_11801) );
na02f80 g558912 ( .a(n_10667), .b(n_10666), .o(n_10668) );
no02f80 g558913 ( .a(n_8875), .b(n_6613), .o(n_11800) );
no02f80 g558914 ( .a(n_11450), .b(n_11449), .o(n_11451) );
in01f80 g558915 ( .a(n_10664), .o(n_10665) );
na02f80 g558916 ( .a(n_8872), .b(n_6605), .o(n_10664) );
na02f80 g558917 ( .a(n_8873), .b(n_6604), .o(n_11799) );
no02f80 g558918 ( .a(n_8969), .b(n_6606), .o(n_9814) );
in01f80 g558919 ( .a(n_10662), .o(n_10663) );
no02f80 g558920 ( .a(n_8870), .b(n_6619), .o(n_10662) );
no02f80 g558921 ( .a(n_8871), .b(n_6620), .o(n_11798) );
in01f80 g558922 ( .a(n_11447), .o(n_11448) );
na02f80 g558923 ( .a(n_9407), .b(n_6635), .o(n_11447) );
na02f80 g558924 ( .a(n_9408), .b(n_6634), .o(n_12441) );
no02f80 g558925 ( .a(n_11687), .b(n_9813), .o(n_11125) );
na02f80 g558926 ( .a(n_10647), .b(n_10646), .o(n_12480) );
oa12f80 g558927 ( .a(n_10719), .b(n_758), .c(FE_OFN352_n_4860), .o(n_10661) );
na02f80 g558928 ( .a(n_9812), .b(n_9811), .o(n_11837) );
in01f80 g558929 ( .a(n_10659), .o(n_10660) );
no02f80 g558930 ( .a(n_9812), .b(n_9811), .o(n_10659) );
no02f80 g558931 ( .a(n_9810), .b(n_9809), .o(n_11794) );
in01f80 g558932 ( .a(n_10657), .o(n_10658) );
no02f80 g558933 ( .a(n_9808), .b(n_9807), .o(n_10657) );
in01f80 g558934 ( .a(n_10655), .o(n_10656) );
no02f80 g558935 ( .a(n_9806), .b(n_9805), .o(n_10655) );
na02f80 g558936 ( .a(n_9806), .b(n_9805), .o(n_11791) );
no02f80 g558937 ( .a(n_8868), .b(n_6614), .o(n_11790) );
in01f80 g558938 ( .a(n_11445), .o(n_11446) );
na02f80 g558939 ( .a(n_8867), .b(n_6625), .o(n_11445) );
na02f80 g558940 ( .a(n_8866), .b(n_6624), .o(n_11789) );
ao12f80 g558941 ( .a(n_8369), .b(n_9544), .c(n_11597), .o(n_11101) );
in01f80 g558942 ( .a(n_10653), .o(n_10654) );
no02f80 g558943 ( .a(n_8864), .b(n_6600), .o(n_10653) );
no02f80 g558944 ( .a(n_8865), .b(n_6601), .o(n_11788) );
in01f80 g558945 ( .a(n_10651), .o(n_10652) );
na02f80 g558946 ( .a(n_8862), .b(n_6622), .o(n_10651) );
na02f80 g558947 ( .a(n_8863), .b(n_6621), .o(n_11787) );
no02f80 g558948 ( .a(n_14855), .b(n_10150), .o(n_10650) );
in01f80 g558949 ( .a(n_11443), .o(n_11444) );
no02f80 g558950 ( .a(n_9405), .b(n_6632), .o(n_11443) );
no02f80 g558951 ( .a(n_9406), .b(n_6633), .o(n_12439) );
na02f80 g558952 ( .a(n_11441), .b(n_11440), .o(n_11442) );
na02f80 g558953 ( .a(n_12314), .b(FE_OFN642_n_12432), .o(n_10649) );
in01f80 g558954 ( .a(n_11819), .o(n_10648) );
no02f80 g558955 ( .a(n_9801), .b(n_9800), .o(n_11819) );
ao12f80 g558956 ( .a(n_8371), .b(n_9545), .c(n_11594), .o(n_11102) );
in01f80 g558957 ( .a(n_11438), .o(n_11439) );
no02f80 g558958 ( .a(n_10647), .b(n_10646), .o(n_11438) );
in01f80 g558959 ( .a(n_12257), .o(n_12258) );
no02f80 g558960 ( .a(n_11437), .b(n_11436), .o(n_12257) );
na02f80 g558961 ( .a(n_11437), .b(n_11436), .o(n_12934) );
in01f80 g558962 ( .a(n_12255), .o(n_12256) );
na02f80 g558963 ( .a(n_11435), .b(n_11434), .o(n_12255) );
no02f80 g558964 ( .a(n_11435), .b(n_11434), .o(n_12933) );
in01f80 g558965 ( .a(n_11432), .o(n_11433) );
no02f80 g558966 ( .a(n_10645), .b(n_10644), .o(n_11432) );
na02f80 g558967 ( .a(n_10645), .b(n_10644), .o(n_12438) );
no02f80 g558968 ( .a(n_11430), .b(n_11429), .o(n_11431) );
no02f80 g558969 ( .a(n_9401), .b(n_6609), .o(n_12437) );
in01f80 g558970 ( .a(n_12253), .o(n_12254) );
na02f80 g558971 ( .a(n_9400), .b(n_6610), .o(n_12253) );
na02f80 g558972 ( .a(n_9399), .b(n_6611), .o(n_12436) );
no02f80 g558973 ( .a(n_10641), .b(n_10640), .o(n_12481) );
in01f80 g558974 ( .a(n_10642), .o(n_10643) );
no02f80 g558975 ( .a(n_8856), .b(n_6617), .o(n_10642) );
no02f80 g558976 ( .a(n_8857), .b(n_6616), .o(n_11781) );
in01f80 g558977 ( .a(n_11427), .o(n_11428) );
na02f80 g558978 ( .a(n_10641), .b(n_10640), .o(n_11427) );
in01f80 g558979 ( .a(n_12251), .o(n_12252) );
na02f80 g558980 ( .a(n_9398), .b(n_5766), .o(n_12251) );
na02f80 g558981 ( .a(n_9397), .b(n_5767), .o(n_12472) );
in01f80 g558982 ( .a(n_12249), .o(n_12250) );
no02f80 g558983 ( .a(n_10329), .b(n_6002), .o(n_12249) );
in01f80 g558984 ( .a(n_10638), .o(n_10639) );
no02f80 g558985 ( .a(n_8853), .b(n_7569), .o(n_10638) );
no02f80 g558986 ( .a(n_10330), .b(n_6003), .o(n_12932) );
no02f80 g558987 ( .a(n_8854), .b(n_7570), .o(n_11780) );
na02f80 g558988 ( .a(n_10637), .b(n_10636), .o(n_12482) );
in01f80 g558989 ( .a(n_11693), .o(n_10635) );
no02f80 g558990 ( .a(n_9804), .b(n_9803), .o(n_11693) );
no02f80 g558991 ( .a(n_10634), .b(n_10633), .o(n_12478) );
in01f80 g558992 ( .a(n_11425), .o(n_11426) );
na02f80 g558993 ( .a(n_10634), .b(n_10633), .o(n_11425) );
in01f80 g558994 ( .a(n_11423), .o(n_11424) );
no02f80 g558995 ( .a(n_10632), .b(n_10631), .o(n_11423) );
in01f80 g558996 ( .a(n_11421), .o(n_11422) );
na02f80 g558997 ( .a(n_10630), .b(n_10629), .o(n_11421) );
in01f80 g558998 ( .a(n_11419), .o(n_11420) );
na02f80 g558999 ( .a(n_10626), .b(n_10625), .o(n_11419) );
na02f80 g559000 ( .a(n_10628), .b(n_10627), .o(n_12475) );
no02f80 g559001 ( .a(n_10626), .b(n_10625), .o(n_12457) );
na02f80 g559002 ( .a(n_10623), .b(n_10622), .o(n_10624) );
in01f80 g559003 ( .a(n_11418), .o(n_12431) );
na02f80 g559004 ( .a(n_10621), .b(n_10620), .o(n_11418) );
oa12f80 g559005 ( .a(n_8607), .b(n_7225), .c(n_6451), .o(n_9802) );
in01f80 g559006 ( .a(n_10618), .o(n_10619) );
na02f80 g559007 ( .a(n_9801), .b(n_9800), .o(n_10618) );
no02f80 g559008 ( .a(n_10616), .b(n_10615), .o(n_10617) );
oa12f80 g559009 ( .a(n_11493), .b(n_479), .c(FE_OFN190_n_28362), .o(n_11417) );
oa12f80 g559010 ( .a(n_11415), .b(n_778), .c(FE_OFN1121_rst), .o(n_11416) );
in01f80 g559011 ( .a(n_10613), .o(n_10614) );
ao22s80 g559012 ( .a(n_7971), .b(n_9621), .c(n_9620), .d(n_6331), .o(n_10613) );
oa12f80 g559013 ( .a(n_11415), .b(n_1585), .c(FE_OFN141_n_27449), .o(n_11414) );
in01f80 g559014 ( .a(n_10611), .o(n_10612) );
ao22s80 g559015 ( .a(n_7969), .b(n_9259), .c(n_9258), .d(n_6332), .o(n_10611) );
no03m80 g559016 ( .a(n_5851), .b(n_9359), .c(n_7653), .o(n_9799) );
in01f80 g559017 ( .a(n_32733), .o(n_10610) );
oa12f80 g559019 ( .a(n_8968), .b(n_7409), .c(n_6082), .o(n_10608) );
in01f80 g559020 ( .a(n_9794), .o(n_9795) );
oa22f80 g559021 ( .a(n_7185), .b(n_9254), .c(n_9255), .d(n_10311), .o(n_9794) );
in01f80 g559022 ( .a(n_10606), .o(n_10607) );
oa22f80 g559023 ( .a(n_7183), .b(n_9793), .c(n_9792), .d(n_12111), .o(n_10606) );
in01f80 g559024 ( .a(n_11372), .o(n_10605) );
oa12f80 g559025 ( .a(n_8611), .b(n_8609), .c(n_8608), .o(n_11372) );
in01f80 g559026 ( .a(n_9790), .o(n_9791) );
oa22f80 g559027 ( .a(n_7181), .b(n_9247), .c(n_10308), .d(n_9248), .o(n_9790) );
in01f80 g559028 ( .a(n_13296), .o(n_10604) );
ao12f80 g559029 ( .a(n_8289), .b(n_9554), .c(n_11548), .o(n_13296) );
in01f80 g559030 ( .a(n_9788), .o(n_9789) );
oa22f80 g559031 ( .a(n_7179), .b(n_9256), .c(n_9257), .d(n_10305), .o(n_9788) );
ao22s80 g559032 ( .a(n_8806), .b(n_4776), .c(n_4952), .d(n_4951), .o(n_9383) );
ao22s80 g559033 ( .a(n_8805), .b(n_4395), .c(n_4965), .d(n_4964), .o(n_9380) );
ao22s80 g559034 ( .a(n_8804), .b(n_4781), .c(n_5349), .d(n_5348), .o(n_9374) );
in01f80 g559035 ( .a(n_10602), .o(n_10603) );
oa22f80 g559036 ( .a(n_9787), .b(n_6503), .c(n_9786), .d(n_12107), .o(n_10602) );
ao12f80 g559037 ( .a(n_5406), .b(n_6400), .c(x_in_41_1), .o(n_13694) );
in01f80 g559038 ( .a(n_13293), .o(n_10601) );
ao12f80 g559039 ( .a(n_8273), .b(n_9558), .c(n_11568), .o(n_13293) );
in01f80 g559040 ( .a(n_13290), .o(n_10600) );
ao12f80 g559041 ( .a(n_8271), .b(n_9557), .c(n_11565), .o(n_13290) );
oa22f80 g559042 ( .a(n_8841), .b(n_5774), .c(n_9409), .d(n_10486), .o(n_11413) );
ao22s80 g559043 ( .a(n_7939), .b(n_6334), .c(n_9225), .d(n_6335), .o(n_11104) );
oa12f80 g559044 ( .a(n_10873), .b(n_13243), .c(n_10872), .o(n_13713) );
ao12f80 g559045 ( .a(n_11997), .b(n_9784), .c(n_9783), .o(n_9785) );
oa12f80 g559046 ( .a(n_8582), .b(n_8581), .c(n_9336), .o(n_11361) );
oa12f80 g559047 ( .a(n_8631), .b(n_9227), .c(n_6337), .o(n_13406) );
no02f80 g559048 ( .a(n_10057), .b(n_5194), .o(n_9782) );
ao12f80 g559049 ( .a(n_8593), .b(n_8463), .c(n_8460), .o(n_12735) );
in01f80 g559050 ( .a(n_10598), .o(n_10599) );
oa22f80 g559051 ( .a(n_7916), .b(n_9781), .c(FE_OFN1232_n_12068), .d(x_in_41_10), .o(n_10598) );
oa22f80 g559052 ( .a(n_7136), .b(n_9341), .c(n_9340), .d(n_5142), .o(n_13391) );
na02f80 g559053 ( .a(n_9156), .b(n_12019), .o(n_10597) );
na02f80 g559054 ( .a(n_8679), .b(n_9684), .o(n_9780) );
ao12f80 g559055 ( .a(FE_OFN1196_n_12016), .b(n_10386), .c(n_10387), .o(n_10596) );
oa22f80 g559056 ( .a(n_8802), .b(n_4747), .c(n_9088), .d(n_5929), .o(n_8803) );
in01f80 g559057 ( .a(n_9778), .o(n_9779) );
oa22f80 g559058 ( .a(n_7128), .b(n_9213), .c(n_9214), .d(n_10302), .o(n_9778) );
in01f80 g559059 ( .a(n_10594), .o(n_10595) );
oa22f80 g559060 ( .a(n_7900), .b(n_9632), .c(n_9633), .d(n_11343), .o(n_10594) );
ao12f80 g559061 ( .a(n_11302), .b(n_9613), .c(x_in_41_8), .o(n_9777) );
ao12f80 g559062 ( .a(n_8563), .b(n_9718), .c(n_8561), .o(n_12078) );
na02f80 g559063 ( .a(n_8717), .b(n_9584), .o(n_9776) );
ao22s80 g559064 ( .a(n_7092), .b(n_8879), .c(n_8878), .d(n_3661), .o(n_9339) );
na02f80 g559065 ( .a(n_8714), .b(n_9581), .o(n_9775) );
ao22s80 g559066 ( .a(n_7876), .b(n_9269), .c(n_9270), .d(n_10299), .o(n_13918) );
oa12f80 g559067 ( .a(n_8964), .b(FE_OFN1083_n_8877), .c(n_8876), .o(n_13168) );
ao22s80 g559068 ( .a(n_7873), .b(n_8516), .c(n_8515), .d(n_10017), .o(n_12765) );
oa12f80 g559069 ( .a(n_8076), .b(n_8523), .c(n_4385), .o(n_12714) );
in01f80 g559070 ( .a(n_12665), .o(n_9774) );
oa12f80 g559071 ( .a(n_6765), .b(n_6774), .c(n_9338), .o(n_12665) );
in01f80 g559072 ( .a(n_9772), .o(n_9773) );
oa22f80 g559073 ( .a(n_9337), .b(n_3094), .c(n_9336), .d(x_in_17_4), .o(n_9772) );
oa12f80 g559074 ( .a(n_7937), .b(n_9138), .c(n_10937), .o(n_10165) );
ao22s80 g559075 ( .a(n_7868), .b(n_8469), .c(n_8468), .d(n_9998), .o(n_13222) );
ao12f80 g559076 ( .a(n_11229), .b(n_9609), .c(x_in_41_12), .o(n_9771) );
in01f80 g559077 ( .a(n_10592), .o(n_10593) );
oa22f80 g559078 ( .a(n_7863), .b(n_9264), .c(n_9265), .d(n_10296), .o(n_10592) );
in01f80 g559079 ( .a(n_9769), .o(n_9770) );
oa22f80 g559080 ( .a(n_7061), .b(n_9234), .c(n_10293), .d(n_9235), .o(n_9769) );
oa12f80 g559081 ( .a(n_11335), .b(n_9335), .c(n_9334), .o(n_10292) );
na02f80 g559082 ( .a(n_8711), .b(n_11327), .o(n_9768) );
ao22s80 g559083 ( .a(n_8357), .b(n_8925), .c(n_8926), .d(n_5600), .o(n_13212) );
in01f80 g559084 ( .a(n_9766), .o(n_9767) );
oa22f80 g559085 ( .a(n_7046), .b(n_9333), .c(n_9332), .d(n_11323), .o(n_9766) );
oa22f80 g559086 ( .a(n_7044), .b(n_8908), .c(n_8909), .d(n_4031), .o(n_9331) );
in01f80 g559087 ( .a(n_9764), .o(n_9765) );
oa22f80 g559088 ( .a(n_7042), .b(n_9262), .c(n_10288), .d(n_9263), .o(n_9764) );
in01f80 g559089 ( .a(n_10590), .o(n_10591) );
oa22f80 g559090 ( .a(n_7851), .b(n_9634), .c(n_9635), .d(n_11317), .o(n_10590) );
in01f80 g559091 ( .a(n_11411), .o(n_11412) );
ao22s80 g559092 ( .a(n_8349), .b(n_9611), .c(n_11134), .d(n_9610), .o(n_11411) );
oa12f80 g559093 ( .a(n_8955), .b(n_8924), .c(n_7840), .o(n_12733) );
in01f80 g559094 ( .a(n_9762), .o(n_9763) );
oa22f80 g559095 ( .a(n_7033), .b(n_9237), .c(n_9238), .d(n_10285), .o(n_9762) );
in01f80 g559096 ( .a(n_9760), .o(n_9761) );
ao22s80 g559097 ( .a(n_7035), .b(n_9330), .c(n_11140), .d(n_9329), .o(n_9760) );
in01f80 g559098 ( .a(n_9758), .o(n_9759) );
ao22s80 g559099 ( .a(n_7034), .b(n_9328), .c(n_11137), .d(n_9327), .o(n_9758) );
ao22s80 g559100 ( .a(n_7839), .b(n_11410), .c(n_12937), .d(n_11409), .o(n_13932) );
in01f80 g559101 ( .a(n_9756), .o(n_9757) );
oa22f80 g559102 ( .a(n_7031), .b(n_9326), .c(n_9325), .d(n_11311), .o(n_9756) );
in01f80 g559103 ( .a(n_9754), .o(n_9755) );
oa22f80 g559104 ( .a(n_7029), .b(n_9324), .c(n_9323), .d(n_11314), .o(n_9754) );
in01f80 g559105 ( .a(n_9752), .o(n_9753) );
oa22f80 g559106 ( .a(n_7027), .b(n_9322), .c(n_9321), .d(n_11308), .o(n_9752) );
in01f80 g559107 ( .a(n_9750), .o(n_9751) );
oa22f80 g559108 ( .a(n_7039), .b(n_9320), .c(n_9319), .d(n_11305), .o(n_9750) );
in01f80 g559109 ( .a(n_9748), .o(n_9749) );
oa22f80 g559110 ( .a(n_7025), .b(n_9228), .c(n_10282), .d(n_9229), .o(n_9748) );
in01f80 g559111 ( .a(n_9746), .o(n_9747) );
oa22f80 g559112 ( .a(n_7037), .b(n_9223), .c(n_10279), .d(n_9224), .o(n_9746) );
na02f80 g559113 ( .a(n_8708), .b(n_9690), .o(n_9745) );
ao22s80 g559114 ( .a(n_9318), .b(n_5158), .c(n_6572), .d(x_in_35_1), .o(n_13174) );
in01f80 g559115 ( .a(n_9743), .o(n_9744) );
oa22f80 g559116 ( .a(n_7018), .b(n_9232), .c(n_9233), .d(n_10276), .o(n_9743) );
in01f80 g559117 ( .a(n_9741), .o(n_9742) );
oa22f80 g559118 ( .a(n_7016), .b(n_9260), .c(n_9261), .d(n_10273), .o(n_9741) );
in01f80 g559119 ( .a(n_9739), .o(n_9740) );
oa22f80 g559120 ( .a(n_7014), .b(n_9317), .c(n_9316), .d(n_11276), .o(n_9739) );
in01f80 g559121 ( .a(n_9737), .o(n_9738) );
oa22f80 g559122 ( .a(n_7010), .b(n_9315), .c(n_9314), .d(n_11288), .o(n_9737) );
in01f80 g559123 ( .a(n_10588), .o(n_10589) );
oa22f80 g559124 ( .a(n_7824), .b(n_9640), .c(n_9641), .d(n_11285), .o(n_10588) );
in01f80 g559125 ( .a(n_9735), .o(n_9736) );
oa22f80 g559126 ( .a(n_7012), .b(n_9313), .c(n_9312), .d(n_11294), .o(n_9735) );
ao22s80 g559127 ( .a(n_8801), .b(n_4663), .c(n_5704), .d(x_in_25_3), .o(n_13132) );
ao12f80 g559128 ( .a(n_7008), .b(n_7007), .c(n_9311), .o(n_13937) );
oa22f80 g559129 ( .a(n_7006), .b(n_9310), .c(n_9309), .d(n_11279), .o(n_13926) );
ao22s80 g559130 ( .a(n_7820), .b(n_9977), .c(n_8448), .d(x_in_11_11), .o(n_13906) );
in01f80 g559131 ( .a(n_9733), .o(n_9734) );
oa22f80 g559132 ( .a(n_7001), .b(n_9281), .c(n_9282), .d(n_10267), .o(n_9733) );
in01f80 g559133 ( .a(n_9731), .o(n_9732) );
oa22f80 g559134 ( .a(n_6990), .b(FE_OFN1206_n_9308), .c(n_9307), .d(n_11264), .o(n_9731) );
in01f80 g559135 ( .a(n_9729), .o(n_9730) );
oa22f80 g559136 ( .a(n_6988), .b(n_9239), .c(n_9240), .d(n_10261), .o(n_9729) );
in01f80 g559137 ( .a(n_9727), .o(n_9728) );
oa22f80 g559138 ( .a(n_9306), .b(n_6996), .c(n_9305), .d(n_11270), .o(n_9727) );
in01f80 g559139 ( .a(n_9725), .o(n_9726) );
oa22f80 g559140 ( .a(n_6998), .b(n_9304), .c(n_9303), .d(n_11267), .o(n_9725) );
in01f80 g559141 ( .a(n_9723), .o(n_9724) );
oa22f80 g559142 ( .a(n_6994), .b(n_9275), .c(n_9276), .d(n_10258), .o(n_9723) );
in01f80 g559143 ( .a(n_9721), .o(n_9722) );
oa22f80 g559144 ( .a(n_6992), .b(n_9219), .c(n_9220), .d(n_10255), .o(n_9721) );
ao12f80 g559145 ( .a(n_11154), .b(n_9647), .c(x_in_17_5), .o(n_9720) );
ao22s80 g559146 ( .a(n_7811), .b(n_9616), .c(n_9617), .d(x_in_51_12), .o(n_9719) );
in01f80 g559147 ( .a(n_10586), .o(n_10587) );
oa12f80 g559148 ( .a(n_8547), .b(n_9718), .c(n_8546), .o(n_10586) );
in01f80 g559149 ( .a(n_10584), .o(n_10585) );
oa22f80 g559150 ( .a(n_7803), .b(n_9644), .c(n_9645), .d(n_11258), .o(n_10584) );
in01f80 g559151 ( .a(n_10582), .o(n_10583) );
oa22f80 g559152 ( .a(n_7797), .b(n_9636), .c(n_9637), .d(n_11255), .o(n_10582) );
ao12f80 g559153 ( .a(n_8556), .b(n_9602), .c(n_6473), .o(n_11107) );
oa22f80 g559154 ( .a(n_6982), .b(n_9302), .c(n_8498), .d(n_9923), .o(n_12783) );
in01f80 g559155 ( .a(n_9716), .o(n_9717) );
oa22f80 g559156 ( .a(n_6980), .b(n_9230), .c(n_9231), .d(n_10247), .o(n_9716) );
ao22s80 g559157 ( .a(n_7785), .b(n_9907), .c(n_8514), .d(x_in_27_11), .o(n_13869) );
na02f80 g559158 ( .a(n_8712), .b(n_11232), .o(n_9715) );
oa12f80 g559159 ( .a(n_8085), .b(n_8467), .c(n_6350), .o(n_12741) );
ao22s80 g559160 ( .a(n_7787), .b(n_9943), .c(n_8444), .d(x_in_43_11), .o(n_13889) );
oa22f80 g559161 ( .a(n_6975), .b(n_9221), .c(n_9222), .d(n_10250), .o(n_13398) );
oa12f80 g559162 ( .a(n_8040), .b(n_8483), .c(n_8482), .o(n_13993) );
oa12f80 g559163 ( .a(n_8027), .b(n_8525), .c(n_8524), .o(n_13977) );
oa12f80 g559164 ( .a(n_9448), .b(n_9437), .c(x_in_21_2), .o(n_14647) );
ao22s80 g559165 ( .a(n_7780), .b(n_9863), .c(n_8521), .d(n_8522), .o(n_13412) );
in01f80 g559166 ( .a(n_10580), .o(n_10581) );
ao22s80 g559167 ( .a(n_7775), .b(n_9665), .c(n_11245), .d(n_9666), .o(n_10580) );
in01f80 g559168 ( .a(n_9713), .o(n_9714) );
oa22f80 g559169 ( .a(n_6962), .b(n_9271), .c(n_10244), .d(n_9272), .o(n_9713) );
na02f80 g559170 ( .a(n_8709), .b(n_11238), .o(n_9712) );
ao12f80 g559171 ( .a(n_9390), .b(n_11381), .c(n_12862), .o(n_13682) );
ao22s80 g559172 ( .a(n_8800), .b(n_5143), .c(n_10218), .d(x_in_53_3), .o(n_13205) );
na02f80 g559173 ( .a(n_8707), .b(n_11214), .o(n_9711) );
na02f80 g559174 ( .a(n_8706), .b(n_11223), .o(n_9710) );
oa12f80 g559175 ( .a(n_8119), .b(n_8464), .c(n_5979), .o(n_12737) );
ao12f80 g559176 ( .a(n_5401), .b(n_9708), .c(n_8032), .o(n_9709) );
ao22s80 g559177 ( .a(n_8335), .b(n_10615), .c(n_8928), .d(n_8929), .o(n_13389) );
in01f80 g559178 ( .a(n_10578), .o(n_10579) );
oa22f80 g559179 ( .a(n_7770), .b(n_9642), .c(n_9643), .d(n_11235), .o(n_10578) );
ao22s80 g559180 ( .a(n_7766), .b(n_9937), .c(n_8907), .d(x_in_19_11), .o(n_14942) );
no02f80 g559181 ( .a(n_9106), .b(n_12053), .o(n_10577) );
ao12f80 g559182 ( .a(n_8540), .b(FE_OFN456_n_8508), .c(x_in_3_11), .o(n_13912) );
oa12f80 g559183 ( .a(n_8548), .b(n_8518), .c(n_8517), .o(n_14000) );
ao22s80 g559184 ( .a(n_7762), .b(n_9972), .c(n_8526), .d(n_8527), .o(n_14011) );
in01f80 g559185 ( .a(n_9706), .o(n_9707) );
ao22s80 g559186 ( .a(n_9301), .b(n_5133), .c(n_6435), .d(n_6434), .o(n_9706) );
in01f80 g559187 ( .a(n_9704), .o(n_9705) );
oa22f80 g559188 ( .a(n_6944), .b(n_9300), .c(n_11220), .d(n_9299), .o(n_9704) );
in01f80 g559189 ( .a(n_11407), .o(n_11408) );
ao22s80 g559190 ( .a(n_8329), .b(n_9217), .c(n_10576), .d(n_9218), .o(n_11407) );
oa22f80 g559191 ( .a(n_6951), .b(n_9878), .c(n_8425), .d(n_8420), .o(n_13949) );
oa22f80 g559192 ( .a(n_6942), .b(n_9298), .c(n_11209), .d(n_9297), .o(n_14902) );
in01f80 g559193 ( .a(n_10574), .o(n_10575) );
ao22s80 g559194 ( .a(n_7753), .b(n_9660), .c(n_11206), .d(FE_OFN761_n_9661), .o(n_10574) );
in01f80 g559195 ( .a(n_10572), .o(n_10573) );
oa22f80 g559196 ( .a(n_7747), .b(n_9250), .c(n_10239), .d(n_9251), .o(n_10572) );
in01f80 g559197 ( .a(n_10570), .o(n_10571) );
oa22f80 g559198 ( .a(n_9703), .b(n_3105), .c(n_12425), .d(n_10486), .o(n_10570) );
in01f80 g559199 ( .a(n_9701), .o(n_9702) );
ao22s80 g559200 ( .a(n_9296), .b(n_2604), .c(n_9295), .d(x_in_9_12), .o(n_9701) );
oa22f80 g559201 ( .a(n_7741), .b(n_9284), .c(n_9285), .d(n_3647), .o(n_13207) );
in01f80 g559202 ( .a(n_11405), .o(n_11406) );
ao22s80 g559203 ( .a(n_8313), .b(n_9671), .c(n_11192), .d(n_9672), .o(n_11405) );
ao22s80 g559204 ( .a(n_8799), .b(n_4625), .c(n_4919), .d(n_4920), .o(n_9368) );
ao22s80 g559205 ( .a(FE_OFN1220_n_8798), .b(n_4249), .c(n_5353), .d(n_5354), .o(n_9377) );
ao22s80 g559206 ( .a(n_8797), .b(n_4628), .c(n_5377), .d(n_5378), .o(n_9371) );
ao12f80 g559207 ( .a(n_8535), .b(FE_OFN763_n_8501), .c(n_6921), .o(n_13351) );
in01f80 g559208 ( .a(n_10568), .o(n_10569) );
oa22f80 g559209 ( .a(n_7727), .b(n_9252), .c(n_9253), .d(n_10231), .o(n_10568) );
oa22f80 g559210 ( .a(n_6918), .b(n_9294), .c(n_11189), .d(n_9293), .o(n_13982) );
oa22f80 g559211 ( .a(n_6916), .b(n_9292), .c(n_6237), .d(n_9291), .o(n_13862) );
in01f80 g559212 ( .a(n_10566), .o(n_10567) );
ao22s80 g559213 ( .a(n_7722), .b(n_9245), .c(n_10228), .d(n_9246), .o(n_10566) );
in01f80 g559214 ( .a(n_10564), .o(n_10565) );
ao22s80 g559215 ( .a(n_7714), .b(n_9669), .c(n_11182), .d(n_9670), .o(n_10564) );
in01f80 g559216 ( .a(n_9699), .o(n_9700) );
oa22f80 g559217 ( .a(n_6888), .b(n_9290), .c(n_11179), .d(n_9289), .o(n_9699) );
in01f80 g559218 ( .a(n_10562), .o(n_10563) );
ao22s80 g559219 ( .a(n_7706), .b(n_9576), .c(n_11176), .d(n_9577), .o(n_10562) );
in01f80 g559220 ( .a(n_12247), .o(n_12248) );
ao12f80 g559221 ( .a(n_9442), .b(n_9436), .c(n_8297), .o(n_12247) );
oa12f80 g559222 ( .a(n_8529), .b(n_8898), .c(n_10214), .o(n_12798) );
oa12f80 g559223 ( .a(n_8933), .b(n_8927), .c(n_7675), .o(n_27429) );
ao22s80 g559224 ( .a(n_9288), .b(n_5136), .c(n_9287), .d(n_11226), .o(n_13352) );
oa22f80 g559225 ( .a(n_8213), .b(FE_OFN157_n_28014), .c(n_1380), .d(FE_OFN336_n_4860), .o(n_10561) );
ao22s80 g559226 ( .a(n_7661), .b(n_9677), .c(n_6245), .d(n_9676), .o(n_13945) );
in01f80 g559227 ( .a(n_12638), .o(n_12614) );
oa12f80 g559228 ( .a(n_8623), .b(n_8622), .c(FE_OFN1091_n_8621), .o(n_12638) );
in01f80 g559229 ( .a(FE_OFN989_n_13374), .o(n_10560) );
ao22s80 g559230 ( .a(n_7462), .b(n_11040), .c(n_7461), .d(x_in_55_10), .o(n_13374) );
ao12f80 g559231 ( .a(n_8154), .b(n_8153), .c(n_8605), .o(n_12198) );
oa22f80 g559232 ( .a(n_8221), .b(n_9786), .c(n_9787), .d(n_6502), .o(n_12108) );
ao22s80 g559233 ( .a(n_9292), .b(n_6915), .c(n_7482), .d(n_9291), .o(n_11187) );
oa22f80 g559234 ( .a(n_7543), .b(n_9319), .c(n_9320), .d(n_7038), .o(n_11306) );
in01f80 g559235 ( .a(n_12691), .o(n_12685) );
oa12f80 g559236 ( .a(n_8676), .b(n_8675), .c(n_8674), .o(n_12691) );
in01f80 g559237 ( .a(n_13091), .o(n_11404) );
ao12f80 g559238 ( .a(n_9084), .b(n_9083), .c(n_9082), .o(n_13091) );
in01f80 g559239 ( .a(n_12185), .o(n_9698) );
oa12f80 g559240 ( .a(n_8164), .b(n_8163), .c(n_8162), .o(n_12185) );
ao22s80 g559241 ( .a(n_10559), .b(n_9783), .c(n_9784), .d(n_10558), .o(n_11998) );
in01f80 g559242 ( .a(n_11171), .o(n_12682) );
oa12f80 g559243 ( .a(n_8620), .b(n_8619), .c(n_8618), .o(n_11171) );
in01f80 g559244 ( .a(n_12191), .o(n_9697) );
ao12f80 g559245 ( .a(n_8161), .b(n_8160), .c(FE_OFN967_n_9286), .o(n_12191) );
in01f80 g559246 ( .a(n_12202), .o(n_9696) );
ao12f80 g559247 ( .a(n_8105), .b(n_8104), .c(n_8103), .o(n_12202) );
oa12f80 g559248 ( .a(n_8094), .b(n_8093), .c(n_8092), .o(n_11375) );
ao22s80 g559249 ( .a(n_10511), .b(n_10557), .c(n_10556), .d(n_10510), .o(n_11986) );
oa22f80 g559250 ( .a(n_9064), .b(n_10555), .c(n_10554), .d(n_9063), .o(n_11977) );
ao22s80 g559251 ( .a(n_7654), .b(n_6368), .c(FE_OFN965_n_9283), .d(n_6369), .o(n_13441) );
ao22s80 g559252 ( .a(n_7668), .b(n_6361), .c(FE_OFN967_n_9286), .d(n_6362), .o(n_13447) );
oa22f80 g559253 ( .a(n_6741), .b(n_9285), .c(n_9284), .d(n_7740), .o(n_10237) );
ao12f80 g559254 ( .a(n_9076), .b(n_9075), .c(n_10553), .o(n_12639) );
no02f80 g559255 ( .a(n_8641), .b(n_11115), .o(n_9695) );
in01f80 g559256 ( .a(n_13085), .o(n_13082) );
oa12f80 g559257 ( .a(n_9074), .b(n_9073), .c(n_9072), .o(n_13085) );
oa22f80 g559258 ( .a(n_6758), .b(n_10142), .c(n_6759), .d(n_10144), .o(n_12205) );
in01f80 g559259 ( .a(n_12695), .o(n_12058) );
oa12f80 g559260 ( .a(n_8684), .b(n_8683), .c(n_8682), .o(n_12695) );
in01f80 g559261 ( .a(n_12148), .o(n_9694) );
ao12f80 g559262 ( .a(n_8128), .b(n_8127), .c(FE_OFN965_n_9283), .o(n_12148) );
oa22f80 g559263 ( .a(n_6675), .b(n_9282), .c(n_9281), .d(n_7000), .o(n_10268) );
in01f80 g559264 ( .a(n_12597), .o(n_10552) );
ao12f80 g559265 ( .a(n_8634), .b(n_8633), .c(n_8632), .o(n_12597) );
oa22f80 g559266 ( .a(n_10551), .b(n_9514), .c(n_9515), .d(n_10550), .o(n_11969) );
ao12f80 g559267 ( .a(n_8767), .b(n_8766), .c(x_in_43_10), .o(n_9693) );
in01f80 g559268 ( .a(n_12200), .o(n_9692) );
ao12f80 g559269 ( .a(n_8122), .b(n_8121), .c(FE_OFN963_n_9280), .o(n_12200) );
ao22s80 g559270 ( .a(n_10549), .b(n_9678), .c(n_9679), .d(n_10548), .o(n_12008) );
ao12f80 g559271 ( .a(n_8773), .b(n_8772), .c(x_in_27_9), .o(n_9691) );
ao12f80 g559272 ( .a(n_9122), .b(n_9121), .c(n_9120), .o(n_11859) );
oa22f80 g559273 ( .a(n_6787), .b(n_10042), .c(n_8802), .d(n_6570), .o(n_10291) );
in01f80 g559274 ( .a(n_11402), .o(n_11403) );
oa12f80 g559275 ( .a(n_9137), .b(n_9136), .c(n_9135), .o(n_11402) );
oa22f80 g559276 ( .a(n_7451), .b(n_9316), .c(n_9317), .d(n_7013), .o(n_11277) );
ao12f80 g559277 ( .a(n_8156), .b(n_8155), .c(n_8603), .o(n_12194) );
oa12f80 g559278 ( .a(n_9148), .b(n_9147), .c(n_9146), .o(n_11941) );
in01f80 g559279 ( .a(n_11400), .o(n_11401) );
oa12f80 g559280 ( .a(n_9134), .b(n_9133), .c(n_9132), .o(n_11400) );
oa12f80 g559281 ( .a(n_8138), .b(n_8137), .c(n_8602), .o(n_12199) );
oa12f80 g559282 ( .a(n_9141), .b(n_9140), .c(n_9139), .o(n_12105) );
oa12f80 g559283 ( .a(n_9189), .b(n_9188), .c(n_9187), .o(n_11861) );
in01f80 g559284 ( .a(n_10208), .o(n_12203) );
oa12f80 g559285 ( .a(n_8159), .b(n_8158), .c(n_8157), .o(n_10208) );
in01f80 g559286 ( .a(n_13521), .o(n_12246) );
ao12f80 g559287 ( .a(n_9522), .b(n_9521), .c(n_9520), .o(n_13521) );
in01f80 g559288 ( .a(n_11398), .o(n_11399) );
ao12f80 g559289 ( .a(n_9093), .b(n_9092), .c(n_9091), .o(n_11398) );
ao22s80 g559290 ( .a(n_9518), .b(n_10547), .c(n_10546), .d(n_9517), .o(n_12002) );
oa12f80 g559291 ( .a(n_8718), .b(n_9690), .c(n_9689), .o(n_11243) );
ao12f80 g559292 ( .a(n_8784), .b(n_8783), .c(x_in_7_8), .o(n_9688) );
in01f80 g559293 ( .a(n_12196), .o(n_11202) );
oa12f80 g559294 ( .a(n_8152), .b(n_8151), .c(n_8599), .o(n_12196) );
oa22f80 g559295 ( .a(n_9279), .b(n_8171), .c(n_6574), .d(n_9278), .o(n_10265) );
no02f80 g559296 ( .a(n_9020), .b(n_11838), .o(n_10545) );
ao22s80 g559297 ( .a(n_9462), .b(n_10544), .c(n_10543), .d(n_9461), .o(n_12028) );
oa22f80 g559298 ( .a(n_9687), .b(n_8715), .c(n_6587), .d(n_9686), .o(n_11292) );
ao12f80 g559299 ( .a(n_9568), .b(n_9567), .c(x_in_39_8), .o(n_11397) );
oa22f80 g559300 ( .a(n_10542), .b(n_10531), .c(n_10532), .d(n_10541), .o(n_12034) );
ao12f80 g559301 ( .a(n_8724), .b(n_8723), .c(n_8722), .o(n_11119) );
oa22f80 g559302 ( .a(n_10540), .b(n_10517), .c(n_10518), .d(n_10539), .o(n_12013) );
oa12f80 g559303 ( .a(n_8678), .b(n_9301), .c(n_8677), .o(n_12674) );
oa12f80 g559304 ( .a(n_8765), .b(n_9685), .c(n_9684), .o(n_11164) );
ao22s80 g559305 ( .a(n_10538), .b(n_9673), .c(n_9674), .d(n_10537), .o(n_11815) );
oa22f80 g559306 ( .a(n_10536), .b(n_9509), .c(n_9510), .d(n_10535), .o(n_12026) );
oa22f80 g559307 ( .a(n_6690), .b(FE_OFN404_n_28303), .c(n_104), .d(FE_OFN136_n_27449), .o(n_9277) );
no02f80 g559308 ( .a(n_9086), .b(n_11973), .o(n_10534) );
oa22f80 g559309 ( .a(n_7468), .b(n_9321), .c(n_9322), .d(n_7026), .o(n_11309) );
ao12f80 g559310 ( .a(n_12033), .b(n_10532), .c(n_10531), .o(n_10533) );
ao22s80 g559311 ( .a(n_10530), .b(n_7396), .c(n_8244), .d(n_10529), .o(n_12020) );
in01f80 g559312 ( .a(n_9682), .o(n_9683) );
ao12f80 g559313 ( .a(n_8168), .b(n_8797), .c(n_8167), .o(n_9682) );
oa22f80 g559314 ( .a(n_6734), .b(n_9276), .c(n_9275), .d(n_6993), .o(n_10259) );
in01f80 g559315 ( .a(n_11218), .o(n_12642) );
oa12f80 g559316 ( .a(n_8657), .b(n_8656), .c(n_8655), .o(n_11218) );
in01f80 g559317 ( .a(n_12187), .o(n_9681) );
ao12f80 g559318 ( .a(n_8149), .b(n_8148), .c(n_8147), .o(n_12187) );
oa22f80 g559319 ( .a(n_6688), .b(FE_OFN406_n_28303), .c(n_713), .d(FE_OFN125_n_27449), .o(n_9274) );
oa12f80 g559320 ( .a(n_12007), .b(n_9679), .c(n_9678), .o(n_9680) );
in01f80 g559321 ( .a(n_13375), .o(n_10528) );
ao12f80 g559322 ( .a(n_8758), .b(n_8757), .c(n_8756), .o(n_13375) );
oa22f80 g559323 ( .a(n_6684), .b(FE_OFN264_n_4280), .c(n_1557), .d(FE_OFN357_n_4860), .o(n_9273) );
oa22f80 g559324 ( .a(n_10527), .b(n_9451), .c(n_9452), .d(n_10526), .o(n_12005) );
ao22s80 g559325 ( .a(n_9503), .b(n_10525), .c(n_10524), .d(n_9502), .o(n_12036) );
oa22f80 g559326 ( .a(n_9677), .b(n_7660), .c(n_7544), .d(n_9676), .o(n_11098) );
no02f80 g559327 ( .a(n_9070), .b(n_11994), .o(n_10523) );
na02f80 g559328 ( .a(n_9069), .b(n_12030), .o(n_10522) );
oa22f80 g559329 ( .a(n_10521), .b(n_3010), .c(n_8216), .d(FE_OFN1256_n_10520), .o(n_11995) );
oa22f80 g559330 ( .a(n_6755), .b(n_9272), .c(n_9271), .d(n_6961), .o(n_10245) );
ao22s80 g559331 ( .a(n_6756), .b(n_9270), .c(n_9269), .d(n_7875), .o(n_10300) );
ao12f80 g559332 ( .a(n_12012), .b(n_10518), .c(n_10517), .o(n_10519) );
oa22f80 g559333 ( .a(n_9080), .b(n_10516), .c(n_10515), .d(n_9079), .o(n_11983) );
ao22s80 g559334 ( .a(n_10514), .b(n_8991), .c(n_8992), .d(n_10513), .o(n_11980) );
oa12f80 g559335 ( .a(n_11814), .b(n_9674), .c(n_9673), .o(n_9675) );
oa12f80 g559336 ( .a(n_8140), .b(n_8800), .c(n_8139), .o(n_10235) );
oa22f80 g559337 ( .a(n_6682), .b(FE_OFN303_n_3069), .c(n_666), .d(n_27709), .o(n_9268) );
ao12f80 g559338 ( .a(n_9108), .b(n_9107), .c(x_in_3_13), .o(n_12011) );
ao22s80 g559339 ( .a(n_7450), .b(n_9672), .c(n_9671), .d(n_8312), .o(n_11193) );
oa22f80 g559340 ( .a(n_7492), .b(n_9293), .c(n_9294), .d(n_6917), .o(n_11190) );
oa22f80 g559341 ( .a(n_7533), .b(n_9299), .c(n_9300), .d(n_6943), .o(n_11221) );
ao12f80 g559342 ( .a(n_11985), .b(n_10511), .c(n_10510), .o(n_10512) );
ao22s80 g559343 ( .a(n_7532), .b(n_9670), .c(n_9669), .d(n_7713), .o(n_11183) );
in01f80 g559344 ( .a(n_13373), .o(n_10509) );
ao22s80 g559345 ( .a(n_7530), .b(n_11037), .c(n_7529), .d(x_in_15_10), .o(n_13373) );
in01f80 g559346 ( .a(n_9667), .o(n_9668) );
ao12f80 g559347 ( .a(n_8136), .b(n_8806), .c(n_8135), .o(n_9667) );
ao22s80 g559348 ( .a(n_7531), .b(n_9666), .c(n_9665), .d(n_7774), .o(n_11246) );
na02f80 g559349 ( .a(n_8670), .b(n_11157), .o(n_9664) );
oa22f80 g559350 ( .a(n_7527), .b(n_9314), .c(n_9315), .d(n_7009), .o(n_11289) );
ao22s80 g559351 ( .a(n_9663), .b(n_5951), .c(n_7526), .d(n_9662), .o(n_11158) );
oa22f80 g559352 ( .a(n_10508), .b(n_9487), .c(n_9488), .d(n_10507), .o(n_11965) );
ao22s80 g559353 ( .a(n_9500), .b(FE_OFN869_n_10506), .c(n_10505), .d(n_9499), .o(n_11962) );
oa22f80 g559354 ( .a(n_10504), .b(n_3299), .c(n_8243), .d(FE_OFN656_n_10503), .o(n_11974) );
oa22f80 g559355 ( .a(n_10502), .b(n_9496), .c(n_9497), .d(FE_OFN865_n_10501), .o(n_11959) );
no02f80 g559356 ( .a(n_9060), .b(n_11952), .o(n_10500) );
ao22s80 g559357 ( .a(n_9494), .b(FE_OFN1240_n_10499), .c(n_10498), .d(n_9493), .o(n_11956) );
ao22s80 g559358 ( .a(n_7644), .b(FE_OFN761_n_9661), .c(n_9660), .d(n_7752), .o(n_11207) );
na02f80 g559359 ( .a(n_9059), .b(n_11949), .o(n_10497) );
oa22f80 g559360 ( .a(n_10496), .b(n_2973), .c(n_8212), .d(FE_OFN863_n_10495), .o(n_11953) );
no02f80 g559361 ( .a(n_9058), .b(n_11946), .o(n_10494) );
ao22s80 g559362 ( .a(n_10493), .b(n_2984), .c(n_8242), .d(FE_OFN861_n_10492), .o(n_11950) );
ao22s80 g559363 ( .a(n_8241), .b(FE_OFN1238_n_10491), .c(n_10490), .d(n_2749), .o(n_11947) );
oa22f80 g559364 ( .a(n_9168), .b(n_10489), .c(n_10488), .d(n_9167), .o(n_11944) );
ao12f80 g559365 ( .a(n_9100), .b(n_9099), .c(n_9098), .o(n_10487) );
in01f80 g559366 ( .a(n_12426), .o(n_11396) );
oa22f80 g559367 ( .a(n_8211), .b(n_10486), .c(n_9703), .d(x_in_45_12), .o(n_12426) );
in01f80 g559368 ( .a(n_12671), .o(n_10485) );
ao12f80 g559369 ( .a(n_8666), .b(n_8665), .c(n_8664), .o(n_12671) );
in01f80 g559370 ( .a(n_13372), .o(n_10484) );
ao22s80 g559371 ( .a(n_7525), .b(n_11034), .c(n_7524), .d(x_in_47_10), .o(n_13372) );
in01f80 g559372 ( .a(n_9658), .o(n_9659) );
ao12f80 g559373 ( .a(n_8132), .b(n_8805), .c(n_8131), .o(n_9658) );
in01f80 g559374 ( .a(n_10482), .o(n_10483) );
oa12f80 g559375 ( .a(n_8566), .b(n_8500), .c(n_9926), .o(n_10482) );
ao22s80 g559376 ( .a(n_7523), .b(n_9287), .c(n_9288), .d(n_5135), .o(n_11227) );
oa22f80 g559377 ( .a(n_7521), .b(x_in_17_12), .c(n_9657), .d(n_5415), .o(n_11328) );
ao22s80 g559378 ( .a(n_9656), .b(n_5418), .c(n_7522), .d(x_in_17_11), .o(n_11239) );
ao22s80 g559379 ( .a(n_9655), .b(n_5359), .c(n_7542), .d(x_in_17_10), .o(n_11233) );
ao22s80 g559380 ( .a(n_9109), .b(n_9654), .c(n_9653), .d(x_in_17_9), .o(n_11253) );
ao22s80 g559381 ( .a(n_9652), .b(n_5360), .c(n_7520), .d(x_in_17_8), .o(n_11215) );
in01f80 g559382 ( .a(n_10480), .o(n_10481) );
ao12f80 g559383 ( .a(n_8771), .b(n_8770), .c(n_8769), .o(n_10480) );
ao22s80 g559384 ( .a(n_9114), .b(n_9651), .c(n_9650), .d(x_in_17_7), .o(n_11331) );
oa12f80 g559385 ( .a(n_8921), .b(n_8919), .c(n_8920), .o(n_12767) );
oa22f80 g559386 ( .a(n_7508), .b(x_in_17_6), .c(n_9649), .d(n_5362), .o(n_11224) );
oa22f80 g559387 ( .a(n_9648), .b(x_in_17_5), .c(n_9647), .d(n_9646), .o(n_11155) );
oa12f80 g559388 ( .a(n_8663), .b(n_9337), .c(n_8662), .o(n_11340) );
oa12f80 g559389 ( .a(n_8780), .b(n_8779), .c(n_8778), .o(n_27213) );
ao22s80 g559390 ( .a(n_7637), .b(n_6357), .c(n_9226), .d(n_6358), .o(n_13400) );
ao12f80 g559391 ( .a(n_8661), .b(n_9318), .c(n_8660), .o(n_11301) );
oa22f80 g559392 ( .a(n_10479), .b(n_10477), .c(n_8238), .d(x_in_17_13), .o(n_12054) );
ao12f80 g559393 ( .a(n_9052), .b(n_10478), .c(FE_OFN554_n_9468), .o(n_11935) );
in01f80 g559394 ( .a(n_11394), .o(n_11395) );
ao22s80 g559395 ( .a(n_8236), .b(x_in_17_13), .c(n_8235), .d(n_10477), .o(n_11394) );
oa22f80 g559396 ( .a(n_7516), .b(n_9645), .c(n_9644), .d(n_7802), .o(n_11259) );
oa22f80 g559397 ( .a(n_7517), .b(n_9643), .c(n_9642), .d(n_7769), .o(n_11236) );
oa22f80 g559398 ( .a(n_10476), .b(n_9484), .c(n_9485), .d(n_10475), .o(n_11933) );
oa22f80 g559399 ( .a(n_7515), .b(n_9641), .c(n_9640), .d(n_7823), .o(n_11286) );
oa12f80 g559400 ( .a(n_9049), .b(n_10474), .c(FE_OFN552_n_9482), .o(n_11931) );
no02f80 g559401 ( .a(n_9071), .b(n_11924), .o(n_10473) );
oa22f80 g559402 ( .a(n_7636), .b(n_9639), .c(n_11903), .d(n_9638), .o(n_14340) );
ao22s80 g559403 ( .a(n_9478), .b(n_10472), .c(n_10471), .d(n_9477), .o(n_11928) );
na02f80 g559404 ( .a(n_9048), .b(n_11921), .o(n_10470) );
oa22f80 g559405 ( .a(n_7514), .b(n_9637), .c(n_9636), .d(n_7796), .o(n_11256) );
ao22s80 g559406 ( .a(n_8232), .b(FE_OFN1214_n_10469), .c(n_10468), .d(n_2978), .o(n_11925) );
no02f80 g559407 ( .a(n_9047), .b(n_11918), .o(n_10467) );
ao22s80 g559408 ( .a(n_10466), .b(n_2977), .c(n_8231), .d(FE_OFN1212_n_10465), .o(n_11922) );
oa22f80 g559409 ( .a(n_7513), .b(n_9635), .c(n_9634), .d(n_7850), .o(n_11318) );
na02f80 g559410 ( .a(n_9004), .b(n_11912), .o(n_10464) );
oa22f80 g559411 ( .a(n_10463), .b(n_2975), .c(n_8230), .d(FE_OFN704_n_10462), .o(n_11919) );
ao12f80 g559412 ( .a(n_9046), .b(n_10461), .c(n_9480), .o(n_11916) );
no02f80 g559413 ( .a(n_9023), .b(n_11909), .o(n_10460) );
oa22f80 g559414 ( .a(n_7512), .b(n_9633), .c(n_9632), .d(n_7899), .o(n_11344) );
ao22s80 g559415 ( .a(n_10459), .b(n_2985), .c(n_8229), .d(FE_OFN1210_n_10458), .o(n_11913) );
in01f80 g559416 ( .a(n_9630), .o(n_9631) );
oa22f80 g559417 ( .a(n_6796), .b(n_9267), .c(n_9266), .d(n_11150), .o(n_9630) );
oa22f80 g559418 ( .a(n_10457), .b(n_3023), .c(n_8228), .d(FE_OFN1208_n_10456), .o(n_11910) );
oa22f80 g559419 ( .a(n_9158), .b(n_10455), .c(n_10454), .d(n_9157), .o(n_11907) );
na02f80 g559420 ( .a(n_9043), .b(n_11900), .o(n_10453) );
oa22f80 g559421 ( .a(n_6677), .b(n_9265), .c(n_9264), .d(n_7862), .o(n_10297) );
oa12f80 g559422 ( .a(n_9476), .b(n_9045), .c(n_9044), .o(n_12128) );
oa22f80 g559423 ( .a(n_8247), .b(n_9638), .c(n_9639), .d(FE_OFN548_n_10452), .o(n_11904) );
no02f80 g559424 ( .a(n_9039), .b(FE_OFN1192_n_11896), .o(n_10451) );
oa22f80 g559425 ( .a(n_7511), .b(n_9266), .c(n_9267), .d(n_6795), .o(n_11151) );
in01f80 g559426 ( .a(FE_OFN1218_n_13369), .o(n_10450) );
ao22s80 g559427 ( .a(n_7549), .b(n_11698), .c(n_7548), .d(x_in_31_10), .o(n_13369) );
ao12f80 g559428 ( .a(n_9037), .b(n_10449), .c(FE_OFN546_n_9036), .o(n_11901) );
in01f80 g559429 ( .a(n_9628), .o(n_9629) );
ao12f80 g559430 ( .a(n_8126), .b(FE_OFN1220_n_8798), .c(n_8125), .o(n_9628) );
na02f80 g559431 ( .a(n_9035), .b(n_11893), .o(n_10448) );
oa12f80 g559432 ( .a(n_9033), .b(n_10447), .c(n_9032), .o(n_11897) );
oa22f80 g559433 ( .a(n_6735), .b(n_9263), .c(n_9262), .d(n_7041), .o(n_10289) );
ao12f80 g559434 ( .a(n_9031), .b(n_10446), .c(FE_OFN544_n_9030), .o(n_11894) );
ao22s80 g559435 ( .a(n_8227), .b(n_9852), .c(n_9853), .d(n_6671), .o(n_12092) );
oa22f80 g559436 ( .a(n_10445), .b(n_9490), .c(n_9491), .d(n_10444), .o(n_11891) );
oa22f80 g559437 ( .a(n_10443), .b(n_9470), .c(n_9471), .d(n_10442), .o(n_11887) );
no02f80 g559438 ( .a(n_9029), .b(n_11882), .o(n_10441) );
in01f80 g559439 ( .a(n_9626), .o(n_9627) );
ao12f80 g559440 ( .a(n_8146), .b(n_8799), .c(n_8145), .o(n_9626) );
ao12f80 g559441 ( .a(n_8764), .b(n_8763), .c(n_8762), .o(n_15538) );
oa22f80 g559442 ( .a(n_8217), .b(x_in_41_10), .c(n_9781), .d(n_7915), .o(n_12069) );
na02f80 g559443 ( .a(n_9028), .b(n_11879), .o(n_10440) );
no02f80 g559444 ( .a(n_9027), .b(n_11876), .o(n_10439) );
ao22s80 g559445 ( .a(n_10438), .b(n_2989), .c(n_8225), .d(n_10437), .o(n_11880) );
oa22f80 g559446 ( .a(n_10436), .b(n_2996), .c(n_8224), .d(n_10435), .o(n_11877) );
oa22f80 g559447 ( .a(n_9161), .b(n_10434), .c(n_10433), .d(n_9160), .o(n_11874) );
in01f80 g559448 ( .a(n_9624), .o(n_9625) );
ao12f80 g559449 ( .a(n_8124), .b(n_8804), .c(n_8123), .o(n_9624) );
ao12f80 g559450 ( .a(n_9125), .b(n_9124), .c(n_9123), .o(n_11849) );
oa22f80 g559451 ( .a(n_10432), .b(n_10426), .c(n_10427), .d(n_10431), .o(n_11871) );
oa22f80 g559452 ( .a(n_9055), .b(n_10430), .c(n_10429), .d(n_9054), .o(n_11864) );
ao12f80 g559453 ( .a(n_11870), .b(n_10427), .c(n_10426), .o(n_10428) );
oa12f80 g559454 ( .a(n_8796), .b(n_8795), .c(x_in_1_6), .o(n_11370) );
oa22f80 g559455 ( .a(n_6754), .b(n_9261), .c(n_9260), .d(n_7015), .o(n_10274) );
in01f80 g559456 ( .a(n_12045), .o(n_11393) );
oa12f80 g559457 ( .a(n_9193), .b(n_9192), .c(n_9191), .o(n_12045) );
ao22s80 g559458 ( .a(n_10425), .b(n_2982), .c(n_8245), .d(FE_OFN658_n_10424), .o(n_12031) );
ao12f80 g559459 ( .a(n_9103), .b(n_9102), .c(n_9101), .o(n_10423) );
in01f80 g559460 ( .a(n_13376), .o(n_10422) );
ao22s80 g559461 ( .a(n_7538), .b(n_11041), .c(n_7537), .d(x_in_23_10), .o(n_13376) );
oa22f80 g559462 ( .a(n_9623), .b(n_2961), .c(n_7587), .d(n_9622), .o(n_12751) );
oa22f80 g559463 ( .a(n_9259), .b(n_7968), .c(n_6676), .d(n_9258), .o(n_10317) );
oa22f80 g559464 ( .a(n_6678), .b(n_9257), .c(n_9256), .d(n_7178), .o(n_10306) );
oa22f80 g559465 ( .a(n_6681), .b(n_9255), .c(n_9254), .d(n_7184), .o(n_10312) );
oa22f80 g559466 ( .a(n_6679), .b(n_9253), .c(n_9252), .d(n_7726), .o(n_10232) );
oa22f80 g559467 ( .a(n_8222), .b(n_9792), .c(n_9793), .d(n_7182), .o(n_12112) );
oa22f80 g559468 ( .a(n_6706), .b(n_9251), .c(n_9250), .d(n_7746), .o(n_10240) );
oa22f80 g559469 ( .a(n_9621), .b(n_7970), .c(n_7494), .d(n_9620), .o(n_11368) );
oa22f80 g559470 ( .a(n_9164), .b(n_10421), .c(n_10420), .d(n_9163), .o(n_11992) );
oa12f80 g559471 ( .a(n_6588), .b(n_10419), .c(n_8284), .o(n_14535) );
in01f80 g559472 ( .a(n_11392), .o(n_12455) );
no02f80 g559473 ( .a(n_9022), .b(n_10419), .o(n_11392) );
oa22f80 g559474 ( .a(n_9025), .b(n_10418), .c(n_10417), .d(n_9024), .o(n_12043) );
ao12f80 g559475 ( .a(n_8120), .b(n_8479), .c(n_9249), .o(n_10195) );
ao12f80 g559476 ( .a(n_8687), .b(n_8686), .c(n_9095), .o(n_11334) );
oa22f80 g559477 ( .a(n_6729), .b(n_9248), .c(n_9247), .d(n_7180), .o(n_10309) );
ao22s80 g559478 ( .a(n_7040), .b(n_9246), .c(n_9245), .d(n_7721), .o(n_10229) );
ao22s80 g559479 ( .a(n_9619), .b(n_5924), .c(n_7433), .d(n_9618), .o(n_20472) );
ao22s80 g559480 ( .a(n_6699), .b(x_in_49_14), .c(n_9244), .d(n_9118), .o(n_10191) );
in01f80 g559481 ( .a(n_12647), .o(n_10416) );
ao12f80 g559482 ( .a(n_8649), .b(n_8648), .c(n_8647), .o(n_12647) );
ao22s80 g559483 ( .a(n_7491), .b(n_9617), .c(n_9616), .d(n_7810), .o(n_11262) );
ao12f80 g559484 ( .a(n_8576), .b(n_8511), .c(x_in_51_10), .o(n_13630) );
oa22f80 g559485 ( .a(n_6977), .b(n_8474), .c(n_8475), .d(n_6351), .o(n_12745) );
ao12f80 g559486 ( .a(n_8584), .b(FE_OFN1248_n_8470), .c(x_in_51_7), .o(n_12743) );
ao12f80 g559487 ( .a(n_8583), .b(n_8465), .c(x_in_51_5), .o(n_12739) );
in01f80 g559488 ( .a(n_12693), .o(n_13094) );
oa12f80 g559489 ( .a(n_8987), .b(n_8986), .c(FE_OFN1089_n_8985), .o(n_12693) );
na02f80 g559490 ( .a(n_9021), .b(n_11866), .o(n_10415) );
oa12f80 g559491 ( .a(n_8595), .b(n_10142), .c(n_6383), .o(n_13429) );
oa22f80 g559492 ( .a(n_10414), .b(n_10392), .c(n_10393), .d(n_10413), .o(n_11851) );
ao22s80 g559493 ( .a(n_7696), .b(n_6375), .c(FE_OFN963_n_9280), .d(n_6376), .o(n_13438) );
oa22f80 g559494 ( .a(n_8220), .b(FE_OFN843_n_10412), .c(n_10411), .d(n_3192), .o(n_11867) );
no02f80 g559495 ( .a(n_9019), .b(n_11844), .o(n_10410) );
in01f80 g559496 ( .a(n_12177), .o(n_11241) );
oa12f80 g559497 ( .a(n_8184), .b(n_8183), .c(n_8182), .o(n_12177) );
oa22f80 g559498 ( .a(n_9296), .b(n_8957), .c(n_7488), .d(x_in_9_12), .o(n_12217) );
in01f80 g559499 ( .a(n_10409), .o(n_12636) );
ao12f80 g559500 ( .a(n_8744), .b(n_8743), .c(n_8742), .o(n_10409) );
na02f80 g559501 ( .a(n_9018), .b(n_11841), .o(n_10408) );
oa22f80 g559502 ( .a(n_10407), .b(n_2831), .c(n_8219), .d(n_10406), .o(n_11845) );
oa22f80 g559503 ( .a(n_8246), .b(n_10405), .c(n_10404), .d(n_2829), .o(n_11842) );
in01f80 g559504 ( .a(n_10403), .o(n_12633) );
ao12f80 g559505 ( .a(n_8746), .b(n_8966), .c(n_8745), .o(n_10403) );
in01f80 g559506 ( .a(n_12174), .o(n_11250) );
oa12f80 g559507 ( .a(n_8178), .b(n_8177), .c(n_8176), .o(n_12174) );
ao22s80 g559508 ( .a(n_9389), .b(n_11409), .c(n_11410), .d(x_in_41_11), .o(n_12938) );
in01f80 g559509 ( .a(n_12180), .o(n_10402) );
ao22s80 g559510 ( .a(n_7441), .b(n_11320), .c(n_7440), .d(n_12606), .o(n_12180) );
oa22f80 g559511 ( .a(n_10401), .b(n_2992), .c(n_8223), .d(n_10400), .o(n_11839) );
in01f80 g559512 ( .a(n_12173), .o(n_9615) );
ao12f80 g559513 ( .a(n_8175), .b(n_8174), .c(n_8173), .o(n_12173) );
ao22s80 g559514 ( .a(n_7497), .b(n_9329), .c(n_9330), .d(x_in_41_9), .o(n_11141) );
oa22f80 g559515 ( .a(n_9614), .b(x_in_41_8), .c(n_9613), .d(n_9612), .o(n_11303) );
in01f80 g559516 ( .a(n_12171), .o(n_11248) );
oa12f80 g559517 ( .a(n_8187), .b(n_8186), .c(n_8185), .o(n_12171) );
oa22f80 g559518 ( .a(n_9611), .b(x_in_41_6), .c(n_7562), .d(n_9610), .o(n_11135) );
in01f80 g559519 ( .a(n_11298), .o(n_12630) );
oa12f80 g559520 ( .a(n_8752), .b(n_8751), .c(n_8750), .o(n_11298) );
in01f80 g559521 ( .a(n_11112), .o(n_12632) );
oa12f80 g559522 ( .a(n_8700), .b(n_8699), .c(n_9338), .o(n_11112) );
ao22s80 g559523 ( .a(n_9609), .b(n_9608), .c(n_9607), .d(x_in_41_12), .o(n_11230) );
no02f80 g559524 ( .a(n_9015), .b(n_11832), .o(n_10399) );
ao12f80 g559525 ( .a(n_8646), .b(n_9606), .c(n_9604), .o(n_11132) );
ao22s80 g559526 ( .a(n_9507), .b(n_10398), .c(n_10397), .d(n_9506), .o(n_12023) );
oa12f80 g559527 ( .a(n_11131), .b(n_7483), .c(n_9604), .o(n_9605) );
ao22s80 g559528 ( .a(n_9455), .b(n_10396), .c(n_10395), .d(n_9454), .o(n_11971) );
ao12f80 g559529 ( .a(n_11850), .b(n_10393), .c(n_10392), .o(n_10394) );
oa22f80 g559530 ( .a(n_10391), .b(n_3000), .c(n_8218), .d(n_10390), .o(n_11833) );
ao22s80 g559531 ( .a(n_7928), .b(n_12697), .c(n_9603), .d(n_10779), .o(n_11129) );
in01f80 g559532 ( .a(n_13928), .o(n_10389) );
ao12f80 g559533 ( .a(n_8755), .b(n_8754), .c(n_8753), .o(n_13928) );
oa12f80 g559534 ( .a(n_8667), .b(n_9335), .c(n_9594), .o(n_11336) );
in01f80 g559535 ( .a(n_11321), .o(n_12605) );
oa12f80 g559536 ( .a(n_8741), .b(n_8740), .c(n_9602), .o(n_11321) );
oa22f80 g559537 ( .a(n_10388), .b(n_10387), .c(n_10386), .d(n_10385), .o(n_12017) );
ao22s80 g559538 ( .a(n_9601), .b(n_2953), .c(n_7573), .d(FE_OFN1272_n_9600), .o(n_12726) );
in01f80 g559539 ( .a(n_12626), .o(n_11391) );
ao12f80 g559540 ( .a(n_9012), .b(n_9011), .c(n_9010), .o(n_12626) );
in01f80 g559541 ( .a(n_13004), .o(n_11390) );
ao12f80 g559542 ( .a(n_9009), .b(n_9008), .c(n_9007), .o(n_13004) );
in01f80 g559543 ( .a(n_11147), .o(n_13007) );
oa12f80 g559544 ( .a(n_8790), .b(n_9342), .c(n_8789), .o(n_11147) );
in01f80 g559545 ( .a(n_12168), .o(n_9599) );
ao12f80 g559546 ( .a(n_8107), .b(n_8801), .c(n_8106), .o(n_12168) );
in01f80 g559547 ( .a(n_13002), .o(n_11389) );
oa12f80 g559548 ( .a(n_9068), .b(n_9067), .c(n_9066), .o(n_13002) );
oa12f80 g559549 ( .a(n_8456), .b(n_8881), .c(n_8880), .o(n_12729) );
in01f80 g559550 ( .a(n_12664), .o(n_10384) );
ao12f80 g559551 ( .a(n_8695), .b(n_8694), .c(n_8693), .o(n_12664) );
ao22s80 g559552 ( .a(n_8989), .b(n_9598), .c(n_9597), .d(n_8988), .o(n_11109) );
in01f80 g559553 ( .a(n_10382), .o(n_10383) );
ao12f80 g559554 ( .a(n_8749), .b(n_8748), .c(n_8747), .o(n_10382) );
oa22f80 g559555 ( .a(n_6686), .b(FE_OFN258_n_4280), .c(n_514), .d(FE_OFN352_n_4860), .o(n_9243) );
in01f80 g559556 ( .a(n_11387), .o(n_11388) );
ao12f80 g559557 ( .a(n_9128), .b(n_9127), .c(n_9126), .o(n_11387) );
oa22f80 g559558 ( .a(n_7473), .b(n_9332), .c(n_9333), .d(n_7045), .o(n_11324) );
in01f80 g559559 ( .a(n_10189), .o(n_12166) );
oa12f80 g559560 ( .a(n_8110), .b(n_8109), .c(n_8108), .o(n_10189) );
oa22f80 g559561 ( .a(n_8112), .b(n_9242), .c(n_8111), .d(n_9241), .o(n_11782) );
oa22f80 g559562 ( .a(n_7476), .b(n_9309), .c(n_9310), .d(n_7005), .o(n_11280) );
in01f80 g559563 ( .a(n_11121), .o(n_12618) );
oa22f80 g559564 ( .a(n_7470), .b(n_4069), .c(n_7471), .d(n_8041), .o(n_11121) );
oa22f80 g559565 ( .a(n_6702), .b(n_9240), .c(n_9239), .d(n_6987), .o(n_10262) );
oa22f80 g559566 ( .a(n_6718), .b(n_9238), .c(n_9237), .d(n_7032), .o(n_10286) );
oa22f80 g559567 ( .a(n_7472), .b(n_9325), .c(n_9326), .d(n_7030), .o(n_11312) );
ao12f80 g559568 ( .a(n_8721), .b(n_8720), .c(n_8719), .o(n_11124) );
oa22f80 g559569 ( .a(n_7469), .b(n_9323), .c(n_9324), .d(n_7028), .o(n_11315) );
ao12f80 g559570 ( .a(n_8733), .b(n_8732), .c(n_8731), .o(n_11161) );
in01f80 g559571 ( .a(n_9595), .o(n_9596) );
ao12f80 g559572 ( .a(n_8197), .b(n_8196), .c(n_8195), .o(n_9595) );
in01f80 g559573 ( .a(n_10380), .o(n_10381) );
oa12f80 g559574 ( .a(n_8727), .b(n_8726), .c(n_8725), .o(n_10380) );
in01f80 g559575 ( .a(n_11196), .o(n_12687) );
oa22f80 g559576 ( .a(n_7564), .b(n_9334), .c(n_7565), .d(n_9594), .o(n_11196) );
oa22f80 g559577 ( .a(n_9593), .b(n_5964), .c(n_7558), .d(n_9592), .o(n_11116) );
oa22f80 g559578 ( .a(n_6712), .b(FE_OFN293_n_3069), .c(n_145), .d(FE_OFN1141_n_27012), .o(n_9236) );
in01f80 g559579 ( .a(n_12443), .o(n_12245) );
no02f80 g559580 ( .a(n_9457), .b(n_9057), .o(n_12443) );
in01f80 g559581 ( .a(n_10378), .o(n_10379) );
ao12f80 g559582 ( .a(n_8739), .b(n_8738), .c(n_8737), .o(n_10378) );
oa22f80 g559583 ( .a(n_6710), .b(n_9235), .c(n_9234), .d(n_7060), .o(n_10294) );
in01f80 g559584 ( .a(n_10376), .o(n_10377) );
oa12f80 g559585 ( .a(n_8736), .b(n_8735), .c(n_8734), .o(n_10376) );
in01f80 g559586 ( .a(n_10374), .o(n_10375) );
ao12f80 g559587 ( .a(n_8730), .b(n_8729), .c(n_8728), .o(n_10374) );
oa12f80 g559588 ( .a(n_8644), .b(n_8643), .c(n_9582), .o(n_11095) );
ao12f80 g559589 ( .a(n_9131), .b(n_9130), .c(n_9129), .o(n_11777) );
oa12f80 g559590 ( .a(n_9173), .b(n_9172), .c(n_9171), .o(n_12118) );
in01f80 g559591 ( .a(n_12617), .o(n_10373) );
oa12f80 g559592 ( .a(n_8638), .b(n_8637), .c(n_8636), .o(n_12617) );
in01f80 g559593 ( .a(n_10371), .o(n_10372) );
oa12f80 g559594 ( .a(n_8703), .b(n_8702), .c(n_8701), .o(n_10371) );
oa12f80 g559595 ( .a(n_8777), .b(n_8776), .c(x_in_5_10), .o(n_11364) );
oa22f80 g559596 ( .a(n_6703), .b(n_9233), .c(n_9232), .d(n_7017), .o(n_10277) );
ao22s80 g559597 ( .a(n_9524), .b(n_10370), .c(n_10369), .d(n_9523), .o(n_11885) );
in01f80 g559598 ( .a(n_12243), .o(n_12244) );
ao12f80 g559599 ( .a(n_9542), .b(n_9541), .c(n_9540), .o(n_12243) );
oa22f80 g559600 ( .a(n_6714), .b(n_9231), .c(n_9230), .d(n_6979), .o(n_10248) );
in01f80 g559601 ( .a(n_12969), .o(n_11386) );
oa12f80 g559602 ( .a(n_8973), .b(n_8972), .c(n_8971), .o(n_12969) );
oa22f80 g559603 ( .a(n_10368), .b(n_2979), .c(n_8226), .d(n_10367), .o(n_11883) );
oa22f80 g559604 ( .a(n_7460), .b(n_9305), .c(n_9306), .d(n_6995), .o(n_11271) );
ao12f80 g559605 ( .a(n_8116), .b(n_8115), .c(n_8114), .o(n_12183) );
oa22f80 g559606 ( .a(n_7459), .b(n_9312), .c(n_9313), .d(n_7011), .o(n_11295) );
ao22s80 g559607 ( .a(n_9002), .b(n_9591), .c(n_9590), .d(n_9001), .o(n_11355) );
in01f80 g559608 ( .a(n_10365), .o(n_10366) );
ao12f80 g559609 ( .a(n_8692), .b(n_8691), .c(n_8690), .o(n_10365) );
oa22f80 g559610 ( .a(n_6700), .b(n_9229), .c(n_9228), .d(n_7024), .o(n_10283) );
in01f80 g559611 ( .a(n_12161), .o(n_9589) );
ao12f80 g559612 ( .a(n_8102), .b(n_8101), .c(FE_OFN787_n_8855), .o(n_12161) );
oa22f80 g559613 ( .a(n_8688), .b(n_9588), .c(n_9587), .d(n_6578), .o(n_11379) );
in01f80 g559614 ( .a(n_12601), .o(n_10364) );
ao12f80 g559615 ( .a(n_8630), .b(n_9396), .c(n_8629), .o(n_12601) );
in01f80 g559616 ( .a(n_12159), .o(n_9586) );
oa12f80 g559617 ( .a(n_8100), .b(n_8099), .c(n_9227), .o(n_12159) );
in01f80 g559618 ( .a(n_10184), .o(n_12156) );
oa12f80 g559619 ( .a(n_8098), .b(n_8097), .c(n_8858), .o(n_10184) );
in01f80 g559620 ( .a(n_10362), .o(n_10363) );
ao12f80 g559621 ( .a(n_8480), .b(n_9249), .c(n_10194), .o(n_10362) );
in01f80 g559622 ( .a(n_12155), .o(n_9585) );
oa12f80 g559623 ( .a(n_8130), .b(n_8129), .c(n_8859), .o(n_12155) );
in01f80 g559624 ( .a(n_12600), .o(n_10361) );
oa12f80 g559625 ( .a(n_8673), .b(n_8672), .c(n_8671), .o(n_12600) );
in01f80 g559626 ( .a(n_12977), .o(n_11385) );
ao12f80 g559627 ( .a(n_8999), .b(n_8998), .c(n_9053), .o(n_12977) );
in01f80 g559628 ( .a(n_13030), .o(n_12980) );
oa12f80 g559629 ( .a(n_9078), .b(n_9077), .c(n_9419), .o(n_13030) );
ao12f80 g559630 ( .a(n_8997), .b(n_8996), .c(n_9403), .o(n_12598) );
in01f80 g559631 ( .a(n_12629), .o(n_11384) );
oa12f80 g559632 ( .a(n_8984), .b(n_8983), .c(n_8982), .o(n_12629) );
in01f80 g559633 ( .a(n_10199), .o(n_12153) );
oa22f80 g559634 ( .a(n_6697), .b(n_11103), .c(n_6698), .d(n_9226), .o(n_10199) );
in01f80 g559635 ( .a(n_12210), .o(n_12150) );
oa12f80 g559636 ( .a(n_8096), .b(n_8095), .c(n_9225), .o(n_12210) );
oa12f80 g559637 ( .a(n_8761), .b(n_9584), .c(n_9583), .o(n_11274) );
in01f80 g559638 ( .a(n_13368), .o(n_10360) );
ao22s80 g559639 ( .a(n_7505), .b(n_11696), .c(n_7504), .d(x_in_63_10), .o(n_13368) );
oa22f80 g559640 ( .a(n_6694), .b(n_9224), .c(n_9223), .d(n_7036), .o(n_10280) );
oa22f80 g559641 ( .a(n_6695), .b(n_9222), .c(n_9221), .d(n_6974), .o(n_10251) );
in01f80 g559642 ( .a(n_10358), .o(n_10359) );
oa12f80 g559643 ( .a(n_8439), .b(n_11094), .c(n_9582), .o(n_10358) );
oa22f80 g559644 ( .a(n_6745), .b(n_9220), .c(n_9219), .d(n_6991), .o(n_10256) );
ao22s80 g559645 ( .a(n_7550), .b(n_9327), .c(n_9328), .d(x_in_41_7), .o(n_11138) );
ao22s80 g559646 ( .a(n_6696), .b(n_9218), .c(n_9217), .d(n_8328), .o(n_10242) );
in01f80 g559647 ( .a(n_10356), .o(n_10357) );
oa12f80 g559648 ( .a(n_8698), .b(n_8697), .c(n_8696), .o(n_10356) );
oa22f80 g559649 ( .a(n_7458), .b(n_9303), .c(n_9304), .d(n_6997), .o(n_11268) );
ao12f80 g559650 ( .a(n_8194), .b(n_8193), .c(n_8192), .o(n_25601) );
oa12f80 g559651 ( .a(n_8759), .b(n_9581), .c(n_9580), .o(n_11283) );
ao22s80 g559652 ( .a(n_9474), .b(n_10355), .c(n_10354), .d(n_9473), .o(n_11889) );
oa22f80 g559653 ( .a(n_9216), .b(n_8169), .c(n_6459), .d(n_9215), .o(n_10271) );
in01f80 g559654 ( .a(n_12587), .o(n_11383) );
oa12f80 g559655 ( .a(n_8979), .b(n_8978), .c(FE_OFN1274_n_8977), .o(n_12587) );
oa22f80 g559656 ( .a(n_7452), .b(n_9307), .c(FE_OFN1206_n_9308), .d(n_6989), .o(n_11265) );
in01f80 g559657 ( .a(n_12641), .o(n_11382) );
oa12f80 g559658 ( .a(n_9090), .b(n_9089), .c(n_9088), .o(n_12641) );
in01f80 g559659 ( .a(n_12583), .o(n_10353) );
oa12f80 g559660 ( .a(n_8626), .b(n_8625), .c(n_8624), .o(n_12583) );
oa22f80 g559661 ( .a(n_7539), .b(n_9289), .c(n_9290), .d(n_6887), .o(n_11180) );
in01f80 g559662 ( .a(n_12580), .o(n_12984) );
oa12f80 g559663 ( .a(n_8976), .b(n_8975), .c(FE_OFN1087_n_8974), .o(n_12580) );
oa12f80 g559664 ( .a(n_8713), .b(n_9311), .c(x_in_41_5), .o(n_11092) );
in01f80 g559665 ( .a(n_12576), .o(n_10352) );
ao12f80 g559666 ( .a(n_8652), .b(n_8651), .c(n_8650), .o(n_12576) );
in01f80 g559667 ( .a(n_12176), .o(n_9579) );
ao12f80 g559668 ( .a(n_8181), .b(n_8180), .c(n_8179), .o(n_12176) );
in01f80 g559669 ( .a(n_12146), .o(n_9578) );
oa12f80 g559670 ( .a(n_8091), .b(n_8090), .c(n_8089), .o(n_12146) );
ao22s80 g559671 ( .a(n_7561), .b(n_9577), .c(n_9576), .d(n_7705), .o(n_11177) );
in01f80 g559672 ( .a(n_12164), .o(n_9575) );
ao12f80 g559673 ( .a(n_8088), .b(n_8087), .c(n_8086), .o(n_12164) );
oa22f80 g559674 ( .a(n_7202), .b(n_9214), .c(n_9213), .d(n_7127), .o(n_10303) );
oa12f80 g559675 ( .a(n_8144), .b(n_8143), .c(n_8142), .o(n_11376) );
oa12f80 g559676 ( .a(n_9182), .b(n_9181), .c(n_9180), .o(n_12114) );
ao22s80 g559677 ( .a(n_9341), .b(n_7135), .c(n_7547), .d(n_9340), .o(n_11347) );
oa22f80 g559678 ( .a(n_7436), .b(n_9297), .c(n_9298), .d(n_6941), .o(n_11210) );
ao22s80 g559679 ( .a(n_9459), .b(n_10351), .c(n_10350), .d(n_9458), .o(n_11835) );
oa22f80 g559680 ( .a(n_6742), .b(FE_OFN234_n_4162), .c(n_1515), .d(FE_OFN101_n_27449), .o(n_9212) );
oa22f80 g559681 ( .a(n_6721), .b(FE_OFN311_n_3069), .c(n_1173), .d(FE_OFN336_n_4860), .o(n_9211) );
oa22f80 g559682 ( .a(n_6757), .b(FE_OFN248_n_4162), .c(n_315), .d(FE_OFN91_n_27449), .o(n_9210) );
ao22s80 g559683 ( .a(n_9155), .b(n_7270), .c(n_8434), .d(n_6021), .o(n_9574) );
ao22s80 g559684 ( .a(n_9153), .b(n_6492), .c(n_8432), .d(n_6023), .o(n_9573) );
ao22s80 g559685 ( .a(n_9154), .b(n_7272), .c(n_8426), .d(n_4523), .o(n_9572) );
ao22s80 g559686 ( .a(n_9152), .b(n_7315), .c(n_8436), .d(n_6022), .o(n_9571) );
ao22s80 g559687 ( .a(n_9151), .b(n_7241), .c(n_8430), .d(n_4498), .o(n_9570) );
ao22s80 g559688 ( .a(n_9150), .b(n_8200), .c(n_8428), .d(n_4884), .o(n_9569) );
ao22s80 g559689 ( .a(n_8458), .b(n_8459), .c(n_9208), .d(n_9207), .o(n_9209) );
ao22s80 g559690 ( .a(n_7898), .b(x_in_17_14), .c(n_7897), .d(n_4794), .o(n_25659) );
no02f80 g559710 ( .a(n_9567), .b(x_in_39_8), .o(n_9568) );
na02f80 g559711 ( .a(n_16002), .b(FE_OFN30_n_13676), .o(n_11415) );
na02f80 g559712 ( .a(n_9206), .b(n_9205), .o(n_14112) );
no02f80 g559713 ( .a(n_11627), .b(n_9543), .o(n_9359) );
no02f80 g559714 ( .a(n_8196), .b(n_8195), .o(n_8197) );
na02f80 g559715 ( .a(n_8795), .b(x_in_1_6), .o(n_8796) );
in01f80 g559716 ( .a(n_9203), .o(n_9204) );
no02f80 g559717 ( .a(n_8788), .b(n_8787), .o(n_9203) );
no02f80 g559718 ( .a(n_8794), .b(n_8588), .o(n_10094) );
no02f80 g559719 ( .a(n_9566), .b(n_8419), .o(n_11522) );
na02f80 g559720 ( .a(n_8792), .b(x_in_4_4), .o(n_10996) );
na02f80 g559721 ( .a(n_8793), .b(x_in_0_4), .o(n_10969) );
in01f80 g559722 ( .a(n_9201), .o(n_9202) );
no02f80 g559723 ( .a(n_8793), .b(x_in_0_4), .o(n_9201) );
in01f80 g559724 ( .a(n_9564), .o(n_9565) );
na02f80 g559725 ( .a(n_9200), .b(n_7957), .o(n_9564) );
in01f80 g559726 ( .a(n_10348), .o(n_10349) );
na02f80 g559727 ( .a(n_9563), .b(n_8403), .o(n_10348) );
na02f80 g559728 ( .a(n_7927), .b(FE_OFN30_n_13676), .o(n_10719) );
na02f80 g559729 ( .a(n_8610), .b(n_6534), .o(n_14073) );
in01f80 g559730 ( .a(n_14147), .o(n_9199) );
na02f80 g559731 ( .a(n_8645), .b(n_2884), .o(n_14147) );
in01f80 g559732 ( .a(n_9197), .o(n_9198) );
no02f80 g559733 ( .a(n_8792), .b(x_in_4_4), .o(n_9197) );
na02f80 g559734 ( .a(n_9562), .b(n_8405), .o(n_19311) );
oa12f80 g559735 ( .a(n_7134), .b(n_8791), .c(n_1980), .o(n_11007) );
na02f80 g559736 ( .a(n_9342), .b(n_8789), .o(n_8790) );
in01f80 g559737 ( .a(n_9195), .o(n_9196) );
na02f80 g559738 ( .a(n_8788), .b(n_8787), .o(n_9195) );
na02f80 g559739 ( .a(n_8386), .b(FE_OFN27_n_13676), .o(n_11493) );
in01f80 g559740 ( .a(n_9194), .o(n_10922) );
na02f80 g559741 ( .a(n_8795), .b(n_521), .o(n_9194) );
na02f80 g559742 ( .a(n_9192), .b(n_9191), .o(n_9193) );
na02f80 g559743 ( .a(n_7563), .b(n_9191), .o(n_10166) );
ao12f80 g559744 ( .a(n_3848), .b(n_5627), .c(x_in_3_13), .o(n_9355) );
na02f80 g559745 ( .a(n_7936), .b(n_9190), .o(n_10987) );
na02f80 g559746 ( .a(n_9188), .b(n_9187), .o(n_9189) );
in01f80 g559747 ( .a(n_11584), .o(n_12867) );
na02f80 g559748 ( .a(n_9567), .b(n_8133), .o(n_11584) );
na02f80 g559749 ( .a(n_9186), .b(n_9185), .o(n_11547) );
in01f80 g559750 ( .a(n_9560), .o(n_9561) );
no02f80 g559751 ( .a(n_9186), .b(n_9185), .o(n_9560) );
no02f80 g559752 ( .a(n_7464), .b(n_6301), .o(n_10962) );
no02f80 g559753 ( .a(n_7463), .b(n_6302), .o(n_10963) );
no02f80 g559754 ( .a(n_8785), .b(n_4656), .o(n_8786) );
na02f80 g559755 ( .a(n_21415), .b(n_7934), .o(n_21106) );
no02f80 g559756 ( .a(n_8783), .b(x_in_7_8), .o(n_8784) );
in01f80 g559757 ( .a(n_9183), .o(n_9184) );
no02f80 g559758 ( .a(n_8782), .b(n_8781), .o(n_9183) );
na02f80 g559759 ( .a(n_8782), .b(n_8781), .o(n_10961) );
ao12f80 g559760 ( .a(n_3847), .b(n_6312), .c(x_in_51_13), .o(n_10089) );
na02f80 g559761 ( .a(n_8779), .b(n_8778), .o(n_8780) );
in01f80 g559762 ( .a(n_10346), .o(n_10347) );
na02f80 g559763 ( .a(n_8389), .b(n_9559), .o(n_10346) );
ao12f80 g559764 ( .a(n_4030), .b(n_4993), .c(x_in_11_13), .o(n_10130) );
no02f80 g559765 ( .a(n_8193), .b(n_8192), .o(n_8194) );
na02f80 g559766 ( .a(n_9181), .b(n_9180), .o(n_9182) );
na02f80 g559767 ( .a(n_9558), .b(n_8274), .o(n_11569) );
na02f80 g559768 ( .a(n_9557), .b(n_8272), .o(n_11566) );
oa12f80 g559769 ( .a(n_9336), .b(n_9179), .c(n_1977), .o(n_10951) );
ao22s80 g559770 ( .a(n_6670), .b(n_6330), .c(n_32730), .d(n_2256), .o(n_15457) );
na02f80 g559771 ( .a(n_9178), .b(n_9177), .o(n_11590) );
in01f80 g559772 ( .a(n_9555), .o(n_9556) );
no02f80 g559773 ( .a(n_9178), .b(n_9177), .o(n_9555) );
oa12f80 g559774 ( .a(n_8191), .b(n_8190), .c(n_2007), .o(n_10065) );
na02f80 g559775 ( .a(n_8776), .b(x_in_5_10), .o(n_8777) );
na02f80 g559776 ( .a(n_8775), .b(n_8774), .o(n_10936) );
in01f80 g559777 ( .a(n_9175), .o(n_9176) );
no02f80 g559778 ( .a(n_8775), .b(n_8774), .o(n_9175) );
na02f80 g559779 ( .a(n_9554), .b(n_8290), .o(n_11549) );
no02f80 g559780 ( .a(n_8772), .b(x_in_27_9), .o(n_8773) );
no02f80 g559781 ( .a(n_8770), .b(n_8769), .o(n_8771) );
no02f80 g559782 ( .a(n_7923), .b(n_9174), .o(n_10945) );
ao12f80 g559783 ( .a(n_3903), .b(n_6448), .c(x_in_35_13), .o(n_10077) );
oa12f80 g559784 ( .a(n_5716), .b(n_8768), .c(n_2026), .o(n_10930) );
ao12f80 g559785 ( .a(n_4080), .b(n_5615), .c(x_in_27_13), .o(n_10126) );
no02f80 g559786 ( .a(n_8766), .b(x_in_43_10), .o(n_8767) );
ao12f80 g559787 ( .a(n_3839), .b(n_5341), .c(x_in_43_13), .o(n_10128) );
na02f80 g559788 ( .a(n_9172), .b(n_9171), .o(n_9173) );
in01f80 g559789 ( .a(n_10052), .o(n_9170) );
na02f80 g559790 ( .a(n_8783), .b(n_7304), .o(n_10052) );
na02f80 g559791 ( .a(n_9553), .b(n_8379), .o(n_15665) );
ao12f80 g559792 ( .a(n_6801), .b(n_5879), .c(n_4377), .o(n_13697) );
no02f80 g559793 ( .a(n_9168), .b(n_9167), .o(n_9169) );
na02f80 g559794 ( .a(n_7913), .b(n_9166), .o(n_10957) );
na02f80 g559795 ( .a(n_9685), .b(n_9684), .o(n_8765) );
na02f80 g559796 ( .a(n_8839), .b(FE_OFN27_n_13676), .o(n_11489) );
no02f80 g559797 ( .a(n_7812), .b(n_9180), .o(n_16132) );
no02f80 g559798 ( .a(n_9164), .b(n_9163), .o(n_9165) );
no02f80 g559799 ( .a(n_9161), .b(n_9160), .o(n_9162) );
no02f80 g559800 ( .a(n_9158), .b(n_9157), .o(n_9159) );
na02f80 g559801 ( .a(n_10530), .b(n_10529), .o(n_9156) );
na02f80 g559802 ( .a(n_8375), .b(n_9552), .o(n_11604) );
in01f80 g559803 ( .a(n_11670), .o(n_9551) );
no02f80 g559804 ( .a(n_9155), .b(x_in_23_8), .o(n_11670) );
in01f80 g559805 ( .a(n_11668), .o(n_9550) );
no02f80 g559806 ( .a(n_9154), .b(x_in_63_8), .o(n_11668) );
in01f80 g559807 ( .a(n_11666), .o(n_9549) );
no02f80 g559808 ( .a(n_9153), .b(x_in_15_8), .o(n_11666) );
in01f80 g559809 ( .a(n_11672), .o(n_9548) );
no02f80 g559810 ( .a(n_9152), .b(x_in_55_8), .o(n_11672) );
in01f80 g559811 ( .a(n_11664), .o(n_9547) );
no02f80 g559812 ( .a(n_9151), .b(x_in_47_8), .o(n_11664) );
in01f80 g559813 ( .a(n_11662), .o(n_9546) );
no02f80 g559814 ( .a(n_9150), .b(x_in_31_8), .o(n_11662) );
no02f80 g559815 ( .a(n_9149), .b(x_in_8_1), .o(n_11053) );
na02f80 g559816 ( .a(n_9149), .b(x_in_8_1), .o(n_11054) );
no02f80 g559817 ( .a(n_8763), .b(n_8762), .o(n_8764) );
na02f80 g559818 ( .a(n_8372), .b(n_9545), .o(n_11595) );
na02f80 g559819 ( .a(n_8186), .b(n_8185), .o(n_8187) );
na02f80 g559820 ( .a(n_9147), .b(n_9146), .o(n_9148) );
in01f80 g559821 ( .a(n_10041), .o(n_9145) );
na02f80 g559822 ( .a(n_8772), .b(n_7289), .o(n_10041) );
na02f80 g559823 ( .a(n_8370), .b(n_9544), .o(n_11598) );
in01f80 g559824 ( .a(n_10023), .o(n_9144) );
na02f80 g559825 ( .a(n_8776), .b(n_5388), .o(n_10023) );
na02f80 g559826 ( .a(n_9584), .b(n_9583), .o(n_8761) );
no02f80 g559827 ( .a(n_7883), .b(n_9143), .o(n_21148) );
no02f80 g559828 ( .a(n_6778), .b(n_6638), .o(n_8760) );
in01f80 g559829 ( .a(n_10016), .o(n_9142) );
na02f80 g559830 ( .a(n_8766), .b(n_6496), .o(n_10016) );
na02f80 g559831 ( .a(n_9581), .b(n_9580), .o(n_8759) );
ao12f80 g559832 ( .a(n_3398), .b(n_6289), .c(x_in_7_13), .o(n_10057) );
no02f80 g559833 ( .a(n_8757), .b(n_8756), .o(n_8758) );
no02f80 g559834 ( .a(n_8292), .b(n_9543), .o(n_11628) );
no02f80 g559835 ( .a(n_8754), .b(n_8753), .o(n_8755) );
na02f80 g559836 ( .a(n_9140), .b(n_9139), .o(n_9141) );
na02f80 g559837 ( .a(n_8751), .b(n_8750), .o(n_8752) );
na02f80 g559838 ( .a(n_7108), .b(n_7111), .o(n_20672) );
no02f80 g559839 ( .a(n_8748), .b(n_8747), .o(n_8749) );
ao12f80 g559840 ( .a(n_3834), .b(n_5595), .c(x_in_59_13), .o(n_9363) );
na02f80 g559841 ( .a(n_8183), .b(n_8182), .o(n_8184) );
no02f80 g559842 ( .a(n_8966), .b(n_8745), .o(n_8746) );
no02f80 g559843 ( .a(n_8180), .b(n_8179), .o(n_8181) );
na02f80 g559844 ( .a(n_8177), .b(n_8176), .o(n_8178) );
no02f80 g559845 ( .a(n_8174), .b(n_8173), .o(n_8175) );
no02f80 g559846 ( .a(n_8743), .b(n_8742), .o(n_8744) );
no02f80 g559847 ( .a(n_10345), .b(n_8835), .o(n_19865) );
no02f80 g559848 ( .a(n_9138), .b(n_7938), .o(n_10938) );
na02f80 g559849 ( .a(n_8740), .b(n_9602), .o(n_8741) );
no02f80 g559850 ( .a(n_9541), .b(n_9540), .o(n_9542) );
na02f80 g559851 ( .a(n_9136), .b(n_9135), .o(n_9137) );
no02f80 g559852 ( .a(n_8738), .b(n_8737), .o(n_8739) );
na02f80 g559853 ( .a(n_8735), .b(n_8734), .o(n_8736) );
na02f80 g559854 ( .a(n_9133), .b(n_9132), .o(n_9134) );
no02f80 g559855 ( .a(n_7853), .b(n_6725), .o(n_9934) );
no02f80 g559856 ( .a(n_8732), .b(n_8731), .o(n_8733) );
no02f80 g559857 ( .a(n_8729), .b(n_8728), .o(n_8730) );
na02f80 g559858 ( .a(n_8726), .b(n_8725), .o(n_8727) );
no02f80 g559859 ( .a(n_9130), .b(n_9129), .o(n_9131) );
no02f80 g559860 ( .a(n_8723), .b(n_8722), .o(n_8724) );
no02f80 g559861 ( .a(n_9127), .b(n_9126), .o(n_9128) );
no02f80 g559862 ( .a(n_9124), .b(n_9123), .o(n_9125) );
no02f80 g559863 ( .a(n_9121), .b(n_9120), .o(n_9122) );
na02f80 g559864 ( .a(n_8901), .b(n_9118), .o(n_9119) );
no02f80 g559865 ( .a(n_8720), .b(n_8719), .o(n_8721) );
na02f80 g559866 ( .a(n_9690), .b(n_9689), .o(n_8718) );
no02f80 g559867 ( .a(n_8171), .b(n_6253), .o(n_8172) );
na02f80 g559868 ( .a(n_9583), .b(n_11273), .o(n_8717) );
no02f80 g559869 ( .a(n_8715), .b(n_6252), .o(n_8716) );
na02f80 g559870 ( .a(n_9580), .b(n_11282), .o(n_8714) );
no02f80 g559871 ( .a(n_8169), .b(n_6246), .o(n_8170) );
na02f80 g559872 ( .a(n_9311), .b(x_in_41_5), .o(n_8713) );
ao12f80 g559873 ( .a(n_3822), .b(n_5770), .c(x_in_61_13), .o(n_10043) );
in01f80 g559874 ( .a(n_9538), .o(n_9539) );
na02f80 g559875 ( .a(n_9117), .b(n_9116), .o(n_9538) );
in01f80 g559876 ( .a(n_9536), .o(n_9537) );
no02f80 g559877 ( .a(n_9117), .b(n_9116), .o(n_9536) );
na02f80 g559878 ( .a(n_9655), .b(x_in_17_10), .o(n_8712) );
na02f80 g559879 ( .a(n_9114), .b(x_in_17_7), .o(n_9115) );
na02f80 g559880 ( .a(n_9657), .b(x_in_17_12), .o(n_8711) );
no02f80 g559881 ( .a(n_8330), .b(n_32735), .o(n_9113) );
in01f80 g559882 ( .a(n_9111), .o(n_9112) );
oa12f80 g559883 ( .a(n_2735), .b(n_8710), .c(n_4153), .o(n_9111) );
na02f80 g559884 ( .a(n_9109), .b(x_in_17_9), .o(n_9110) );
no02f80 g559885 ( .a(n_9107), .b(x_in_3_13), .o(n_9108) );
na02f80 g559886 ( .a(n_9656), .b(x_in_17_11), .o(n_8709) );
na02f80 g559887 ( .a(n_9689), .b(n_11682), .o(n_8708) );
na02f80 g559888 ( .a(n_9652), .b(x_in_17_8), .o(n_8707) );
na02f80 g559889 ( .a(n_9649), .b(x_in_17_6), .o(n_8706) );
no02f80 g559890 ( .a(n_8832), .b(n_9535), .o(n_15231) );
no02f80 g559891 ( .a(n_10479), .b(x_in_17_13), .o(n_9106) );
no02f80 g559892 ( .a(n_8705), .b(n_8704), .o(n_10789) );
in01f80 g559893 ( .a(n_9104), .o(n_9105) );
na02f80 g559894 ( .a(n_8705), .b(n_8704), .o(n_9104) );
no02f80 g559895 ( .a(n_9534), .b(n_8333), .o(n_16476) );
na02f80 g559896 ( .a(n_8702), .b(n_8701), .o(n_8703) );
no02f80 g559897 ( .a(n_9102), .b(n_9101), .o(n_9103) );
no02f80 g559898 ( .a(n_9099), .b(n_9098), .o(n_9100) );
na02f80 g559899 ( .a(n_8699), .b(n_9338), .o(n_8700) );
na02f80 g559900 ( .a(n_8831), .b(n_10344), .o(n_14484) );
na02f80 g559901 ( .a(n_8323), .b(n_9533), .o(n_14019) );
na02f80 g559902 ( .a(n_9097), .b(n_9096), .o(n_11520) );
in01f80 g559903 ( .a(n_9531), .o(n_9532) );
no02f80 g559904 ( .a(n_9097), .b(n_9096), .o(n_9531) );
na02f80 g559905 ( .a(n_8697), .b(n_8696), .o(n_8698) );
in01f80 g559906 ( .a(n_9529), .o(n_9530) );
na02f80 g559907 ( .a(n_7432), .b(n_7499), .o(n_9529) );
na02f80 g559908 ( .a(n_7431), .b(n_7498), .o(n_10814) );
na02f80 g559909 ( .a(n_9528), .b(n_8315), .o(n_17409) );
no02f80 g559910 ( .a(n_8694), .b(n_8693), .o(n_8695) );
no02f80 g559911 ( .a(n_8691), .b(n_8690), .o(n_8692) );
na02f80 g559912 ( .a(n_8310), .b(n_9527), .o(n_20459) );
no02f80 g559913 ( .a(n_8688), .b(n_6249), .o(n_8689) );
no02f80 g559914 ( .a(n_8827), .b(n_9526), .o(n_19350) );
no02f80 g559915 ( .a(n_8686), .b(n_9095), .o(n_8687) );
no02f80 g559916 ( .a(n_7484), .b(n_9095), .o(n_14017) );
na02f80 g559917 ( .a(n_11381), .b(n_9391), .o(n_12863) );
no02f80 g559918 ( .a(n_7719), .b(n_9094), .o(n_20834) );
no02f80 g559919 ( .a(n_9092), .b(n_9091), .o(n_9093) );
no02f80 g559920 ( .a(n_8826), .b(n_10343), .o(n_15594) );
na02f80 g559921 ( .a(n_9089), .b(n_9088), .o(n_9090) );
no02f80 g559922 ( .a(n_8797), .b(n_8167), .o(n_8168) );
oa12f80 g559923 ( .a(n_8680), .b(n_724), .c(n_27449), .o(n_8685) );
na02f80 g559924 ( .a(n_9524), .b(n_9523), .o(n_9525) );
na02f80 g559925 ( .a(n_9601), .b(FE_OFN1272_n_9600), .o(n_9087) );
na02f80 g559926 ( .a(n_8812), .b(n_6471), .o(n_12259) );
no02f80 g559927 ( .a(n_10504), .b(FE_OFN656_n_10503), .o(n_9086) );
in01f80 g559928 ( .a(n_11678), .o(n_14881) );
na02f80 g559929 ( .a(n_8615), .b(n_8614), .o(n_11678) );
no02f80 g559930 ( .a(n_7486), .b(n_2697), .o(n_14432) );
in01f80 g559931 ( .a(n_11090), .o(n_9085) );
no02f80 g559932 ( .a(n_7495), .b(n_3002), .o(n_11090) );
no02f80 g559933 ( .a(n_9521), .b(n_9520), .o(n_9522) );
no02f80 g559934 ( .a(n_9083), .b(n_9082), .o(n_9084) );
na02f80 g559935 ( .a(n_8163), .b(n_8162), .o(n_8164) );
no02f80 g559936 ( .a(n_9080), .b(n_9079), .o(n_9081) );
no02f80 g559937 ( .a(n_8160), .b(FE_OFN967_n_9286), .o(n_8161) );
na02f80 g559938 ( .a(n_9077), .b(n_9419), .o(n_9078) );
na02f80 g559939 ( .a(n_8683), .b(n_8682), .o(n_8684) );
no02f80 g559940 ( .a(n_9075), .b(n_10553), .o(n_9076) );
no02f80 g559941 ( .a(n_7496), .b(n_3003), .o(n_10178) );
na02f80 g559942 ( .a(n_9073), .b(n_9072), .o(n_9074) );
na02f80 g559943 ( .a(n_9518), .b(n_9517), .o(n_9519) );
na02f80 g559944 ( .a(n_8158), .b(n_8157), .o(n_8159) );
no02f80 g559945 ( .a(n_8155), .b(n_8603), .o(n_8156) );
na02f80 g559946 ( .a(n_9515), .b(n_9514), .o(n_9516) );
no02f80 g559947 ( .a(n_10468), .b(FE_OFN1214_n_10469), .o(n_9071) );
in01f80 g559948 ( .a(n_15647), .o(n_9513) );
ao12f80 g559949 ( .a(n_13335), .b(n_7981), .c(n_7980), .o(n_15647) );
in01f80 g559950 ( .a(n_15285), .o(n_9512) );
ao12f80 g559951 ( .a(n_13338), .b(n_7992), .c(n_7991), .o(n_15285) );
no02f80 g559952 ( .a(n_8153), .b(n_8605), .o(n_8154) );
na02f80 g559953 ( .a(n_8151), .b(n_8599), .o(n_8152) );
oa12f80 g559954 ( .a(n_8680), .b(n_1654), .c(n_25680), .o(n_8681) );
no02f80 g559955 ( .a(n_10521), .b(FE_OFN1256_n_10520), .o(n_9070) );
na02f80 g559956 ( .a(n_10425), .b(FE_OFN658_n_10424), .o(n_9069) );
na02f80 g559957 ( .a(n_9685), .b(n_11163), .o(n_8679) );
no02f80 g559958 ( .a(n_7509), .b(n_6515), .o(n_13943) );
na02f80 g559959 ( .a(n_9510), .b(n_9509), .o(n_9511) );
na02f80 g559960 ( .a(n_9301), .b(n_8677), .o(n_8678) );
no02f80 g559961 ( .a(n_7510), .b(n_6516), .o(n_10149) );
ao22s80 g559962 ( .a(n_9396), .b(n_5658), .c(n_6340), .d(n_6339), .o(n_13453) );
no02f80 g559963 ( .a(n_7534), .b(n_2785), .o(n_14323) );
na02f80 g559964 ( .a(n_9067), .b(n_9066), .o(n_9068) );
na02f80 g559965 ( .a(n_9507), .b(n_9506), .o(n_9508) );
in01f80 g559966 ( .a(n_8150), .o(n_9366) );
oa12f80 g559967 ( .a(n_2265), .b(n_7206), .c(n_3256), .o(n_8150) );
no02f80 g559968 ( .a(n_8148), .b(n_8147), .o(n_8149) );
in01f80 g559969 ( .a(n_10153), .o(n_10152) );
ao12f80 g559970 ( .a(n_4003), .b(n_5382), .c(n_4822), .o(n_10153) );
no02f80 g559971 ( .a(n_7487), .b(n_2698), .o(n_10176) );
no02f80 g559972 ( .a(n_8799), .b(n_8145), .o(n_8146) );
na02f80 g559973 ( .a(n_8675), .b(n_8674), .o(n_8676) );
in01f80 g559974 ( .a(n_15340), .o(n_9505) );
ao12f80 g559975 ( .a(n_13344), .b(n_7996), .c(n_7995), .o(n_15340) );
na02f80 g559976 ( .a(n_8143), .b(n_8142), .o(n_8144) );
in01f80 g559977 ( .a(n_8141), .o(n_9361) );
oa12f80 g559978 ( .a(n_2171), .b(n_7205), .c(n_2813), .o(n_8141) );
na02f80 g559979 ( .a(n_8800), .b(n_8139), .o(n_8140) );
no02f80 g559980 ( .a(n_9064), .b(n_9063), .o(n_9065) );
na02f80 g559981 ( .a(n_8672), .b(n_8671), .o(n_8673) );
na02f80 g559982 ( .a(n_9503), .b(n_9502), .o(n_9504) );
no02f80 g559983 ( .a(n_7535), .b(n_2786), .o(n_10172) );
na02f80 g559984 ( .a(n_8137), .b(n_8602), .o(n_8138) );
no02f80 g559985 ( .a(n_8806), .b(n_8135), .o(n_8136) );
na02f80 g559986 ( .a(n_9663), .b(n_9662), .o(n_8670) );
in01f80 g559987 ( .a(n_11035), .o(n_11036) );
no02f80 g559988 ( .a(n_8669), .b(n_8668), .o(n_11035) );
in01f80 g559989 ( .a(n_9061), .o(n_9062) );
na02f80 g559990 ( .a(n_8669), .b(n_8668), .o(n_9061) );
in01f80 g559991 ( .a(n_15672), .o(n_11654) );
ao12f80 g559992 ( .a(n_13331), .b(n_7990), .c(n_7989), .o(n_15672) );
na02f80 g559993 ( .a(n_9500), .b(n_9499), .o(n_9501) );
na02f80 g559994 ( .a(n_9497), .b(n_9496), .o(n_9498) );
na02f80 g559995 ( .a(n_9494), .b(n_9493), .o(n_9495) );
no02f80 g559996 ( .a(n_10496), .b(FE_OFN863_n_10495), .o(n_9060) );
na02f80 g559997 ( .a(n_10493), .b(FE_OFN861_n_10492), .o(n_9059) );
no02f80 g559998 ( .a(n_10490), .b(FE_OFN1238_n_10491), .o(n_9058) );
no02f80 g559999 ( .a(n_8239), .b(n_3006), .o(n_14389) );
no02f80 g560000 ( .a(n_8240), .b(n_3007), .o(n_11083) );
na02f80 g560001 ( .a(n_9335), .b(n_9594), .o(n_8667) );
no02f80 g560002 ( .a(n_8665), .b(n_8664), .o(n_8666) );
na02f80 g560003 ( .a(n_9491), .b(n_9490), .o(n_9492) );
na02f80 g560004 ( .a(n_9488), .b(n_9487), .o(n_9489) );
no02f80 g560005 ( .a(n_8805), .b(n_8131), .o(n_8132) );
na02f80 g560006 ( .a(n_9485), .b(n_9484), .o(n_9486) );
na02f80 g560007 ( .a(n_9337), .b(n_8662), .o(n_8663) );
no02f80 g560008 ( .a(n_8209), .b(n_5144), .o(n_9057) );
no02f80 g560009 ( .a(n_9318), .b(n_8660), .o(n_8661) );
no02f80 g560010 ( .a(n_9055), .b(n_9054), .o(n_9056) );
in01f80 g560011 ( .a(n_15662), .o(n_11651) );
ao12f80 g560012 ( .a(n_13314), .b(n_7988), .c(n_7987), .o(n_15662) );
no02f80 g560013 ( .a(n_8237), .b(FE_OFN552_n_9482), .o(n_9483) );
ao22s80 g560014 ( .a(n_9053), .b(n_7210), .c(n_7429), .d(n_7430), .o(n_13456) );
no02f80 g560015 ( .a(n_10478), .b(FE_OFN554_n_9468), .o(n_9052) );
na02f80 g560016 ( .a(n_7572), .b(n_9050), .o(n_9051) );
na02f80 g560017 ( .a(n_8129), .b(n_8859), .o(n_8130) );
in01f80 g560018 ( .a(n_15641), .o(n_11648) );
ao12f80 g560019 ( .a(n_13322), .b(n_7979), .c(n_7978), .o(n_15641) );
no02f80 g560020 ( .a(n_8233), .b(n_9480), .o(n_9481) );
na02f80 g560021 ( .a(n_9478), .b(n_9477), .o(n_9479) );
na02f80 g560022 ( .a(n_10474), .b(FE_OFN552_n_9482), .o(n_9049) );
na02f80 g560023 ( .a(n_10466), .b(FE_OFN1212_n_10465), .o(n_9048) );
no02f80 g560024 ( .a(n_10463), .b(FE_OFN704_n_10462), .o(n_9047) );
no02f80 g560025 ( .a(n_10461), .b(n_9480), .o(n_9046) );
in01f80 g560026 ( .a(n_9476), .o(n_14338) );
na02f80 g560027 ( .a(n_9045), .b(n_9044), .o(n_9476) );
na02f80 g560028 ( .a(n_10449), .b(n_9042), .o(n_9043) );
in01f80 g560029 ( .a(n_11699), .o(n_14879) );
na02f80 g560030 ( .a(n_8659), .b(n_8658), .o(n_11699) );
in01f80 g560031 ( .a(n_9040), .o(n_9041) );
no02f80 g560032 ( .a(n_8659), .b(n_8658), .o(n_9040) );
no02f80 g560033 ( .a(n_10447), .b(n_9038), .o(n_9039) );
no02f80 g560034 ( .a(n_8127), .b(FE_OFN965_n_9283), .o(n_8128) );
no02f80 g560035 ( .a(n_10449), .b(FE_OFN546_n_9036), .o(n_9037) );
no02f80 g560036 ( .a(FE_OFN1220_n_8798), .b(n_8125), .o(n_8126) );
na02f80 g560037 ( .a(n_10446), .b(n_9034), .o(n_9035) );
na02f80 g560038 ( .a(n_10447), .b(n_9032), .o(n_9033) );
no02f80 g560039 ( .a(n_10446), .b(FE_OFN544_n_9030), .o(n_9031) );
in01f80 g560040 ( .a(n_15287), .o(n_11645) );
ao12f80 g560041 ( .a(n_13317), .b(n_7986), .c(n_7985), .o(n_15287) );
na02f80 g560042 ( .a(n_9474), .b(n_9473), .o(n_9475) );
na02f80 g560043 ( .a(n_9471), .b(n_9470), .o(n_9472) );
oa12f80 g560044 ( .a(n_14509), .b(n_7198), .c(n_7197), .o(n_10100) );
no02f80 g560045 ( .a(n_10368), .b(n_10367), .o(n_9029) );
na02f80 g560046 ( .a(n_10438), .b(n_10437), .o(n_9028) );
na02f80 g560047 ( .a(n_8656), .b(n_8655), .o(n_8657) );
no02f80 g560048 ( .a(n_10436), .b(n_10435), .o(n_9027) );
no02f80 g560049 ( .a(n_7506), .b(n_3004), .o(n_14332) );
no02f80 g560050 ( .a(n_9025), .b(n_9024), .o(n_9026) );
no02f80 g560051 ( .a(n_8804), .b(n_8123), .o(n_8124) );
no02f80 g560052 ( .a(n_8234), .b(FE_OFN554_n_9468), .o(n_9469) );
no02f80 g560053 ( .a(n_7507), .b(n_3005), .o(n_10170) );
in01f80 g560054 ( .a(n_8654), .o(n_10168) );
oa12f80 g560055 ( .a(n_7976), .b(n_6432), .c(n_5399), .o(n_8654) );
no02f80 g560056 ( .a(n_9623), .b(n_9622), .o(n_8653) );
ao12f80 g560057 ( .a(n_4611), .b(n_7953), .c(n_6203), .o(n_8809) );
no02f80 g560058 ( .a(n_10457), .b(FE_OFN1208_n_10456), .o(n_9023) );
no02f80 g560059 ( .a(n_8121), .b(FE_OFN963_n_9280), .o(n_8122) );
na02f80 g560060 ( .a(n_8283), .b(n_6589), .o(n_9022) );
no02f80 g560061 ( .a(n_8479), .b(n_9249), .o(n_8120) );
no02f80 g560062 ( .a(n_8260), .b(FE_OFN484_n_12038), .o(n_9467) );
no02f80 g560063 ( .a(n_8651), .b(n_8650), .o(n_8652) );
no02f80 g560064 ( .a(n_8648), .b(n_8647), .o(n_8649) );
in01f80 g560065 ( .a(n_15247), .o(n_11641) );
ao12f80 g560066 ( .a(n_13262), .b(n_7994), .c(n_7993), .o(n_15247) );
no02f80 g560067 ( .a(n_8277), .b(n_9466), .o(n_17120) );
na02f80 g560068 ( .a(n_8824), .b(n_10342), .o(n_18048) );
no02f80 g560069 ( .a(n_8279), .b(n_9465), .o(n_19021) );
oa12f80 g560070 ( .a(n_8118), .b(n_8117), .c(x_in_51_4), .o(n_8119) );
ao12f80 g560071 ( .a(n_9798), .b(n_8415), .c(n_8414), .o(n_11639) );
ao12f80 g560072 ( .a(n_11638), .b(n_8417), .c(n_8416), .o(n_11637) );
na02f80 g560073 ( .a(n_8813), .b(n_6470), .o(n_12260) );
ao12f80 g560074 ( .a(n_11636), .b(n_8413), .c(n_8412), .o(n_11635) );
ao12f80 g560075 ( .a(n_11634), .b(n_8411), .c(n_8410), .o(n_11633) );
ao12f80 g560076 ( .a(n_11632), .b(n_8409), .c(n_8408), .o(n_11631) );
ao12f80 g560077 ( .a(n_11630), .b(n_8407), .c(n_8406), .o(n_11626) );
no02f80 g560078 ( .a(n_8270), .b(n_9464), .o(n_17452) );
na02f80 g560079 ( .a(n_10411), .b(FE_OFN843_n_10412), .o(n_9021) );
no02f80 g560080 ( .a(n_10401), .b(n_10400), .o(n_9020) );
no02f80 g560081 ( .a(n_10407), .b(n_10406), .o(n_9019) );
na02f80 g560082 ( .a(n_10404), .b(n_10405), .o(n_9018) );
no02f80 g560083 ( .a(n_8262), .b(n_9016), .o(n_9017) );
na02f80 g560084 ( .a(n_9462), .b(n_9461), .o(n_9463) );
no02f80 g560085 ( .a(n_9606), .b(n_9604), .o(n_8646) );
no02f80 g560086 ( .a(n_10391), .b(n_10390), .o(n_9015) );
no02f80 g560087 ( .a(n_8115), .b(n_8114), .o(n_8116) );
na02f80 g560088 ( .a(n_9459), .b(n_9458), .o(n_9460) );
na02f80 g560089 ( .a(n_8263), .b(n_9013), .o(n_9014) );
no02f80 g560090 ( .a(n_8822), .b(FE_OFN1200_n_10340), .o(n_10341) );
no02f80 g560091 ( .a(n_9011), .b(n_9010), .o(n_9012) );
oa12f80 g560092 ( .a(n_8645), .b(n_7194), .c(n_7193), .o(n_10122) );
na02f80 g560093 ( .a(n_8643), .b(n_9582), .o(n_8644) );
no02f80 g560094 ( .a(n_9008), .b(n_9007), .o(n_9009) );
no02f80 g560095 ( .a(n_8112), .b(n_8111), .o(n_8113) );
na02f80 g560096 ( .a(n_8109), .b(n_8108), .o(n_8110) );
oa12f80 g560097 ( .a(FE_OFN398_n_8616), .b(n_1277), .c(FE_OFN1174_n_4860), .o(n_8642) );
oa12f80 g560098 ( .a(n_10109), .b(n_7165), .c(n_8191), .o(n_10096) );
no02f80 g560099 ( .a(n_8801), .b(n_8106), .o(n_8107) );
no02f80 g560100 ( .a(n_9593), .b(n_9592), .o(n_8641) );
in01f80 g560101 ( .a(n_11684), .o(n_14876) );
na02f80 g560102 ( .a(n_8640), .b(n_8639), .o(n_11684) );
in01f80 g560103 ( .a(n_9005), .o(n_9006) );
no02f80 g560104 ( .a(n_8640), .b(n_8639), .o(n_9005) );
no02f80 g560105 ( .a(n_8104), .b(n_8103), .o(n_8105) );
no02f80 g560106 ( .a(n_8210), .b(n_7571), .o(n_9457) );
na02f80 g560107 ( .a(n_8637), .b(n_8636), .o(n_8638) );
in01f80 g560108 ( .a(n_8635), .o(n_10167) );
oa12f80 g560109 ( .a(n_7972), .b(n_6328), .c(n_5400), .o(n_8635) );
na02f80 g560110 ( .a(n_10459), .b(FE_OFN1210_n_10458), .o(n_9004) );
no02f80 g560111 ( .a(n_8633), .b(n_8632), .o(n_8634) );
no02f80 g560112 ( .a(n_8816), .b(n_5966), .o(n_11543) );
na02f80 g560113 ( .a(n_9002), .b(n_9001), .o(n_9003) );
no02f80 g560114 ( .a(n_8817), .b(n_5965), .o(n_12267) );
no02f80 g560115 ( .a(n_7500), .b(n_5975), .o(n_14855) );
no02f80 g560116 ( .a(n_7501), .b(n_5976), .o(n_10150) );
no02f80 g560117 ( .a(n_8101), .b(FE_OFN787_n_8855), .o(n_8102) );
oa12f80 g560118 ( .a(n_6338), .b(n_8442), .c(n_6336), .o(n_8631) );
in01f80 g560119 ( .a(n_14014), .o(n_9000) );
ao22s80 g560120 ( .a(FE_OFN787_n_8855), .b(n_5655), .c(n_6345), .d(n_6344), .o(n_14014) );
no02f80 g560121 ( .a(n_9396), .b(n_8629), .o(n_8630) );
na02f80 g560122 ( .a(n_8099), .b(n_9227), .o(n_8100) );
ao12f80 g560123 ( .a(n_7610), .b(n_6341), .c(n_6342), .o(n_13462) );
na02f80 g560124 ( .a(n_8097), .b(n_8858), .o(n_8098) );
ao12f80 g560125 ( .a(n_7609), .b(n_6449), .c(n_6450), .o(n_13459) );
no02f80 g560126 ( .a(n_8998), .b(n_9053), .o(n_8999) );
no02f80 g560127 ( .a(n_8996), .b(n_9403), .o(n_8997) );
na02f80 g560128 ( .a(n_8628), .b(n_8627), .o(n_10768) );
in01f80 g560129 ( .a(n_8994), .o(n_8995) );
no02f80 g560130 ( .a(n_8628), .b(n_8627), .o(n_8994) );
na02f80 g560131 ( .a(n_8095), .b(n_9225), .o(n_8096) );
no02f80 g560132 ( .a(n_8992), .b(n_8991), .o(n_8993) );
na02f80 g560133 ( .a(n_8989), .b(n_8988), .o(n_8990) );
na02f80 g560134 ( .a(n_8214), .b(n_5972), .o(n_13874) );
na02f80 g560135 ( .a(n_8986), .b(FE_OFN1089_n_8985), .o(n_8987) );
na02f80 g560136 ( .a(n_8215), .b(n_5973), .o(n_11691) );
na02f80 g560137 ( .a(n_8983), .b(n_8982), .o(n_8984) );
na02f80 g560138 ( .a(n_7568), .b(n_8980), .o(n_8981) );
na02f80 g560139 ( .a(n_8978), .b(FE_OFN1274_n_8977), .o(n_8979) );
na02f80 g560140 ( .a(n_8625), .b(n_8624), .o(n_8626) );
na02f80 g560141 ( .a(n_8093), .b(n_8092), .o(n_8094) );
na02f80 g560142 ( .a(n_8622), .b(FE_OFN1091_n_8621), .o(n_8623) );
na02f80 g560143 ( .a(n_8975), .b(FE_OFN1087_n_8974), .o(n_8976) );
na02f80 g560144 ( .a(n_8972), .b(n_8971), .o(n_8973) );
na02f80 g560145 ( .a(n_8090), .b(n_8089), .o(n_8091) );
na02f80 g560146 ( .a(n_9455), .b(n_9454), .o(n_9456) );
no02f80 g560147 ( .a(n_8087), .b(n_8086), .o(n_8088) );
na02f80 g560148 ( .a(n_8619), .b(n_8618), .o(n_8620) );
oa12f80 g560149 ( .a(FE_OFN398_n_8616), .b(n_1046), .c(FE_OFN1174_n_4860), .o(n_8617) );
in01f80 g560150 ( .a(n_8969), .o(n_8970) );
no02f80 g560151 ( .a(n_8615), .b(n_8614), .o(n_8969) );
na02f80 g560152 ( .a(n_9452), .b(n_9451), .o(n_9453) );
ao22s80 g560153 ( .a(n_8613), .b(n_4778), .c(n_8612), .d(n_10970), .o(n_11430) );
na03f80 g560154 ( .a(n_6538), .b(n_10050), .c(n_8484), .o(n_9450) );
ao12f80 g560155 ( .a(n_8610), .b(n_8609), .c(n_8608), .o(n_8611) );
ao22s80 g560156 ( .a(n_6298), .b(FE_OFN1181_rst), .c(x_out_44_19), .d(FE_OFN279_n_16656), .o(n_8607) );
ao22s80 g560157 ( .a(n_7219), .b(FE_OFN1111_rst), .c(x_out_37_19), .d(n_16656), .o(n_8968) );
oa12f80 g560158 ( .a(n_8084), .b(n_8083), .c(x_in_51_6), .o(n_8085) );
oa12f80 g560159 ( .a(n_6343), .b(n_8185), .c(x_in_33_5), .o(n_8082) );
oa12f80 g560160 ( .a(n_6680), .b(n_8742), .c(x_in_33_11), .o(n_8606) );
oa12f80 g560161 ( .a(n_6352), .b(n_8173), .c(x_in_33_6), .o(n_8081) );
ao22s80 g560162 ( .a(n_8605), .b(n_5696), .c(n_6388), .d(n_7734), .o(n_13435) );
ao12f80 g560163 ( .a(n_10111), .b(n_7123), .c(n_7122), .o(n_10082) );
ao12f80 g560164 ( .a(n_10113), .b(n_7117), .c(n_7116), .o(n_10112) );
ao12f80 g560165 ( .a(n_10117), .b(n_7121), .c(n_7120), .o(n_10116) );
ao12f80 g560166 ( .a(n_10115), .b(n_7119), .c(n_7118), .o(n_10114) );
oa12f80 g560167 ( .a(n_6348), .b(n_8966), .c(x_in_33_9), .o(n_8967) );
ao12f80 g560168 ( .a(n_10119), .b(n_7107), .c(n_7106), .o(n_10118) );
oa12f80 g560169 ( .a(n_6347), .b(n_8179), .c(x_in_33_8), .o(n_8080) );
oa12f80 g560170 ( .a(n_6346), .b(n_8176), .c(x_in_33_7), .o(n_8079) );
in01f80 g560171 ( .a(n_9365), .o(n_8604) );
oa12f80 g560172 ( .a(n_6647), .b(n_8394), .c(n_4963), .o(n_9365) );
ao22s80 g560173 ( .a(n_8603), .b(n_5634), .c(n_6379), .d(n_2388), .o(n_13421) );
oa12f80 g560174 ( .a(n_6349), .b(n_8182), .c(x_in_33_10), .o(n_8078) );
in01f80 g560175 ( .a(n_11657), .o(n_10339) );
ao12f80 g560176 ( .a(n_14466), .b(n_8368), .c(n_8367), .o(n_11657) );
oa12f80 g560177 ( .a(n_7201), .b(n_8750), .c(x_in_33_4), .o(n_8077) );
ao12f80 g560178 ( .a(n_9449), .b(n_8366), .c(n_8365), .o(n_11623) );
oa22f80 g560179 ( .a(n_8602), .b(n_4859), .c(n_6377), .d(n_6378), .o(n_13417) );
oa12f80 g560180 ( .a(n_5631), .b(n_8601), .c(n_5630), .o(n_12809) );
oa12f80 g560181 ( .a(n_5628), .b(n_8600), .c(n_5629), .o(n_13396) );
in01f80 g560182 ( .a(n_10075), .o(n_8965) );
ao12f80 g560183 ( .a(n_13243), .b(n_7196), .c(n_7195), .o(n_10075) );
na02f80 g560184 ( .a(n_7874), .b(n_10902), .o(n_8964) );
ao12f80 g560185 ( .a(n_11622), .b(n_7094), .c(n_7093), .o(n_10120) );
oa22f80 g560186 ( .a(n_8599), .b(n_4855), .c(n_6365), .d(n_8598), .o(n_13432) );
ao22s80 g560187 ( .a(n_8597), .b(n_6442), .c(n_8596), .d(n_10882), .o(n_13103) );
oa12f80 g560188 ( .a(n_8075), .b(n_8074), .c(n_10004), .o(n_8076) );
oa12f80 g560189 ( .a(n_6384), .b(n_10144), .c(n_6382), .o(n_8595) );
oa12f80 g560190 ( .a(n_8963), .b(n_7869), .c(n_12425), .o(n_12343) );
ao22s80 g560191 ( .a(n_6309), .b(n_10553), .c(n_7559), .d(n_7560), .o(n_14449) );
oa22f80 g560192 ( .a(n_8594), .b(n_3158), .c(n_3756), .d(n_3755), .o(n_13450) );
ao12f80 g560193 ( .a(n_4762), .b(n_8073), .c(n_4761), .o(n_12781) );
ao12f80 g560194 ( .a(n_9834), .b(n_8461), .c(n_8462), .o(n_8593) );
in01f80 g560195 ( .a(FE_OFN574_n_10137), .o(n_8592) );
ao22s80 g560196 ( .a(n_8072), .b(n_4104), .c(n_8071), .d(n_4405), .o(n_10137) );
in01f80 g560197 ( .a(n_10134), .o(n_8591) );
ao22s80 g560198 ( .a(FE_OFN873_n_8070), .b(n_4117), .c(n_8069), .d(n_4596), .o(n_10134) );
in01f80 g560199 ( .a(n_11029), .o(n_8590) );
ao22s80 g560200 ( .a(FE_OFN1280_n_8068), .b(n_4107), .c(n_8067), .d(n_4415), .o(n_11029) );
oa22f80 g560201 ( .a(n_9419), .b(n_6305), .c(n_7456), .d(n_7455), .o(n_14240) );
in01f80 g560202 ( .a(n_8961), .o(n_8962) );
ao12f80 g560203 ( .a(n_8589), .b(n_8588), .c(n_7043), .o(n_8961) );
ao22s80 g560204 ( .a(n_8066), .b(n_4756), .c(n_8065), .d(n_10053), .o(n_12724) );
in01f80 g560205 ( .a(n_10140), .o(n_8587) );
ao22s80 g560206 ( .a(n_8064), .b(n_3509), .c(n_8063), .d(n_4416), .o(n_10140) );
in01f80 g560207 ( .a(n_10146), .o(n_8586) );
ao22s80 g560208 ( .a(n_8062), .b(n_3699), .c(n_8061), .d(n_4424), .o(n_10146) );
in01f80 g560209 ( .a(n_11032), .o(n_8585) );
ao22s80 g560210 ( .a(FE_OFN708_n_8059), .b(n_3696), .c(n_8058), .d(n_4518), .o(n_11032) );
no02f80 g560211 ( .a(n_6969), .b(n_8471), .o(n_8584) );
ao22s80 g560212 ( .a(n_5598), .b(n_8650), .c(n_6730), .d(n_6731), .o(n_14219) );
ao22s80 g560213 ( .a(n_8055), .b(n_2104), .c(x_in_5_4), .d(x_in_5_3), .o(n_9812) );
no02f80 g560214 ( .a(n_6973), .b(n_8466), .o(n_8583) );
ao22s80 g560215 ( .a(n_4913), .b(n_8103), .c(n_6385), .d(n_6386), .o(n_13409) );
ao22s80 g560216 ( .a(n_4730), .b(n_8054), .c(n_10045), .d(n_8503), .o(n_12796) );
oa12f80 g560217 ( .a(n_7837), .b(n_7021), .c(n_7020), .o(n_10110) );
oa22f80 g560218 ( .a(n_4845), .b(n_8162), .c(n_6354), .d(n_6355), .o(n_14455) );
ao12f80 g560219 ( .a(n_7838), .b(n_8581), .c(n_9336), .o(n_8582) );
in01f80 g560220 ( .a(n_8579), .o(n_8580) );
ao22s80 g560221 ( .a(n_4713), .b(n_8053), .c(n_10036), .d(n_8502), .o(n_8579) );
in01f80 g560222 ( .a(n_8577), .o(n_8578) );
ao22s80 g560223 ( .a(n_4174), .b(n_8052), .c(n_10033), .d(n_5246), .o(n_8577) );
no02f80 g560224 ( .a(n_6978), .b(n_8512), .o(n_8576) );
ao22s80 g560225 ( .a(n_4709), .b(n_8051), .c(n_10030), .d(n_4902), .o(n_12785) );
ao12f80 g560226 ( .a(n_6392), .b(n_6364), .c(n_6363), .o(n_14262) );
in01f80 g560227 ( .a(n_8574), .o(n_8575) );
ao22s80 g560228 ( .a(n_4704), .b(n_8050), .c(n_10024), .d(n_5239), .o(n_8574) );
ao22s80 g560229 ( .a(n_8573), .b(n_3660), .c(n_4401), .d(n_8539), .o(n_13934) );
oa12f80 g560230 ( .a(n_8261), .b(n_7555), .c(n_7554), .o(n_14396) );
in01f80 g560231 ( .a(n_8571), .o(n_8572) );
ao22s80 g560232 ( .a(n_4705), .b(n_8049), .c(n_10027), .d(n_10222), .o(n_8571) );
oa22f80 g560233 ( .a(n_3552), .b(n_8048), .c(n_2863), .d(n_8047), .o(n_12722) );
in01f80 g560234 ( .a(n_8959), .o(n_8960) );
oa22f80 g560235 ( .a(n_8570), .b(n_4978), .c(n_8569), .d(n_5730), .o(n_8959) );
oa22f80 g560236 ( .a(n_5182), .b(n_8046), .c(n_3061), .d(n_11166), .o(n_12794) );
in01f80 g560237 ( .a(n_8567), .o(n_8568) );
ao22s80 g560238 ( .a(n_4359), .b(n_8045), .c(n_10010), .d(n_8044), .o(n_8567) );
na02f80 g560239 ( .a(n_6983), .b(n_8499), .o(n_8566) );
oa22f80 g560240 ( .a(n_3958), .b(n_8043), .c(n_3058), .d(n_8042), .o(n_12720) );
ao22s80 g560241 ( .a(n_5573), .b(n_8041), .c(n_6717), .d(n_6716), .o(n_13414) );
oa12f80 g560242 ( .a(n_9929), .b(n_8039), .c(x_in_59_11), .o(n_8040) );
ao22s80 g560243 ( .a(n_8565), .b(n_4164), .c(n_10817), .d(n_8564), .o(n_13144) );
oa12f80 g560244 ( .a(n_8562), .b(n_9718), .c(n_8561), .o(n_8563) );
in01f80 g560245 ( .a(n_8559), .o(n_8560) );
ao22s80 g560246 ( .a(n_4290), .b(n_8037), .c(n_10001), .d(n_8036), .o(n_8559) );
oa22f80 g560247 ( .a(n_8558), .b(n_1984), .c(n_8557), .d(n_6781), .o(n_10620) );
ao12f80 g560248 ( .a(n_6474), .b(n_8440), .c(n_6472), .o(n_8556) );
in01f80 g560249 ( .a(n_8554), .o(n_8555) );
ao22s80 g560250 ( .a(n_4689), .b(n_8035), .c(n_9995), .d(n_8034), .o(n_8554) );
oa12f80 g560251 ( .a(n_7586), .b(n_5823), .c(n_8957), .o(n_8958) );
no03m80 g560252 ( .a(n_7914), .b(n_5984), .c(n_8032), .o(n_8033) );
in01f80 g560253 ( .a(n_8552), .o(n_8553) );
ao22s80 g560254 ( .a(n_4686), .b(n_8031), .c(n_9992), .d(n_2775), .o(n_8552) );
in01f80 g560255 ( .a(n_8550), .o(n_8551) );
ao22s80 g560256 ( .a(n_4265), .b(n_8030), .c(n_9989), .d(n_8029), .o(n_8550) );
in01f80 g560257 ( .a(n_10143), .o(n_8549) );
ao22s80 g560258 ( .a(n_8147), .b(n_5568), .c(n_6381), .d(n_3042), .o(n_10143) );
na02f80 g560259 ( .a(n_6950), .b(n_9910), .o(n_8548) );
ao22s80 g560260 ( .a(n_9403), .b(n_6669), .c(n_7453), .d(n_7454), .o(n_14237) );
oa12f80 g560261 ( .a(n_7566), .b(n_8562), .c(n_8598), .o(n_15261) );
ao12f80 g560262 ( .a(n_11625), .b(n_8401), .c(n_8400), .o(n_12237) );
oa22f80 g560263 ( .a(n_8956), .b(n_3506), .c(n_5260), .d(n_5342), .o(n_10734) );
ao12f80 g560264 ( .a(n_8562), .b(n_9718), .c(n_8546), .o(n_8547) );
na02f80 g560265 ( .a(n_7841), .b(n_10714), .o(n_8955) );
oa22f80 g560266 ( .a(n_8492), .b(n_5781), .c(n_8491), .d(n_9969), .o(n_12771) );
oa12f80 g560267 ( .a(n_9883), .b(n_8026), .c(x_in_35_11), .o(n_8027) );
ao12f80 g560268 ( .a(n_6260), .b(n_8545), .c(n_6261), .o(n_13427) );
ao22s80 g560269 ( .a(n_8025), .b(n_4670), .c(n_5307), .d(x_in_57_5), .o(n_9822) );
ao22s80 g560270 ( .a(n_8490), .b(n_5802), .c(n_8489), .d(n_3644), .o(n_12769) );
ao22s80 g560271 ( .a(n_8024), .b(n_5150), .c(n_8023), .d(n_4082), .o(n_12777) );
in01f80 g560272 ( .a(n_8543), .o(n_8544) );
ao22s80 g560273 ( .a(n_4661), .b(n_8022), .c(n_9949), .d(n_8021), .o(n_8543) );
oa22f80 g560274 ( .a(n_8493), .b(n_5800), .c(n_8494), .d(n_9946), .o(n_12775) );
oa22f80 g560275 ( .a(n_8495), .b(n_5798), .c(n_8496), .d(n_9940), .o(n_12779) );
ao22s80 g560276 ( .a(n_8542), .b(n_5181), .c(n_3360), .d(n_8541), .o(n_10718) );
oa12f80 g560277 ( .a(n_8326), .b(n_8954), .c(n_7751), .o(n_20071) );
na02f80 g560278 ( .a(n_8339), .b(n_11449), .o(n_9448) );
in01f80 g560279 ( .a(n_9446), .o(n_9447) );
ao22s80 g560280 ( .a(n_6226), .b(n_8953), .c(n_8952), .d(x_in_53_13), .o(n_9446) );
no02f80 g560281 ( .a(n_6960), .b(n_9875), .o(n_8540) );
oa12f80 g560282 ( .a(n_6794), .b(n_6751), .c(n_8539), .o(n_10678) );
ao22s80 g560283 ( .a(n_8020), .b(n_4954), .c(n_4078), .d(n_8019), .o(n_12773) );
in01f80 g560284 ( .a(n_9444), .o(n_9445) );
ao22s80 g560285 ( .a(n_7207), .b(n_8488), .c(n_9855), .d(n_10477), .o(n_9444) );
oa12f80 g560286 ( .a(n_8320), .b(n_8951), .c(n_7743), .o(n_16304) );
oa12f80 g560287 ( .a(n_8318), .b(n_8950), .c(n_7742), .o(n_19679) );
in01f80 g560288 ( .a(n_8948), .o(n_8949) );
oa12f80 g560289 ( .a(n_6786), .b(n_6719), .c(FE_OFN674_n_6720), .o(n_8948) );
in01f80 g560290 ( .a(n_8946), .o(n_8947) );
oa22f80 g560291 ( .a(n_8538), .b(n_4263), .c(n_10879), .d(n_8537), .o(n_8946) );
ao12f80 g560292 ( .a(n_6656), .b(n_6658), .c(n_8536), .o(n_11521) );
in01f80 g560293 ( .a(n_14090), .o(n_9443) );
oa12f80 g560294 ( .a(n_8945), .b(n_8944), .c(n_8932), .o(n_14090) );
ao22s80 g560295 ( .a(n_8017), .b(n_4318), .c(n_6750), .d(n_5337), .o(n_10692) );
oa12f80 g560296 ( .a(n_8307), .b(n_8943), .c(n_7720), .o(n_18354) );
no02f80 g560297 ( .a(n_6922), .b(n_9868), .o(n_8535) );
in01f80 g560299 ( .a(n_8941), .o(n_8942) );
oa22f80 g560300 ( .a(n_6212), .b(n_8478), .c(n_9840), .d(n_8477), .o(n_8941) );
in01f80 g560301 ( .a(n_8939), .o(n_8940) );
oa22f80 g560302 ( .a(n_8534), .b(n_5045), .c(n_10861), .d(n_8851), .o(n_8939) );
in01f80 g560303 ( .a(n_8937), .o(n_8938) );
ao22s80 g560304 ( .a(n_8533), .b(n_4614), .c(n_8532), .d(n_10793), .o(n_8937) );
oa12f80 g560305 ( .a(n_8293), .b(n_8936), .c(n_7686), .o(n_16590) );
in01f80 g560306 ( .a(n_8934), .o(n_8935) );
oa22f80 g560307 ( .a(n_8531), .b(n_3900), .c(n_8530), .d(n_10790), .o(n_8934) );
no02f80 g560308 ( .a(n_11440), .b(n_8298), .o(n_9442) );
oa12f80 g560309 ( .a(n_10754), .b(n_8528), .c(n_10212), .o(n_8529) );
na02f80 g560310 ( .a(n_7676), .b(n_10746), .o(n_8933) );
in01f80 g560311 ( .a(n_11055), .o(n_9441) );
ao12f80 g560312 ( .a(n_7911), .b(n_8932), .c(n_8376), .o(n_11055) );
in01f80 g560313 ( .a(n_12365), .o(n_8931) );
oa12f80 g560314 ( .a(n_7140), .b(n_7139), .c(n_7138), .o(n_12365) );
ao12f80 g560315 ( .a(n_6886), .b(n_6885), .c(n_6884), .o(n_9887) );
oa12f80 g560316 ( .a(n_7921), .b(n_7920), .c(n_7919), .o(n_10623) );
ao12f80 g560317 ( .a(n_7778), .b(n_7777), .c(n_7776), .o(n_10811) );
ao22s80 g560318 ( .a(n_7761), .b(n_8527), .c(n_8526), .d(n_7760), .o(n_9973) );
oa12f80 g560319 ( .a(n_7783), .b(n_7782), .c(n_7781), .o(n_10743) );
oa12f80 g560320 ( .a(n_8342), .b(n_8341), .c(n_8340), .o(n_11509) );
oa12f80 g560321 ( .a(n_6407), .b(n_6406), .c(n_6405), .o(n_9346) );
ao12f80 g560322 ( .a(n_8338), .b(n_8337), .c(n_8336), .o(n_11496) );
oa12f80 g560323 ( .a(n_7692), .b(n_7691), .c(n_7690), .o(n_10630) );
ao12f80 g560324 ( .a(n_6411), .b(n_6410), .c(n_6409), .o(n_9344) );
oa12f80 g560325 ( .a(n_7849), .b(n_7848), .c(n_7847), .o(n_10886) );
ao22s80 g560326 ( .a(n_8525), .b(x_in_35_11), .c(n_8026), .d(n_8524), .o(n_9884) );
ao22s80 g560327 ( .a(n_8523), .b(n_8075), .c(n_8074), .d(n_4550), .o(n_10005) );
in01f80 g560328 ( .a(n_10158), .o(n_8930) );
oa12f80 g560329 ( .a(n_6863), .b(n_8064), .c(n_6862), .o(n_10158) );
oa12f80 g560330 ( .a(n_8393), .b(n_8392), .c(n_9440), .o(n_11526) );
ao22s80 g560331 ( .a(n_7779), .b(n_8522), .c(n_8521), .d(x_in_7_4), .o(n_9864) );
ao22s80 g560332 ( .a(n_8520), .b(n_7723), .c(n_7724), .d(n_8519), .o(n_12747) );
oa12f80 g560333 ( .a(n_8012), .b(n_8011), .c(n_8010), .o(n_10634) );
ao22s80 g560334 ( .a(n_8518), .b(n_2410), .c(n_5960), .d(n_8517), .o(n_9911) );
in01f80 g560335 ( .a(n_9438), .o(n_9439) );
oa12f80 g560336 ( .a(n_7657), .b(n_7656), .c(n_7655), .o(n_9438) );
ao12f80 g560337 ( .a(n_7056), .b(n_7055), .c(n_7054), .o(n_10072) );
oa22f80 g560338 ( .a(n_6454), .b(n_12172), .c(n_6455), .d(x_in_33_6), .o(n_10776) );
ao12f80 g560339 ( .a(n_7664), .b(n_7663), .c(n_7662), .o(n_11006) );
oa12f80 g560340 ( .a(n_7149), .b(n_7148), .c(n_7147), .o(n_9988) );
ao12f80 g560341 ( .a(n_7890), .b(n_8601), .c(n_7889), .o(n_10895) );
ao22s80 g560342 ( .a(n_9437), .b(n_7434), .c(n_7400), .d(x_in_21_2), .o(n_11450) );
ao22s80 g560343 ( .a(n_7872), .b(n_8516), .c(n_8515), .d(n_4256), .o(n_10018) );
ao22s80 g560344 ( .a(n_7784), .b(x_in_27_11), .c(n_8514), .d(n_8513), .o(n_9908) );
ao12f80 g560345 ( .a(n_7098), .b(n_8512), .c(n_8511), .o(n_9919) );
oa12f80 g560346 ( .a(n_7405), .b(n_8594), .c(n_7404), .o(n_11153) );
oa12f80 g560347 ( .a(n_6968), .b(n_6967), .c(n_6966), .o(n_9957) );
oa22f80 g560348 ( .a(n_8510), .b(n_7844), .c(n_7845), .d(n_8509), .o(n_10179) );
oa12f80 g560349 ( .a(n_8296), .b(n_9436), .c(n_8295), .o(n_11441) );
ao22s80 g560350 ( .a(n_8334), .b(n_8929), .c(n_8928), .d(x_in_61_4), .o(n_10616) );
ao12f80 g560351 ( .a(n_7640), .b(n_8791), .c(n_7639), .o(n_10968) );
oa12f80 g560352 ( .a(n_7817), .b(n_7816), .c(n_7815), .o(n_10840) );
oa22f80 g560353 ( .a(FE_OFN456_n_8508), .b(n_6380), .c(n_5842), .d(x_in_3_11), .o(n_9876) );
oa22f80 g560354 ( .a(n_8507), .b(n_6963), .c(n_6964), .d(n_8506), .o(n_12712) );
oa12f80 g560355 ( .a(n_7647), .b(n_7646), .c(n_7645), .o(n_10846) );
ao12f80 g560356 ( .a(n_7699), .b(n_7698), .c(n_7697), .o(n_10901) );
ao12f80 g560357 ( .a(n_7678), .b(n_8927), .c(n_7677), .o(n_10747) );
oa12f80 g560358 ( .a(n_7382), .b(n_7381), .c(n_7380), .o(n_10824) );
ao12f80 g560359 ( .a(n_7667), .b(n_7666), .c(n_7665), .o(n_10910) );
ao12f80 g560360 ( .a(n_7792), .b(n_7791), .c(n_7790), .o(n_10788) );
oa12f80 g560361 ( .a(n_6934), .b(n_6933), .c(n_6932), .o(n_9889) );
oa22f80 g560362 ( .a(n_8926), .b(n_5079), .c(n_8356), .d(n_8925), .o(n_10870) );
oa22f80 g560363 ( .a(n_8505), .b(n_6970), .c(n_6971), .d(n_8504), .o(n_12708) );
oa12f80 g560364 ( .a(n_6799), .b(n_6798), .c(n_6797), .o(n_9953) );
ao12f80 g560365 ( .a(n_7843), .b(n_8924), .c(n_7842), .o(n_10715) );
ao12f80 g560366 ( .a(n_7685), .b(n_7684), .c(n_7683), .o(n_10647) );
ao12f80 g560367 ( .a(n_7733), .b(n_7732), .c(n_7731), .o(n_10876) );
ao12f80 g560368 ( .a(n_7164), .b(n_7163), .c(n_7162), .o(n_10106) );
ao22s80 g560369 ( .a(n_5954), .b(n_8503), .c(n_8054), .d(n_11148), .o(n_10046) );
in01f80 g560370 ( .a(n_10157), .o(n_8923) );
oa12f80 g560371 ( .a(n_6859), .b(n_8072), .c(n_6858), .o(n_10157) );
ao22s80 g560372 ( .a(n_5950), .b(n_8502), .c(n_8053), .d(n_11168), .o(n_10037) );
oa12f80 g560373 ( .a(n_7857), .b(n_7856), .c(n_7855), .o(n_10850) );
ao22s80 g560374 ( .a(n_5949), .b(n_10222), .c(n_8049), .d(n_10220), .o(n_10028) );
ao12f80 g560375 ( .a(n_6857), .b(n_8052), .c(n_6856), .o(n_10034) );
ao22s80 g560376 ( .a(n_6579), .b(n_8596), .c(n_8597), .d(n_6441), .o(n_10883) );
ao12f80 g560377 ( .a(n_6855), .b(n_8050), .c(FE_OFN971_n_6854), .o(n_10025) );
ao12f80 g560378 ( .a(n_6823), .b(n_8051), .c(FE_OFN973_n_6822), .o(n_10031) );
in01f80 g560379 ( .a(n_10156), .o(n_8922) );
oa12f80 g560380 ( .a(n_6853), .b(FE_OFN873_n_8070), .c(n_6852), .o(n_10156) );
oa22f80 g560381 ( .a(n_8022), .b(n_4660), .c(n_5947), .d(n_8021), .o(n_9950) );
oa12f80 g560382 ( .a(n_6920), .b(FE_OFN763_n_8501), .c(n_6919), .o(n_9869) );
oa12f80 g560383 ( .a(n_7085), .b(n_8500), .c(n_8499), .o(n_9927) );
in01f80 g560384 ( .a(n_10337), .o(n_10338) );
ao12f80 g560385 ( .a(n_8362), .b(n_8361), .c(n_8360), .o(n_10337) );
ao22s80 g560386 ( .a(n_8498), .b(n_8497), .c(n_6981), .d(n_9302), .o(n_9924) );
oa12f80 g560387 ( .a(n_7087), .b(n_8073), .c(n_7086), .o(n_9985) );
oa22f80 g560388 ( .a(n_5946), .b(n_8496), .c(n_8495), .d(n_5797), .o(n_9941) );
ao22s80 g560389 ( .a(n_7399), .b(n_8952), .c(n_8953), .d(n_6225), .o(n_11528) );
oa22f80 g560390 ( .a(n_8024), .b(n_5149), .c(n_5945), .d(n_8023), .o(n_9959) );
oa22f80 g560391 ( .a(n_5865), .b(n_8494), .c(n_8493), .d(n_5799), .o(n_9947) );
ao22s80 g560392 ( .a(n_8492), .b(n_5780), .c(n_5738), .d(n_8491), .o(n_9970) );
na02f80 g560393 ( .a(n_7638), .b(n_10751), .o(n_8921) );
oa22f80 g560394 ( .a(n_8490), .b(n_5801), .c(n_5944), .d(n_8489), .o(n_9962) );
oa22f80 g560395 ( .a(n_6575), .b(n_8920), .c(n_8919), .d(n_4379), .o(n_10752) );
in01f80 g560396 ( .a(n_10335), .o(n_10336) );
oa12f80 g560397 ( .a(n_8346), .b(n_8345), .c(x_in_35_1), .o(n_10335) );
ao22s80 g560398 ( .a(n_5739), .b(n_10477), .c(n_8488), .d(x_in_17_13), .o(n_9856) );
oa22f80 g560399 ( .a(n_8020), .b(n_4953), .c(n_5967), .d(n_8019), .o(n_9897) );
in01f80 g560400 ( .a(n_10334), .o(n_12282) );
ao12f80 g560401 ( .a(n_8288), .b(n_9179), .c(n_8287), .o(n_10334) );
ao12f80 g560402 ( .a(n_6851), .b(n_6850), .c(n_6849), .o(n_10950) );
in01f80 g560403 ( .a(n_9434), .o(n_9435) );
oa12f80 g560404 ( .a(n_7730), .b(n_7729), .c(n_7728), .o(n_9434) );
in01f80 g560405 ( .a(n_8917), .o(n_8918) );
ao12f80 g560406 ( .a(n_6931), .b(n_6930), .c(n_6929), .o(n_8917) );
ao12f80 g560407 ( .a(n_6871), .b(n_6870), .c(n_6869), .o(n_9981) );
oa12f80 g560408 ( .a(n_6900), .b(n_6899), .c(n_6898), .o(n_9872) );
ao12f80 g560409 ( .a(n_6848), .b(n_6847), .c(n_6846), .o(n_9936) );
in01f80 g560410 ( .a(n_8915), .o(n_8916) );
ao12f80 g560411 ( .a(n_6880), .b(n_6879), .c(n_6878), .o(n_8915) );
ao12f80 g560412 ( .a(n_6903), .b(n_6902), .c(n_6901), .o(n_9922) );
in01f80 g560413 ( .a(n_8913), .o(n_8914) );
ao12f80 g560414 ( .a(n_6874), .b(n_6873), .c(n_6872), .o(n_8913) );
ao12f80 g560415 ( .a(n_7059), .b(n_7058), .c(n_7057), .o(n_9965) );
ao12f80 g560416 ( .a(n_6845), .b(n_6844), .c(n_6843), .o(n_9904) );
oa12f80 g560417 ( .a(n_6937), .b(n_6936), .c(n_6935), .o(n_9892) );
oa12f80 g560418 ( .a(n_6891), .b(n_6890), .c(n_6889), .o(n_9820) );
ao12f80 g560419 ( .a(n_7155), .b(n_7154), .c(n_7153), .o(n_9386) );
ao12f80 g560420 ( .a(n_7756), .b(n_7755), .c(n_7754), .o(n_10857) );
in01f80 g560421 ( .a(n_10155), .o(n_8912) );
oa12f80 g560422 ( .a(n_6865), .b(FE_OFN708_n_8059), .c(n_6864), .o(n_10155) );
oa22f80 g560423 ( .a(n_8487), .b(n_6947), .c(n_6948), .d(n_8486), .o(n_12759) );
oa22f80 g560424 ( .a(n_5935), .b(n_11166), .c(n_8046), .d(n_8485), .o(n_10014) );
ao22s80 g560425 ( .a(n_5846), .b(n_8484), .c(n_5845), .d(n_4006), .o(n_11697) );
ao12f80 g560426 ( .a(n_7152), .b(n_7151), .c(n_7150), .o(n_10098) );
oa22f80 g560427 ( .a(n_8911), .b(n_5768), .c(n_6520), .d(n_8910), .o(n_22570) );
ao12f80 g560428 ( .a(n_7926), .b(n_7925), .c(n_8846), .o(n_10831) );
ao12f80 g560429 ( .a(n_7768), .b(n_7767), .c(x_in_19_11), .o(n_10813) );
ao12f80 g560430 ( .a(n_7892), .b(n_8600), .c(n_7891), .o(n_10890) );
ao12f80 g560431 ( .a(n_7834), .b(n_7833), .c(x_in_19_10), .o(n_10805) );
oa12f80 g560432 ( .a(n_7832), .b(n_7831), .c(x_in_19_9), .o(n_10740) );
ao12f80 g560433 ( .a(n_7830), .b(n_7829), .c(x_in_19_8), .o(n_10738) );
oa12f80 g560434 ( .a(n_7828), .b(n_7827), .c(x_in_19_7), .o(n_10782) );
in01f80 g560435 ( .a(n_9432), .o(n_9433) );
ao12f80 g560436 ( .a(n_7826), .b(n_7825), .c(x_in_19_6), .o(n_9432) );
in01f80 g560437 ( .a(n_9430), .o(n_9431) );
ao12f80 g560438 ( .a(n_7822), .b(n_7821), .c(x_in_19_5), .o(n_9430) );
ao12f80 g560439 ( .a(n_7789), .b(n_7788), .c(x_in_19_4), .o(n_10736) );
ao12f80 g560440 ( .a(n_6839), .b(n_6838), .c(n_6837), .o(n_10733) );
oa12f80 g560441 ( .a(n_8286), .b(n_8956), .c(n_8285), .o(n_11525) );
ao22s80 g560442 ( .a(n_6569), .b(n_8909), .c(n_8908), .d(n_8907), .o(n_10867) );
oa12f80 g560443 ( .a(n_7910), .b(n_7909), .c(x_in_1_5), .o(n_10989) );
ao22s80 g560444 ( .a(n_7383), .b(n_9429), .c(n_9428), .d(n_3221), .o(n_12442) );
ao22s80 g560445 ( .a(n_8483), .b(x_in_59_11), .c(n_8039), .d(n_8482), .o(n_9930) );
ao22s80 g560446 ( .a(n_6631), .b(n_8906), .c(n_8905), .d(n_8904), .o(n_10763) );
ao12f80 g560447 ( .a(n_7104), .b(n_7103), .c(n_7102), .o(n_8481) );
ao12f80 g560448 ( .a(n_7635), .b(n_8903), .c(n_7634), .o(n_10730) );
oa12f80 g560449 ( .a(n_7946), .b(n_7945), .c(n_7944), .o(n_10693) );
ao22s80 g560450 ( .a(n_6549), .b(n_8810), .c(n_8811), .d(n_7199), .o(n_10835) );
oa12f80 g560451 ( .a(n_7896), .b(n_8903), .c(n_7895), .o(n_10949) );
oa22f80 g560452 ( .a(n_6545), .b(n_8537), .c(n_8538), .d(x_in_29_10), .o(n_10880) );
no02f80 g560453 ( .a(n_6866), .b(n_8479), .o(n_8480) );
in01f80 g560454 ( .a(n_8902), .o(n_11676) );
oa12f80 g560455 ( .a(n_7115), .b(n_7114), .c(n_7113), .o(n_8902) );
in01f80 g560456 ( .a(n_11365), .o(n_11362) );
ao12f80 g560457 ( .a(n_7955), .b(n_7954), .c(n_7953), .o(n_11365) );
oa12f80 g560458 ( .a(n_7759), .b(n_7758), .c(n_7757), .o(n_10888) );
oa12f80 g560459 ( .a(n_7861), .b(n_7860), .c(x_in_49_1), .o(n_10921) );
oa12f80 g560460 ( .a(n_8282), .b(n_7633), .c(n_7632), .o(n_10726) );
ao12f80 g560461 ( .a(n_7631), .b(n_6836), .c(n_6835), .o(n_9847) );
oa12f80 g560462 ( .a(n_10725), .b(n_6868), .c(n_6867), .o(n_9849) );
oa12f80 g560463 ( .a(n_9848), .b(n_6834), .c(n_6833), .o(n_9859) );
ao12f80 g560464 ( .a(n_7643), .b(n_6861), .c(n_6860), .o(n_9804) );
ao12f80 g560465 ( .a(n_9803), .b(n_6793), .c(n_6792), .o(n_9845) );
ao12f80 g560466 ( .a(n_7146), .b(n_7145), .c(n_7924), .o(n_9976) );
ao12f80 g560467 ( .a(n_7023), .b(n_7022), .c(n_9975), .o(n_11047) );
oa12f80 g560468 ( .a(n_8901), .b(n_7630), .c(n_7629), .o(n_10722) );
in01f80 g560469 ( .a(n_8899), .o(n_8900) );
ao12f80 g560470 ( .a(n_7084), .b(n_7083), .c(n_7082), .o(n_8899) );
oa22f80 g560471 ( .a(n_8478), .b(n_7581), .c(n_6316), .d(n_8477), .o(n_9841) );
oa12f80 g560472 ( .a(n_7836), .b(n_8545), .c(n_7835), .o(n_10766) );
oa22f80 g560473 ( .a(n_8528), .b(n_10214), .c(n_8898), .d(n_10212), .o(n_10755) );
in01f80 g560474 ( .a(n_8897), .o(n_10984) );
oa12f80 g560475 ( .a(n_7063), .b(n_7062), .c(x_in_49_1), .o(n_8897) );
oa22f80 g560476 ( .a(n_6566), .b(n_8896), .c(n_8015), .d(n_5792), .o(n_20989) );
in01f80 g560477 ( .a(n_8895), .o(n_10690) );
ao12f80 g560478 ( .a(n_7066), .b(n_7065), .c(n_7064), .o(n_8895) );
ao12f80 g560479 ( .a(n_7177), .b(n_7176), .c(n_8476), .o(n_9901) );
ao22s80 g560480 ( .a(n_8475), .b(n_6290), .c(n_6976), .d(n_8474), .o(n_9917) );
in01f80 g560481 ( .a(n_8472), .o(n_8473) );
ao12f80 g560482 ( .a(n_6418), .b(n_6417), .c(n_6416), .o(n_8472) );
ao12f80 g560483 ( .a(n_7137), .b(n_8471), .c(FE_OFN1248_n_8470), .o(n_9899) );
ao22s80 g560484 ( .a(n_7867), .b(n_8469), .c(n_8468), .d(n_4551), .o(n_9999) );
ao12f80 g560485 ( .a(n_6413), .b(n_7206), .c(n_6412), .o(n_8008) );
ao22s80 g560486 ( .a(n_6565), .b(n_8541), .c(n_8542), .d(n_6359), .o(n_10821) );
ao22s80 g560487 ( .a(n_8084), .b(n_8467), .c(n_5259), .d(n_8083), .o(n_9915) );
ao12f80 g560488 ( .a(n_7975), .b(n_7974), .c(n_7973), .o(n_10717) );
ao12f80 g560489 ( .a(n_7158), .b(n_7157), .c(n_7156), .o(n_10108) );
oa12f80 g560490 ( .a(n_7131), .b(n_8466), .c(n_8465), .o(n_9913) );
ao22s80 g560491 ( .a(n_8464), .b(n_8118), .c(n_8117), .d(n_5266), .o(n_9894) );
ao22s80 g560492 ( .a(n_8463), .b(n_8462), .c(n_8461), .d(n_8460), .o(n_9835) );
ao22s80 g560493 ( .a(n_6514), .b(n_8564), .c(n_8565), .d(n_4163), .o(n_10818) );
in01f80 g560494 ( .a(n_8893), .o(n_8894) );
ao12f80 g560495 ( .a(n_7192), .b(n_8457), .c(n_7191), .o(n_8893) );
ao22s80 g560496 ( .a(n_5909), .b(n_8459), .c(n_8458), .d(n_5208), .o(n_9388) );
ao12f80 g560497 ( .a(n_7966), .b(n_7965), .c(n_7964), .o(n_10873) );
ao12f80 g560498 ( .a(n_8309), .b(n_9427), .c(n_9426), .o(n_16538) );
ao12f80 g560499 ( .a(n_6830), .b(n_6829), .c(n_6828), .o(n_9832) );
ao12f80 g560500 ( .a(n_8265), .b(n_9425), .c(n_9424), .o(n_18309) );
ao12f80 g560501 ( .a(n_8384), .b(n_9423), .c(n_9422), .o(n_20342) );
oa22f80 g560502 ( .a(n_8344), .b(n_8557), .c(n_7389), .d(x_in_21_4), .o(n_11616) );
in01f80 g560503 ( .a(n_9420), .o(n_9421) );
ao12f80 g560504 ( .a(n_7737), .b(n_7736), .c(n_7735), .o(n_9420) );
oa12f80 g560505 ( .a(n_8304), .b(n_9419), .c(n_8303), .o(n_11435) );
in01f80 g560506 ( .a(n_9417), .o(n_9418) );
ao12f80 g560507 ( .a(n_7871), .b(n_7870), .c(x_in_41_2), .o(n_9417) );
ao12f80 g560508 ( .a(n_6946), .b(n_8457), .c(n_6945), .o(n_10060) );
oa22f80 g560509 ( .a(n_6564), .b(n_8892), .c(n_8891), .d(n_5124), .o(n_17402) );
ao12f80 g560510 ( .a(n_7623), .b(n_8573), .c(n_7622), .o(n_11071) );
in01f80 g560511 ( .a(n_9415), .o(n_9416) );
ao12f80 g560512 ( .a(n_7963), .b(n_7962), .c(n_7961), .o(n_9415) );
ao12f80 g560513 ( .a(n_7618), .b(n_7617), .c(FE_OFN845_n_7616), .o(n_10703) );
ao12f80 g560514 ( .a(n_7621), .b(n_7620), .c(n_7619), .o(n_8890) );
ao12f80 g560515 ( .a(n_8396), .b(n_8395), .c(n_8394), .o(n_12310) );
in01f80 g560516 ( .a(n_12627), .o(n_8889) );
oa12f80 g560517 ( .a(n_6906), .b(n_6905), .c(n_6904), .o(n_12627) );
in01f80 g560518 ( .a(n_13117), .o(n_9414) );
oa12f80 g560519 ( .a(n_7949), .b(n_7948), .c(n_7947), .o(n_13117) );
ao12f80 g560520 ( .a(n_7886), .b(n_7885), .c(n_7884), .o(n_10830) );
ao12f80 g560521 ( .a(n_7161), .b(n_7160), .c(n_7159), .o(n_10102) );
in01f80 g560522 ( .a(n_11823), .o(n_10333) );
oa12f80 g560523 ( .a(n_8399), .b(n_8398), .c(n_8397), .o(n_11823) );
oa12f80 g560524 ( .a(n_7081), .b(n_7080), .c(n_7079), .o(n_9830) );
oa12f80 g560525 ( .a(n_6705), .b(n_8017), .c(n_6704), .o(n_10080) );
ao12f80 g560526 ( .a(n_7069), .b(n_7068), .c(n_7067), .o(n_9828) );
oa12f80 g560527 ( .a(n_7072), .b(n_7071), .c(n_7070), .o(n_11687) );
in01f80 g560528 ( .a(n_8887), .o(n_8888) );
oa12f80 g560529 ( .a(n_7090), .b(n_7089), .c(n_7088), .o(n_8887) );
oa12f80 g560530 ( .a(n_7800), .b(n_7799), .c(x_in_33_4), .o(n_10677) );
oa22f80 g560531 ( .a(n_6556), .b(x_in_33_5), .c(n_6557), .d(n_11297), .o(n_10688) );
in01f80 g560532 ( .a(n_8886), .o(n_10685) );
ao12f80 g560533 ( .a(n_7126), .b(n_7125), .c(n_7124), .o(n_8886) );
ao22s80 g560534 ( .a(n_6586), .b(x_in_33_7), .c(n_6585), .d(n_8885), .o(n_10774) );
oa22f80 g560535 ( .a(n_6536), .b(n_12175), .c(n_6537), .d(x_in_33_8), .o(n_10799) );
in01f80 g560536 ( .a(n_9412), .o(n_9413) );
ao22s80 g560537 ( .a(n_6552), .b(x_in_33_9), .c(n_6551), .d(n_8884), .o(n_9412) );
oa22f80 g560538 ( .a(n_6546), .b(n_12634), .c(n_6547), .d(x_in_33_10), .o(n_10786) );
in01f80 g560539 ( .a(n_8882), .o(n_8883) );
oa22f80 g560540 ( .a(n_5910), .b(x_in_33_11), .c(n_5911), .d(n_12178), .o(n_8882) );
ao22s80 g560541 ( .a(n_8881), .b(n_8454), .c(n_8455), .d(n_8880), .o(n_10680) );
oa12f80 g560542 ( .a(n_10679), .b(n_8455), .c(n_8454), .o(n_8456) );
in01f80 g560543 ( .a(n_9410), .o(n_9411) );
oa12f80 g560544 ( .a(n_7649), .b(n_8710), .c(n_7648), .o(n_9410) );
ao22s80 g560545 ( .a(n_5899), .b(n_8065), .c(n_8066), .d(n_4755), .o(n_10054) );
oa22f80 g560546 ( .a(n_5898), .b(n_8047), .c(n_8048), .d(n_3551), .o(n_10021) );
ao22s80 g560547 ( .a(n_8879), .b(n_7091), .c(n_6550), .d(n_8878), .o(n_10898) );
ao22s80 g560548 ( .a(n_5897), .b(n_8044), .c(n_8045), .d(n_4358), .o(n_10011) );
ao22s80 g560549 ( .a(n_8043), .b(n_3957), .c(n_5896), .d(n_8042), .o(n_10008) );
ao12f80 g560550 ( .a(n_7190), .b(n_7189), .c(n_8453), .o(n_10086) );
ao22s80 g560551 ( .a(n_5927), .b(n_8036), .c(n_8037), .d(n_4289), .o(n_10002) );
ao22s80 g560552 ( .a(n_5895), .b(n_8034), .c(n_8035), .d(n_4688), .o(n_9996) );
ao22s80 g560553 ( .a(n_5894), .b(n_8029), .c(n_8030), .d(n_4264), .o(n_9990) );
oa12f80 g560554 ( .a(n_6825), .b(n_8031), .c(FE_OFN676_n_6824), .o(n_9993) );
in01f80 g560555 ( .a(n_10331), .o(n_10332) );
oa22f80 g560556 ( .a(n_8840), .b(n_6554), .c(n_9409), .d(n_6555), .o(n_10331) );
ao22s80 g560557 ( .a(FE_OFN1083_n_8877), .b(n_4553), .c(n_6518), .d(n_8876), .o(n_10903) );
oa22f80 g560558 ( .a(n_8452), .b(n_7807), .c(n_7808), .d(n_8451), .o(n_10205) );
ao12f80 g560559 ( .a(n_6404), .b(n_7205), .c(n_6403), .o(n_8006) );
ao12f80 g560560 ( .a(n_6821), .b(n_8190), .c(n_6820), .o(n_9968) );
ao12f80 g560561 ( .a(n_7188), .b(n_8025), .c(n_7187), .o(n_10066) );
ao12f80 g560562 ( .a(n_6940), .b(n_6939), .c(n_6938), .o(n_9821) );
ao12f80 g560563 ( .a(n_6894), .b(n_6893), .c(n_6892), .o(n_9818) );
in01f80 g560564 ( .a(n_12313), .o(n_11580) );
ao12f80 g560565 ( .a(n_7960), .b(n_7959), .c(n_7958), .o(n_12313) );
oa12f80 g560566 ( .a(n_6819), .b(n_6818), .c(n_6817), .o(n_9851) );
ao12f80 g560567 ( .a(n_6816), .b(n_6815), .c(n_6814), .o(n_9816) );
in01f80 g560568 ( .a(n_8874), .o(n_8875) );
ao12f80 g560569 ( .a(n_6813), .b(n_6812), .c(n_6811), .o(n_8874) );
in01f80 g560570 ( .a(n_8872), .o(n_8873) );
oa12f80 g560571 ( .a(n_6883), .b(n_6882), .c(n_6881), .o(n_8872) );
oa22f80 g560572 ( .a(n_8450), .b(n_7002), .c(n_7003), .d(n_8449), .o(n_12716) );
in01f80 g560573 ( .a(n_8870), .o(n_8871) );
ao12f80 g560574 ( .a(n_6914), .b(n_6913), .c(n_6912), .o(n_8870) );
ao22s80 g560575 ( .a(n_7819), .b(x_in_11_11), .c(n_8448), .d(n_7818), .o(n_9978) );
in01f80 g560576 ( .a(n_9407), .o(n_9408) );
oa12f80 g560577 ( .a(n_7704), .b(n_7703), .c(n_7702), .o(n_9407) );
ao22s80 g560578 ( .a(n_6539), .b(n_8532), .c(n_8533), .d(n_4613), .o(n_10794) );
ao12f80 g560579 ( .a(n_7168), .b(n_7167), .c(n_7166), .o(n_10074) );
ao12f80 g560580 ( .a(n_6827), .b(n_8055), .c(n_6826), .o(n_9983) );
ao12f80 g560581 ( .a(n_7101), .b(n_7100), .c(n_7099), .o(n_8447) );
oa12f80 g560582 ( .a(n_6810), .b(n_6809), .c(n_6808), .o(n_9811) );
oa12f80 g560583 ( .a(n_6954), .b(n_6953), .c(n_6952), .o(n_9810) );
ao12f80 g560584 ( .a(n_6928), .b(n_6927), .c(n_6926), .o(n_9808) );
oa12f80 g560585 ( .a(n_6877), .b(n_6876), .c(n_6875), .o(n_9861) );
ao12f80 g560586 ( .a(n_6909), .b(n_6908), .c(n_6907), .o(n_9806) );
in01f80 g560587 ( .a(n_8868), .o(n_8869) );
oa12f80 g560588 ( .a(n_6897), .b(n_6896), .c(n_6895), .o(n_8868) );
in01f80 g560589 ( .a(n_8866), .o(n_8867) );
ao12f80 g560590 ( .a(n_6807), .b(n_6806), .c(n_6805), .o(n_8866) );
in01f80 g560591 ( .a(n_8864), .o(n_8865) );
ao12f80 g560592 ( .a(n_6804), .b(n_6803), .c(n_6802), .o(n_8864) );
in01f80 g560593 ( .a(n_8862), .o(n_8863) );
oa12f80 g560594 ( .a(n_6925), .b(n_6924), .c(n_6923), .o(n_8862) );
in01f80 g560595 ( .a(n_9405), .o(n_9406) );
ao12f80 g560596 ( .a(n_7615), .b(n_7614), .c(n_7613), .o(n_9405) );
oa12f80 g560597 ( .a(n_7709), .b(n_7708), .c(n_7707), .o(n_12314) );
oa22f80 g560598 ( .a(n_6544), .b(n_8530), .c(n_8531), .d(n_3899), .o(n_10791) );
in01f80 g560599 ( .a(n_9404), .o(n_11610) );
oa12f80 g560600 ( .a(n_7859), .b(n_7858), .c(x_in_29_1), .o(n_9404) );
oa12f80 g560601 ( .a(n_7612), .b(n_8570), .c(n_7611), .o(n_10976) );
oa12f80 g560602 ( .a(n_7773), .b(n_7772), .c(n_7771), .o(n_11106) );
oa22f80 g560603 ( .a(n_8446), .b(n_6464), .c(n_6465), .d(n_8445), .o(n_12710) );
ao22s80 g560604 ( .a(n_7786), .b(x_in_43_11), .c(n_8444), .d(n_8443), .o(n_9944) );
oa12f80 g560605 ( .a(n_7750), .b(n_7749), .c(n_7748), .o(n_10758) );
ao12f80 g560606 ( .a(n_9844), .b(n_6832), .c(n_6831), .o(n_10062) );
ao12f80 g560607 ( .a(n_6957), .b(n_6956), .c(n_6955), .o(n_9882) );
ao22s80 g560608 ( .a(n_6560), .b(n_8861), .c(n_8860), .d(n_3278), .o(n_10708) );
oa12f80 g560609 ( .a(n_7952), .b(n_7951), .c(n_7950), .o(n_10667) );
ao12f80 g560610 ( .a(n_7607), .b(n_7606), .c(n_7605), .o(n_10931) );
oa22f80 g560611 ( .a(n_8613), .b(n_4777), .c(n_6548), .d(n_8612), .o(n_10971) );
ao12f80 g560612 ( .a(n_8300), .b(n_9403), .c(n_8299), .o(n_11437) );
oa12f80 g560613 ( .a(n_7695), .b(n_7694), .c(n_7693), .o(n_10641) );
ao12f80 g560614 ( .a(n_7682), .b(n_9053), .c(n_7681), .o(n_10645) );
in01f80 g560615 ( .a(n_9401), .o(n_9402) );
oa12f80 g560616 ( .a(n_7680), .b(n_8859), .c(n_7679), .o(n_9401) );
ao12f80 g560617 ( .a(n_8268), .b(n_8267), .c(n_8266), .o(n_11429) );
in01f80 g560618 ( .a(n_9399), .o(n_9400) );
ao12f80 g560619 ( .a(n_7701), .b(n_8858), .c(n_7700), .o(n_9399) );
in01f80 g560620 ( .a(n_8856), .o(n_8857) );
ao22s80 g560621 ( .a(n_9227), .b(n_5408), .c(n_8442), .d(n_3095), .o(n_8856) );
in01f80 g560622 ( .a(n_9397), .o(n_9398) );
ao12f80 g560623 ( .a(n_7659), .b(FE_OFN787_n_8855), .c(n_7658), .o(n_9397) );
ao12f80 g560624 ( .a(n_7712), .b(n_7711), .c(n_7710), .o(n_10637) );
in01f80 g560625 ( .a(n_10329), .o(n_10330) );
ao12f80 g560626 ( .a(n_8306), .b(n_9396), .c(n_8305), .o(n_10329) );
ao22s80 g560627 ( .a(n_9226), .b(n_6766), .c(n_11103), .d(n_2632), .o(n_10893) );
ao12f80 g560628 ( .a(n_6506), .b(n_6505), .c(n_6504), .o(n_10104) );
in01f80 g560629 ( .a(n_8853), .o(n_8854) );
ao12f80 g560630 ( .a(n_6800), .b(n_9225), .c(n_8441), .o(n_8853) );
in01f80 g560631 ( .a(n_9394), .o(n_9395) );
oa12f80 g560632 ( .a(n_7528), .b(n_3866), .c(n_8441), .o(n_9394) );
in01f80 g560633 ( .a(n_10154), .o(n_8852) );
oa12f80 g560634 ( .a(n_6842), .b(FE_OFN1280_n_8068), .c(n_6841), .o(n_10154) );
ao12f80 g560635 ( .a(n_7652), .b(n_7651), .c(n_7650), .o(n_10632) );
ao12f80 g560636 ( .a(n_6986), .b(n_6985), .c(n_6984), .o(n_9905) );
ao12f80 g560637 ( .a(n_7050), .b(n_7049), .c(n_7048), .o(n_10064) );
ao12f80 g560638 ( .a(n_7604), .b(n_7603), .c(n_7602), .o(n_10852) );
ao12f80 g560639 ( .a(n_7795), .b(n_7794), .c(n_7793), .o(n_10713) );
ao12f80 g560640 ( .a(n_7671), .b(n_7670), .c(n_7669), .o(n_10906) );
oa12f80 g560641 ( .a(n_7717), .b(n_7716), .c(n_7715), .o(n_10626) );
ao12f80 g560642 ( .a(n_7689), .b(n_7688), .c(n_7687), .o(n_10628) );
ao12f80 g560643 ( .a(n_7674), .b(n_7673), .c(n_7672), .o(n_10621) );
oa22f80 g560644 ( .a(n_6559), .b(n_8851), .c(n_8534), .d(x_in_39_10), .o(n_10862) );
oa12f80 g560645 ( .a(n_7642), .b(n_8558), .c(n_7641), .o(n_10848) );
ao12f80 g560646 ( .a(n_8844), .b(n_8843), .c(n_8842), .o(n_10328) );
oa22f80 g560647 ( .a(n_9602), .b(n_3044), .c(n_8440), .d(n_6773), .o(n_9801) );
na02f80 g560648 ( .a(n_6840), .b(n_8643), .o(n_8439) );
oa12f80 g560649 ( .a(n_7075), .b(n_7074), .c(n_7073), .o(n_9826) );
ao12f80 g560650 ( .a(n_7143), .b(n_7142), .c(n_7141), .o(n_9954) );
in01f80 g560651 ( .a(n_11052), .o(n_9393) );
ao12f80 g560652 ( .a(n_7814), .b(n_8536), .c(n_7813), .o(n_11052) );
ao12f80 g560653 ( .a(n_7078), .b(n_7077), .c(n_7076), .o(n_10092) );
in01f80 g560654 ( .a(n_10159), .o(n_8850) );
oa12f80 g560655 ( .a(n_6791), .b(n_8062), .c(n_6790), .o(n_10159) );
oa12f80 g560656 ( .a(n_7608), .b(n_8768), .c(n_8569), .o(n_10778) );
ao12f80 g560657 ( .a(n_7053), .b(n_7052), .c(n_7051), .o(n_10070) );
ao22s80 g560658 ( .a(n_8849), .b(n_7879), .c(n_7880), .d(n_8848), .o(n_12706) );
oa22f80 g560659 ( .a(n_5262), .b(FE_OFN308_n_3069), .c(n_293), .d(FE_OFN91_n_27449), .o(n_8004) );
ao22s80 g560660 ( .a(n_6999), .b(n_8438), .c(n_8536), .d(x_in_28_1), .o(n_10039) );
oa22f80 g560661 ( .a(n_5258), .b(FE_OFN294_n_3069), .c(n_1064), .d(FE_OFN21_n_27452), .o(n_8003) );
ao22s80 g560662 ( .a(n_8932), .b(n_8847), .c(n_8377), .d(x_in_38_1), .o(n_10907) );
oa22f80 g560663 ( .a(n_7457), .b(n_26454), .c(n_34), .d(FE_OFN1111_rst), .o(n_8001) );
oa22f80 g560664 ( .a(n_5370), .b(FE_OFN267_n_4280), .c(n_181), .d(FE_OFN60_n_27012), .o(n_8000) );
oa22f80 g560665 ( .a(FE_OFN474_n_5257), .b(n_21988), .c(n_636), .d(FE_OFN96_n_27449), .o(n_7999) );
oa22f80 g560666 ( .a(n_5323), .b(FE_OFN295_n_3069), .c(n_1392), .d(FE_OFN127_n_27449), .o(n_7998) );
ao22s80 g560667 ( .a(n_8436), .b(n_3349), .c(x_out_59_23), .d(n_16893), .o(n_8437) );
ao22s80 g560668 ( .a(n_8434), .b(n_2860), .c(x_out_58_23), .d(FE_OFN280_n_16656), .o(n_8435) );
ao22s80 g560669 ( .a(n_8432), .b(n_4202), .c(x_out_60_23), .d(n_27400), .o(n_8433) );
ao22s80 g560670 ( .a(n_8430), .b(n_4296), .c(x_out_61_23), .d(FE_OFN306_n_3069), .o(n_8431) );
ao22s80 g560671 ( .a(n_8428), .b(n_4212), .c(x_out_62_23), .d(n_16028), .o(n_8429) );
ao22s80 g560672 ( .a(n_8426), .b(n_2797), .c(x_out_63_23), .d(FE_OFN274_n_16893), .o(n_8427) );
oa22f80 g560673 ( .a(n_8842), .b(n_4162), .c(n_910), .d(FE_OFN129_n_27449), .o(n_7997) );
oa22f80 g560674 ( .a(n_8421), .b(n_6959), .c(n_8425), .d(n_6958), .o(n_9838) );
oa22f80 g560675 ( .a(n_7105), .b(n_6000), .c(n_6280), .d(x_in_5_9), .o(n_10093) );
ao22s80 g560676 ( .a(n_5744), .b(x_in_43_9), .c(n_7095), .d(n_7268), .o(n_8424) );
ao22s80 g560677 ( .a(n_6281), .b(x_in_27_8), .c(n_7112), .d(n_7287), .o(n_8423) );
ao12f80 g560678 ( .a(n_7864), .b(n_8846), .c(x_in_19_12), .o(n_13260) );
ao22s80 g560679 ( .a(n_6306), .b(x_in_7_7), .c(n_6511), .d(n_6494), .o(n_8422) );
ao22s80 g560680 ( .a(n_7426), .b(x_in_39_7), .c(n_8391), .d(n_7325), .o(n_9392) );
ao22s80 g560681 ( .a(n_8845), .b(n_8497), .c(n_7930), .d(n_9302), .o(n_12791) );
oa22f80 g560682 ( .a(n_8421), .b(n_8420), .c(n_8425), .d(x_in_51_11), .o(n_9879) );
ao22s80 g560683 ( .a(n_8909), .b(x_in_19_11), .c(n_8907), .d(n_7765), .o(n_9938) );
no02f80 g560702 ( .a(n_7996), .b(n_7995), .o(n_13344) );
no02f80 g560703 ( .a(n_9180), .b(x_in_28_2), .o(n_9566) );
no02f80 g560704 ( .a(n_7994), .b(n_7993), .o(n_13262) );
no02f80 g560705 ( .a(n_7992), .b(n_7991), .o(n_13338) );
in01f80 g560706 ( .a(n_8418), .o(n_8419) );
na02f80 g560707 ( .a(n_9180), .b(x_in_28_2), .o(n_8418) );
no02f80 g560708 ( .a(n_7990), .b(n_7989), .o(n_13331) );
no02f80 g560709 ( .a(n_7988), .b(n_7987), .o(n_13314) );
no02f80 g560710 ( .a(n_7986), .b(n_7985), .o(n_13317) );
no02f80 g560711 ( .a(n_6417), .b(n_5970), .o(n_13308) );
na02f80 g560712 ( .a(n_7983), .b(n_7982), .o(n_7984) );
in01f80 g560713 ( .a(n_9149), .o(n_15228) );
no02f80 g560714 ( .a(n_7983), .b(n_7982), .o(n_9149) );
no02f80 g560715 ( .a(n_8417), .b(n_8416), .o(n_11638) );
no02f80 g560716 ( .a(n_8415), .b(n_8414), .o(n_9798) );
no02f80 g560717 ( .a(n_8413), .b(n_8412), .o(n_11636) );
no02f80 g560718 ( .a(n_8411), .b(n_8410), .o(n_11634) );
no02f80 g560719 ( .a(n_8409), .b(n_8408), .o(n_11632) );
no02f80 g560720 ( .a(n_8407), .b(n_8406), .o(n_11630) );
na02f80 g560721 ( .a(n_7866), .b(n_7865), .o(n_9562) );
in01f80 g560722 ( .a(n_8404), .o(n_8405) );
no02f80 g560723 ( .a(n_7866), .b(n_7865), .o(n_8404) );
no02f80 g560724 ( .a(n_7981), .b(n_7980), .o(n_13335) );
na02f80 g560725 ( .a(n_7199), .b(n_5311), .o(n_7200) );
na02f80 g560726 ( .a(n_7220), .b(n_8842), .o(n_10973) );
no02f80 g560727 ( .a(n_7979), .b(n_7978), .o(n_13322) );
na02f80 g560728 ( .a(n_7198), .b(n_7197), .o(n_14509) );
na03f80 g560729 ( .a(n_5222), .b(n_13251), .c(n_16909), .o(n_8680) );
no02f80 g560730 ( .a(n_7196), .b(n_7195), .o(n_13243) );
in01f80 g560731 ( .a(n_8794), .o(n_7977) );
na02f80 g560732 ( .a(n_5857), .b(n_7947), .o(n_8794) );
in01f80 g560733 ( .a(n_8402), .o(n_8403) );
no02f80 g560734 ( .a(n_7967), .b(x_in_0_3), .o(n_8402) );
na02f80 g560735 ( .a(n_7976), .b(n_6433), .o(n_9102) );
no02f80 g560736 ( .a(n_7974), .b(n_7973), .o(n_7975) );
na02f80 g560737 ( .a(n_6329), .b(n_7972), .o(n_9099) );
na02f80 g560738 ( .a(n_7970), .b(n_11367), .o(n_7971) );
na02f80 g560739 ( .a(n_7968), .b(n_10316), .o(n_7969) );
no02f80 g560740 ( .a(n_6417), .b(n_6416), .o(n_6418) );
no02f80 g560741 ( .a(n_8401), .b(n_8400), .o(n_11625) );
na02f80 g560742 ( .a(n_7967), .b(x_in_0_3), .o(n_9563) );
no02f80 g560743 ( .a(n_7965), .b(n_7964), .o(n_7966) );
na02f80 g560744 ( .a(n_7194), .b(n_7193), .o(n_8645) );
no02f80 g560745 ( .a(n_7962), .b(n_7961), .o(n_7963) );
no02f80 g560746 ( .a(n_8457), .b(n_7191), .o(n_7192) );
na02f80 g560747 ( .a(n_8398), .b(n_8397), .o(n_8399) );
no02f80 g560748 ( .a(n_7189), .b(n_8453), .o(n_7190) );
na03f80 g560749 ( .a(n_5220), .b(n_13246), .c(FE_OFN422_n_16909), .o(n_8616) );
no02f80 g560750 ( .a(n_7959), .b(n_7958), .o(n_7960) );
no02f80 g560751 ( .a(n_8025), .b(n_7187), .o(n_7188) );
in01f80 g560752 ( .a(n_7956), .o(n_7957) );
no02f80 g560753 ( .a(n_7186), .b(x_in_4_3), .o(n_7956) );
no02f80 g560754 ( .a(n_7954), .b(n_7953), .o(n_7955) );
na02f80 g560755 ( .a(n_7186), .b(x_in_4_3), .o(n_9200) );
na02f80 g560756 ( .a(n_7951), .b(n_7950), .o(n_7952) );
no02f80 g560757 ( .a(n_8843), .b(n_8842), .o(n_8844) );
na02f80 g560758 ( .a(n_7948), .b(n_7947), .o(n_7949) );
no02f80 g560759 ( .a(n_7184), .b(n_6327), .o(n_7185) );
no02f80 g560760 ( .a(n_7182), .b(n_6436), .o(n_7183) );
no02f80 g560761 ( .a(n_7180), .b(n_6322), .o(n_7181) );
na02f80 g560762 ( .a(n_7945), .b(n_7944), .o(n_7946) );
no02f80 g560763 ( .a(n_6321), .b(x_in_1_5), .o(n_8795) );
no02f80 g560764 ( .a(n_7178), .b(n_5921), .o(n_7179) );
no02f80 g560765 ( .a(n_6502), .b(n_6320), .o(n_6503) );
no02f80 g560766 ( .a(n_8395), .b(n_8394), .o(n_8396) );
na02f80 g560767 ( .a(n_5233), .b(n_10085), .o(n_5782) );
no02f80 g560768 ( .a(n_7176), .b(n_8476), .o(n_7177) );
na02f80 g560769 ( .a(n_7942), .b(n_7941), .o(n_9206) );
no02f80 g560770 ( .a(n_7942), .b(n_7941), .o(n_7943) );
in01f80 g560771 ( .a(n_13719), .o(n_7940) );
no02f80 g560772 ( .a(n_5438), .b(n_4824), .o(n_13719) );
no02f80 g560773 ( .a(n_8840), .b(x_in_45_12), .o(n_8841) );
na02f80 g560774 ( .a(n_5875), .b(n_6333), .o(n_7939) );
na02f80 g560775 ( .a(n_8392), .b(n_9440), .o(n_8393) );
no02f80 g560776 ( .a(n_7175), .b(n_7174), .o(n_9138) );
in01f80 g560777 ( .a(n_7937), .o(n_7938) );
na02f80 g560778 ( .a(n_7175), .b(n_7174), .o(n_7937) );
in01f80 g560779 ( .a(n_7935), .o(n_7936) );
no02f80 g560780 ( .a(n_7173), .b(n_7172), .o(n_7935) );
na02f80 g560781 ( .a(n_7173), .b(n_7172), .o(n_9190) );
no02f80 g560782 ( .a(n_8391), .b(x_in_39_7), .o(n_9567) );
na02f80 g560783 ( .a(n_7171), .b(n_7170), .o(n_21415) );
in01f80 g560784 ( .a(n_8785), .o(n_7934) );
no02f80 g560785 ( .a(n_7171), .b(n_7170), .o(n_8785) );
na02f80 g560786 ( .a(n_5255), .b(n_8562), .o(n_13347) );
na02f80 g560787 ( .a(n_9428), .b(n_9429), .o(n_8390) );
na02f80 g560788 ( .a(n_7933), .b(n_7932), .o(n_9559) );
in01f80 g560789 ( .a(n_8388), .o(n_8389) );
no02f80 g560790 ( .a(n_7933), .b(n_7932), .o(n_8388) );
na02f80 g560791 ( .a(n_7930), .b(n_8497), .o(n_7931) );
ao12f80 g560792 ( .a(n_8387), .b(n_4773), .c(x_in_17_1), .o(n_16002) );
in01f80 g560793 ( .a(n_15638), .o(n_8386) );
na02f80 g560794 ( .a(n_7929), .b(n_4829), .o(n_15638) );
in01f80 g560795 ( .a(n_8839), .o(n_15184) );
ao12f80 g560796 ( .a(n_8385), .b(n_3990), .c(x_in_3_1), .o(n_8839) );
in01f80 g560797 ( .a(n_9603), .o(n_7928) );
na02f80 g560798 ( .a(n_5441), .b(n_3143), .o(n_9603) );
in01f80 g560799 ( .a(n_15007), .o(n_7927) );
oa12f80 g560800 ( .a(n_7169), .b(n_4019), .c(x_in_49_2), .o(n_15007) );
no02f80 g560801 ( .a(n_7167), .b(n_7166), .o(n_7168) );
na02f80 g560802 ( .a(n_7165), .b(n_8191), .o(n_10109) );
no02f80 g560803 ( .a(n_6505), .b(n_6504), .o(n_6506) );
no02f80 g560804 ( .a(n_7163), .b(n_7162), .o(n_7164) );
no02f80 g560805 ( .a(n_7160), .b(n_7159), .o(n_7161) );
no02f80 g560806 ( .a(n_7157), .b(n_7156), .o(n_7158) );
no02f80 g560807 ( .a(n_7154), .b(n_7153), .o(n_7155) );
no02f80 g560808 ( .a(n_7151), .b(n_7150), .o(n_7152) );
na02f80 g560809 ( .a(n_7148), .b(n_7147), .o(n_7149) );
no02f80 g560810 ( .a(n_7925), .b(n_8846), .o(n_7926) );
no02f80 g560811 ( .a(n_7145), .b(n_7924), .o(n_7146) );
no02f80 g560812 ( .a(n_5917), .b(n_7924), .o(n_10061) );
no02f80 g560813 ( .a(n_9423), .b(n_9422), .o(n_8384) );
in01f80 g560814 ( .a(n_7922), .o(n_7923) );
na02f80 g560815 ( .a(n_6510), .b(n_6509), .o(n_7922) );
no02f80 g560816 ( .a(n_6510), .b(n_6509), .o(n_9174) );
oa22f80 g560817 ( .a(n_4322), .b(FE_OFN1188_n_5249), .c(n_3557), .d(n_7144), .o(n_13722) );
na02f80 g560818 ( .a(n_7920), .b(n_7919), .o(n_7921) );
oa12f80 g560819 ( .a(n_6527), .b(n_5175), .c(FE_OFN306_n_3069), .o(n_8383) );
oa12f80 g560820 ( .a(n_6523), .b(n_5172), .c(FE_OFN235_n_4162), .o(n_8382) );
oa12f80 g560821 ( .a(FE_OFN1149_n_6525), .b(n_5174), .c(n_22019), .o(n_8381) );
oa12f80 g560822 ( .a(n_6531), .b(n_5173), .c(FE_OFN404_n_28303), .o(n_8380) );
oa12f80 g560823 ( .a(FE_OFN82_n_6529), .b(n_5055), .c(n_29033), .o(n_8208) );
oa12f80 g560824 ( .a(n_4922), .b(n_5038), .c(FE_OFN405_n_28303), .o(n_7373) );
no02f80 g560825 ( .a(n_6511), .b(x_in_7_7), .o(n_8783) );
na02f80 g560826 ( .a(n_7918), .b(n_7917), .o(n_9553) );
in01f80 g560827 ( .a(n_8378), .o(n_8379) );
no02f80 g560828 ( .a(n_7918), .b(n_7917), .o(n_8378) );
no02f80 g560829 ( .a(n_7142), .b(n_7141), .o(n_7143) );
na02f80 g560830 ( .a(n_7139), .b(n_7138), .o(n_7140) );
no02f80 g560831 ( .a(n_6004), .b(n_7915), .o(n_7916) );
na02f80 g560832 ( .a(n_5985), .b(n_7914), .o(n_9708) );
no02f80 g560833 ( .a(n_8471), .b(FE_OFN1248_n_8470), .o(n_7137) );
no02f80 g560834 ( .a(n_7135), .b(n_11346), .o(n_7136) );
in01f80 g560835 ( .a(n_7912), .o(n_7913) );
no02f80 g560836 ( .a(n_7133), .b(n_7134), .o(n_7912) );
no02f80 g560837 ( .a(n_8932), .b(n_8376), .o(n_7911) );
na02f80 g560838 ( .a(n_7909), .b(x_in_1_5), .o(n_7910) );
no02f80 g560839 ( .a(n_8377), .b(n_8376), .o(n_12288) );
na02f80 g560840 ( .a(n_7133), .b(n_7134), .o(n_9166) );
in01f80 g560841 ( .a(n_8374), .o(n_8375) );
no02f80 g560842 ( .a(n_7908), .b(n_7907), .o(n_8374) );
na02f80 g560843 ( .a(n_7908), .b(n_7907), .o(n_9552) );
na02f80 g560844 ( .a(n_8434), .b(n_7906), .o(n_9155) );
na02f80 g560845 ( .a(n_8436), .b(n_7905), .o(n_9152) );
na02f80 g560846 ( .a(n_8432), .b(n_7904), .o(n_9153) );
na02f80 g560847 ( .a(n_8426), .b(n_7903), .o(n_9154) );
na02f80 g560848 ( .a(n_8428), .b(n_7902), .o(n_9150) );
na02f80 g560849 ( .a(n_8430), .b(n_7901), .o(n_9151) );
no02f80 g560850 ( .a(n_7176), .b(x_in_51_9), .o(n_7132) );
na02f80 g560851 ( .a(n_8466), .b(n_8465), .o(n_7131) );
na02f80 g560852 ( .a(n_7130), .b(n_7129), .o(n_9797) );
in01f80 g560853 ( .a(n_9387), .o(n_9796) );
no02f80 g560854 ( .a(n_7130), .b(n_7129), .o(n_9387) );
oa12f80 g560855 ( .a(n_6533), .b(n_5198), .c(n_27681), .o(n_8373) );
no02f80 g560856 ( .a(n_7127), .b(n_6284), .o(n_7128) );
in01f80 g560857 ( .a(n_9390), .o(n_9391) );
no02f80 g560858 ( .a(n_8838), .b(n_8837), .o(n_9390) );
no02f80 g560859 ( .a(n_7899), .b(n_5731), .o(n_7900) );
na02f80 g560860 ( .a(n_8838), .b(n_8837), .o(n_11381) );
in01f80 g560861 ( .a(n_7897), .o(n_7898) );
oa12f80 g560862 ( .a(n_5396), .b(n_4715), .c(n_10477), .o(n_7897) );
na02f80 g560863 ( .a(n_8903), .b(n_7895), .o(n_7896) );
in01f80 g560864 ( .a(n_8371), .o(n_8372) );
no02f80 g560865 ( .a(n_7894), .b(n_7893), .o(n_8371) );
na02f80 g560866 ( .a(n_7894), .b(n_7893), .o(n_9545) );
no02f80 g560867 ( .a(n_7125), .b(n_7124), .o(n_7126) );
no02f80 g560868 ( .a(n_8600), .b(n_7891), .o(n_7892) );
no02f80 g560869 ( .a(n_7123), .b(n_7122), .o(n_10111) );
no02f80 g560870 ( .a(n_7121), .b(n_7120), .o(n_10117) );
no02f80 g560871 ( .a(n_7119), .b(n_7118), .o(n_10115) );
no02f80 g560872 ( .a(n_7117), .b(n_7116), .o(n_10113) );
na02f80 g560873 ( .a(n_7114), .b(n_7113), .o(n_7115) );
no02f80 g560874 ( .a(n_7920), .b(n_4771), .o(n_13254) );
no02f80 g560875 ( .a(n_8601), .b(n_7889), .o(n_7890) );
no02f80 g560876 ( .a(n_7112), .b(x_in_27_8), .o(n_8772) );
in01f80 g560877 ( .a(n_7110), .o(n_7111) );
no02f80 g560878 ( .a(n_6415), .b(n_6414), .o(n_7110) );
in01f80 g560879 ( .a(n_7108), .o(n_7109) );
na02f80 g560880 ( .a(n_6415), .b(n_6414), .o(n_7108) );
no02f80 g560881 ( .a(n_7107), .b(n_7106), .o(n_10119) );
na02f80 g560882 ( .a(n_7888), .b(n_7887), .o(n_9544) );
in01f80 g560883 ( .a(n_8369), .o(n_8370) );
no02f80 g560884 ( .a(n_7888), .b(n_7887), .o(n_8369) );
no02f80 g560885 ( .a(n_7105), .b(x_in_5_9), .o(n_8776) );
no02f80 g560886 ( .a(n_7885), .b(n_7884), .o(n_7886) );
no02f80 g560887 ( .a(n_7103), .b(n_7102), .o(n_7104) );
no02f80 g560888 ( .a(n_8368), .b(n_8367), .o(n_14466) );
oa12f80 g560889 ( .a(n_6040), .b(n_4712), .c(n_4017), .o(n_15186) );
no02f80 g560890 ( .a(n_7100), .b(n_7099), .o(n_7101) );
no02f80 g560891 ( .a(n_8512), .b(n_8511), .o(n_7098) );
in01f80 g560892 ( .a(n_9449), .o(n_8836) );
no02f80 g560893 ( .a(n_8366), .b(n_8365), .o(n_9449) );
in01f80 g560894 ( .a(n_7882), .o(n_7883) );
na02f80 g560895 ( .a(n_7097), .b(n_7096), .o(n_7882) );
no02f80 g560896 ( .a(n_7097), .b(n_7096), .o(n_9143) );
no02f80 g560897 ( .a(n_8392), .b(x_in_51_11), .o(n_8364) );
no02f80 g560898 ( .a(n_7095), .b(x_in_43_9), .o(n_8766) );
no02f80 g560899 ( .a(n_7094), .b(n_7093), .o(n_11622) );
na02f80 g560900 ( .a(n_7880), .b(n_7879), .o(n_7881) );
na02f80 g560901 ( .a(n_7091), .b(n_10897), .o(n_7092) );
in01f80 g560902 ( .a(n_12834), .o(n_8363) );
no02f80 g560903 ( .a(n_7878), .b(n_7877), .o(n_12834) );
na02f80 g560904 ( .a(n_7875), .b(n_2900), .o(n_7876) );
na02f80 g560905 ( .a(FE_OFN1083_n_8877), .b(n_8876), .o(n_7874) );
na02f80 g560906 ( .a(n_7872), .b(n_2922), .o(n_7873) );
na02f80 g560907 ( .a(n_5234), .b(n_4575), .o(n_8754) );
na02f80 g560908 ( .a(n_7089), .b(n_7088), .o(n_7090) );
na02f80 g560909 ( .a(n_8073), .b(n_7086), .o(n_7087) );
no02f80 g560910 ( .a(n_7206), .b(n_6412), .o(n_6413) );
na02f80 g560911 ( .a(n_8500), .b(n_8499), .o(n_7085) );
no02f80 g560912 ( .a(n_7083), .b(n_7082), .o(n_7084) );
na02f80 g560913 ( .a(n_7080), .b(n_7079), .o(n_7081) );
no02f80 g560914 ( .a(n_7870), .b(x_in_41_2), .o(n_7871) );
no02f80 g560915 ( .a(n_7077), .b(n_7076), .o(n_7078) );
no02f80 g560916 ( .a(n_8361), .b(n_8360), .o(n_8362) );
na02f80 g560917 ( .a(n_7074), .b(n_7073), .o(n_7075) );
na02f80 g560918 ( .a(n_7869), .b(n_12425), .o(n_8963) );
na02f80 g560919 ( .a(n_7867), .b(n_3312), .o(n_7868) );
na02f80 g560920 ( .a(n_7071), .b(n_7070), .o(n_7072) );
in01f80 g560921 ( .a(n_8834), .o(n_8835) );
na02f80 g560922 ( .a(n_8359), .b(n_8358), .o(n_8834) );
no02f80 g560923 ( .a(n_8359), .b(n_8358), .o(n_10345) );
no02f80 g560924 ( .a(n_7925), .b(n_2352), .o(n_7864) );
no02f80 g560925 ( .a(n_7862), .b(n_6274), .o(n_7863) );
no02f80 g560926 ( .a(n_7068), .b(n_7067), .o(n_7069) );
no02f80 g560927 ( .a(n_7065), .b(n_7064), .o(n_7066) );
na02f80 g560928 ( .a(n_7860), .b(x_in_49_1), .o(n_7861) );
na02f80 g560929 ( .a(n_7858), .b(x_in_29_1), .o(n_7859) );
na02f80 g560930 ( .a(n_7062), .b(x_in_49_1), .o(n_7063) );
no02f80 g560931 ( .a(n_7060), .b(n_6273), .o(n_7061) );
na02f80 g560932 ( .a(n_7856), .b(n_7855), .o(n_7857) );
na02f80 g560933 ( .a(n_8356), .b(n_10869), .o(n_8357) );
no02f80 g560934 ( .a(n_7058), .b(n_7057), .o(n_7059) );
no02f80 g560935 ( .a(n_7055), .b(n_7054), .o(n_7056) );
no02f80 g560936 ( .a(n_7052), .b(n_7051), .o(n_7053) );
no02f80 g560937 ( .a(n_7049), .b(n_7048), .o(n_7050) );
na02f80 g560938 ( .a(n_6663), .b(n_7904), .o(n_8355) );
na02f80 g560939 ( .a(n_6664), .b(n_7903), .o(n_8354) );
na02f80 g560940 ( .a(n_6665), .b(n_7905), .o(n_8353) );
na02f80 g560941 ( .a(n_6666), .b(n_7906), .o(n_8352) );
in01f80 g560942 ( .a(n_7853), .o(n_7854) );
no02f80 g560943 ( .a(n_7047), .b(n_9295), .o(n_7853) );
no02f80 g560944 ( .a(n_7045), .b(n_6270), .o(n_7046) );
no02f80 g560945 ( .a(n_8907), .b(n_10866), .o(n_7044) );
in01f80 g560946 ( .a(n_8589), .o(n_7852) );
no02f80 g560947 ( .a(n_8588), .b(n_7043), .o(n_8589) );
na02f80 g560948 ( .a(n_6661), .b(n_7902), .o(n_8351) );
na02f80 g560949 ( .a(n_6662), .b(n_7901), .o(n_8350) );
no02f80 g560950 ( .a(n_7041), .b(n_6160), .o(n_7042) );
no02f80 g560951 ( .a(n_7850), .b(n_6269), .o(n_7851) );
na02f80 g560952 ( .a(n_6016), .b(n_12817), .o(n_10050) );
na02f80 g560953 ( .a(n_7848), .b(n_7847), .o(n_7849) );
na02f80 g560954 ( .a(n_6623), .b(x_in_41_6), .o(n_8349) );
na02f80 g560955 ( .a(n_7845), .b(n_7844), .o(n_7846) );
no02f80 g560956 ( .a(n_8924), .b(n_7842), .o(n_7843) );
na02f80 g560957 ( .a(n_8924), .b(n_7840), .o(n_7841) );
no02f80 g560958 ( .a(n_7038), .b(n_6262), .o(n_7039) );
no02f80 g560959 ( .a(n_7036), .b(n_6267), .o(n_7037) );
na02f80 g560960 ( .a(n_5906), .b(x_in_41_9), .o(n_7035) );
na02f80 g560961 ( .a(n_5981), .b(x_in_41_7), .o(n_7034) );
na02f80 g560962 ( .a(n_6561), .b(x_in_41_11), .o(n_7839) );
no02f80 g560963 ( .a(n_7032), .b(n_6266), .o(n_7033) );
no02f80 g560964 ( .a(n_7030), .b(n_6265), .o(n_7031) );
no02f80 g560965 ( .a(n_7028), .b(n_6264), .o(n_7029) );
no02f80 g560966 ( .a(n_7026), .b(n_6263), .o(n_7027) );
no02f80 g560967 ( .a(n_7024), .b(n_6310), .o(n_7025) );
no02f80 g560968 ( .a(n_7022), .b(n_9975), .o(n_7023) );
ao12f80 g560969 ( .a(n_3063), .b(n_4731), .c(x_in_19_13), .o(n_8763) );
in01f80 g560970 ( .a(n_8347), .o(n_8348) );
na02f80 g560971 ( .a(n_8581), .b(n_7838), .o(n_8347) );
in01f80 g560972 ( .a(n_7837), .o(n_10081) );
na02f80 g560973 ( .a(n_7021), .b(n_7020), .o(n_7837) );
oa22f80 g560974 ( .a(n_4382), .b(FE_OFN1073_n_6399), .c(n_3768), .d(n_6693), .o(n_13691) );
na02f80 g560975 ( .a(n_8545), .b(n_7835), .o(n_7836) );
no02f80 g560976 ( .a(n_7384), .b(x_in_35_1), .o(n_11300) );
na02f80 g560977 ( .a(n_8345), .b(x_in_35_1), .o(n_8346) );
no02f80 g560978 ( .a(n_7833), .b(x_in_19_10), .o(n_7834) );
na02f80 g560979 ( .a(n_7831), .b(x_in_19_9), .o(n_7832) );
no02f80 g560980 ( .a(n_7829), .b(x_in_19_8), .o(n_7830) );
na02f80 g560981 ( .a(n_7827), .b(x_in_19_7), .o(n_7828) );
no02f80 g560982 ( .a(n_7825), .b(x_in_19_6), .o(n_7826) );
no02f80 g560983 ( .a(n_7017), .b(n_6256), .o(n_7018) );
no02f80 g560984 ( .a(n_7015), .b(n_6255), .o(n_7016) );
no02f80 g560985 ( .a(n_7013), .b(n_6247), .o(n_7014) );
no02f80 g560986 ( .a(n_7011), .b(n_6250), .o(n_7012) );
no02f80 g560987 ( .a(n_7009), .b(n_6251), .o(n_7010) );
no02f80 g560988 ( .a(n_7823), .b(n_6258), .o(n_7824) );
no02f80 g560989 ( .a(n_7821), .b(x_in_19_5), .o(n_7822) );
na02f80 g560990 ( .a(n_7819), .b(n_7818), .o(n_7820) );
no02f80 g560991 ( .a(n_11091), .b(x_in_41_5), .o(n_7008) );
na02f80 g560992 ( .a(n_11091), .b(x_in_41_5), .o(n_7007) );
no02f80 g560993 ( .a(n_7005), .b(n_6419), .o(n_7006) );
no02f80 g560994 ( .a(n_7003), .b(n_7002), .o(n_7004) );
no02f80 g560995 ( .a(n_7000), .b(n_6248), .o(n_7001) );
na02f80 g560996 ( .a(n_7816), .b(n_7815), .o(n_7817) );
no02f80 g560997 ( .a(n_8536), .b(n_7813), .o(n_7814) );
in01f80 g560998 ( .a(n_7812), .o(n_9181) );
na02f80 g560999 ( .a(n_6999), .b(n_7813), .o(n_7812) );
no02f80 g561000 ( .a(n_6997), .b(n_6421), .o(n_6998) );
no02f80 g561001 ( .a(n_6995), .b(n_6241), .o(n_6996) );
no02f80 g561002 ( .a(n_6993), .b(n_6242), .o(n_6994) );
no02f80 g561003 ( .a(n_6991), .b(n_6243), .o(n_6992) );
no02f80 g561004 ( .a(n_6989), .b(n_6238), .o(n_6990) );
no02f80 g561005 ( .a(n_6987), .b(n_6244), .o(n_6988) );
no02f80 g561006 ( .a(n_6985), .b(n_6984), .o(n_6986) );
no02f80 g561007 ( .a(n_6410), .b(n_6409), .o(n_6411) );
na02f80 g561008 ( .a(n_7810), .b(n_6420), .o(n_7811) );
na02f80 g561009 ( .a(n_8344), .b(x_in_21_4), .o(n_13685) );
na02f80 g561010 ( .a(n_7808), .b(n_7807), .o(n_7809) );
na02f80 g561011 ( .a(n_6019), .b(n_11040), .o(n_7806) );
na02f80 g561012 ( .a(n_6020), .b(n_11041), .o(n_7805) );
na02f80 g561013 ( .a(n_7203), .b(n_11037), .o(n_8343) );
na02f80 g561014 ( .a(n_6018), .b(n_11698), .o(n_7804) );
no02f80 g561015 ( .a(n_7802), .b(n_6233), .o(n_7803) );
na02f80 g561016 ( .a(n_6024), .b(n_11034), .o(n_7801) );
na02f80 g561017 ( .a(n_7799), .b(x_in_33_4), .o(n_7800) );
na02f80 g561018 ( .a(n_6025), .b(n_11696), .o(n_7798) );
na02f80 g561019 ( .a(n_8341), .b(n_8340), .o(n_8342) );
no02f80 g561020 ( .a(n_7796), .b(n_6257), .o(n_7797) );
no02f80 g561021 ( .a(n_7794), .b(n_7793), .o(n_7795) );
na02f80 g561022 ( .a(n_8500), .b(n_9926), .o(n_6983) );
no02f80 g561023 ( .a(n_6981), .b(n_4023), .o(n_6982) );
no02f80 g561024 ( .a(n_7791), .b(n_7790), .o(n_7792) );
no02f80 g561025 ( .a(n_7788), .b(x_in_19_4), .o(n_7789) );
no02f80 g561026 ( .a(n_6979), .b(n_6229), .o(n_6980) );
no02f80 g561027 ( .a(n_8511), .b(x_in_51_10), .o(n_6978) );
no02f80 g561028 ( .a(n_6976), .b(x_in_51_8), .o(n_6977) );
no02f80 g561029 ( .a(n_6465), .b(n_6464), .o(n_6466) );
na02f80 g561030 ( .a(n_7786), .b(n_8443), .o(n_7787) );
no02f80 g561031 ( .a(n_6974), .b(n_6228), .o(n_6975) );
no02f80 g561032 ( .a(n_8465), .b(x_in_51_5), .o(n_6973) );
no02f80 g561033 ( .a(n_6971), .b(n_6970), .o(n_6972) );
na02f80 g561034 ( .a(n_7784), .b(n_8513), .o(n_7785) );
na02f80 g561035 ( .a(n_6406), .b(n_6405), .o(n_6407) );
na02f80 g561036 ( .a(n_9437), .b(x_in_21_2), .o(n_8339) );
na02f80 g561037 ( .a(n_7782), .b(n_7781), .o(n_7783) );
no02f80 g561038 ( .a(FE_OFN1248_n_8470), .b(x_in_51_7), .o(n_6969) );
na02f80 g561039 ( .a(n_7779), .b(x_in_7_4), .o(n_7780) );
na02f80 g561040 ( .a(n_6967), .b(n_6966), .o(n_6968) );
no02f80 g561041 ( .a(n_7777), .b(n_7776), .o(n_7778) );
na02f80 g561042 ( .a(n_7774), .b(n_6275), .o(n_7775) );
no02f80 g561043 ( .a(n_6964), .b(n_6963), .o(n_6965) );
no02f80 g561044 ( .a(n_6961), .b(n_6227), .o(n_6962) );
no02f80 g561045 ( .a(FE_OFN456_n_8508), .b(x_in_3_11), .o(n_6960) );
na02f80 g561046 ( .a(n_7772), .b(n_7771), .o(n_7773) );
no02f80 g561047 ( .a(n_6956), .b(n_6955), .o(n_6957) );
no02f80 g561048 ( .a(n_8337), .b(n_8336), .o(n_8338) );
na02f80 g561049 ( .a(n_8334), .b(x_in_61_4), .o(n_8335) );
na02f80 g561050 ( .a(n_6953), .b(n_6952), .o(n_6954) );
in01f80 g561051 ( .a(n_8832), .o(n_8833) );
no02f80 g561052 ( .a(n_6568), .b(n_4933), .o(n_8832) );
no02f80 g561053 ( .a(n_6567), .b(n_4934), .o(n_9535) );
no02f80 g561054 ( .a(n_7769), .b(n_6222), .o(n_7770) );
no02f80 g561055 ( .a(n_7767), .b(x_in_19_11), .o(n_7768) );
na02f80 g561056 ( .a(n_8909), .b(n_7765), .o(n_7766) );
in01f80 g561057 ( .a(n_12167), .o(n_12169) );
na02f80 g561058 ( .a(n_7142), .b(n_2948), .o(n_12167) );
no02f80 g561059 ( .a(n_8421), .b(x_in_51_11), .o(n_6951) );
na02f80 g561060 ( .a(n_8518), .b(n_8517), .o(n_6950) );
in01f80 g561061 ( .a(n_8332), .o(n_8333) );
na02f80 g561062 ( .a(n_7764), .b(n_7763), .o(n_8332) );
no02f80 g561063 ( .a(n_7764), .b(n_7763), .o(n_9534) );
no02f80 g561064 ( .a(n_6948), .b(n_6947), .o(n_6949) );
na02f80 g561065 ( .a(n_7761), .b(n_7760), .o(n_7762) );
no02f80 g561066 ( .a(n_8457), .b(n_6945), .o(n_6946) );
na02f80 g561067 ( .a(n_7758), .b(n_7757), .o(n_7759) );
in01f80 g561068 ( .a(n_8330), .o(n_8331) );
na02f80 g561069 ( .a(n_6427), .b(n_9891), .o(n_8330) );
no02f80 g561070 ( .a(n_6426), .b(n_6943), .o(n_6944) );
no02f80 g561071 ( .a(n_7205), .b(n_6403), .o(n_6404) );
na02f80 g561072 ( .a(n_5834), .b(n_9888), .o(n_24515) );
na02f80 g561073 ( .a(n_6618), .b(n_8328), .o(n_8329) );
no02f80 g561074 ( .a(n_7755), .b(n_7754), .o(n_7756) );
no02f80 g561075 ( .a(n_5419), .b(n_2842), .o(n_12053) );
no02f80 g561076 ( .a(n_6268), .b(n_6941), .o(n_6942) );
na02f80 g561077 ( .a(n_6041), .b(n_7752), .o(n_7753) );
in01f80 g561078 ( .a(n_8326), .o(n_8327) );
na02f80 g561079 ( .a(n_8954), .b(n_7751), .o(n_8326) );
no02f80 g561080 ( .a(n_6939), .b(n_6938), .o(n_6940) );
ao12f80 g561081 ( .a(n_3022), .b(n_4219), .c(n_5938), .o(n_13228) );
na02f80 g561082 ( .a(n_7749), .b(n_7748), .o(n_7750) );
no02f80 g561083 ( .a(n_6239), .b(n_7746), .o(n_7747) );
in01f80 g561084 ( .a(n_8830), .o(n_8831) );
no02f80 g561085 ( .a(n_8325), .b(n_8324), .o(n_8830) );
na02f80 g561086 ( .a(n_8325), .b(n_8324), .o(n_10344) );
na02f80 g561087 ( .a(n_7745), .b(n_7744), .o(n_9533) );
in01f80 g561088 ( .a(n_8322), .o(n_8323) );
no02f80 g561089 ( .a(n_7745), .b(n_7744), .o(n_8322) );
na02f80 g561090 ( .a(n_6936), .b(n_6935), .o(n_6937) );
na02f80 g561091 ( .a(n_6933), .b(n_6932), .o(n_6934) );
in01f80 g561092 ( .a(n_8320), .o(n_8321) );
na02f80 g561093 ( .a(n_8951), .b(n_7743), .o(n_8320) );
in01f80 g561094 ( .a(n_8318), .o(n_8319) );
na02f80 g561095 ( .a(n_8950), .b(n_7742), .o(n_8318) );
in01f80 g561096 ( .a(n_13277), .o(n_8829) );
no02f80 g561097 ( .a(n_8317), .b(n_8316), .o(n_13277) );
no02f80 g561098 ( .a(n_7740), .b(n_10236), .o(n_7741) );
na02f80 g561099 ( .a(n_7739), .b(n_7738), .o(n_9528) );
in01f80 g561100 ( .a(n_8314), .o(n_8315) );
no02f80 g561101 ( .a(n_7739), .b(n_7738), .o(n_8314) );
no02f80 g561102 ( .a(n_6930), .b(n_6929), .o(n_6931) );
no02f80 g561103 ( .a(n_7736), .b(n_7735), .o(n_7737) );
no02f80 g561104 ( .a(n_6927), .b(n_6926), .o(n_6928) );
no02f80 g561105 ( .a(n_5955), .b(n_7734), .o(n_10234) );
no02f80 g561106 ( .a(n_7732), .b(n_7731), .o(n_7733) );
na02f80 g561107 ( .a(n_7729), .b(n_7728), .o(n_7730) );
na02f80 g561108 ( .a(n_6924), .b(n_6923), .o(n_6925) );
na02f80 g561109 ( .a(n_6650), .b(n_8312), .o(n_8313) );
in01f80 g561110 ( .a(n_8310), .o(n_8311) );
na02f80 g561111 ( .a(n_6462), .b(n_7475), .o(n_8310) );
na02f80 g561112 ( .a(n_6463), .b(n_7474), .o(n_9527) );
no02f80 g561113 ( .a(FE_OFN763_n_8501), .b(n_6921), .o(n_6922) );
na02f80 g561114 ( .a(FE_OFN763_n_8501), .b(n_6919), .o(n_6920) );
oa12f80 g561115 ( .a(n_3050), .b(n_4679), .c(n_3734), .o(n_11327) );
no02f80 g561116 ( .a(n_7726), .b(n_6649), .o(n_7727) );
oa12f80 g561117 ( .a(n_3046), .b(n_4360), .c(n_3760), .o(n_11330) );
na02f80 g561118 ( .a(n_7381), .b(n_7380), .o(n_7382) );
in01f80 g561119 ( .a(n_8827), .o(n_8828) );
no02f80 g561120 ( .a(n_6453), .b(n_5118), .o(n_8827) );
no02f80 g561121 ( .a(n_6452), .b(n_5119), .o(n_9526) );
na02f80 g561122 ( .a(n_7724), .b(n_7723), .o(n_7725) );
no02f80 g561123 ( .a(n_9427), .b(n_9426), .o(n_8309) );
no02f80 g561124 ( .a(n_6259), .b(n_6917), .o(n_6918) );
no02f80 g561125 ( .a(n_11186), .b(n_6915), .o(n_6916) );
no02f80 g561126 ( .a(n_6913), .b(n_6912), .o(n_6914) );
na02f80 g561127 ( .a(n_6236), .b(n_7721), .o(n_7722) );
in01f80 g561128 ( .a(n_8307), .o(n_8308) );
na02f80 g561129 ( .a(n_8943), .b(n_7720), .o(n_8307) );
in01f80 g561130 ( .a(n_7718), .o(n_7719) );
na02f80 g561131 ( .a(n_6911), .b(n_6910), .o(n_7718) );
no02f80 g561132 ( .a(n_6911), .b(n_6910), .o(n_9094) );
no02f80 g561133 ( .a(n_6908), .b(n_6907), .o(n_6909) );
na02f80 g561134 ( .a(n_6905), .b(n_6904), .o(n_6906) );
na02f80 g561135 ( .a(n_7716), .b(n_7715), .o(n_7717) );
na02f80 g561136 ( .a(n_6370), .b(n_7713), .o(n_7714) );
no02f80 g561137 ( .a(n_6902), .b(n_6901), .o(n_6903) );
no02f80 g561138 ( .a(n_9396), .b(n_8305), .o(n_8306) );
na02f80 g561139 ( .a(n_9419), .b(n_8303), .o(n_8304) );
na02f80 g561140 ( .a(n_6899), .b(n_6898), .o(n_6900) );
in01f80 g561141 ( .a(n_8825), .o(n_8826) );
na02f80 g561142 ( .a(n_8302), .b(n_8301), .o(n_8825) );
no02f80 g561143 ( .a(n_8302), .b(n_8301), .o(n_10343) );
na02f80 g561144 ( .a(n_6896), .b(n_6895), .o(n_6897) );
no02f80 g561145 ( .a(n_6893), .b(n_6892), .o(n_6894) );
na02f80 g561146 ( .a(n_6890), .b(n_6889), .o(n_6891) );
no02f80 g561147 ( .a(n_6240), .b(n_6887), .o(n_6888) );
no02f80 g561148 ( .a(n_6885), .b(n_6884), .o(n_6886) );
no02f80 g561149 ( .a(n_9403), .b(n_8299), .o(n_8300) );
no02f80 g561150 ( .a(n_7711), .b(n_7710), .o(n_7712) );
na02f80 g561151 ( .a(n_7708), .b(n_7707), .o(n_7709) );
na02f80 g561152 ( .a(n_6254), .b(n_7705), .o(n_7706) );
na02f80 g561153 ( .a(n_7703), .b(n_7702), .o(n_7704) );
na02f80 g561154 ( .a(n_6882), .b(n_6881), .o(n_6883) );
no02f80 g561155 ( .a(n_9436), .b(n_8297), .o(n_8298) );
na02f80 g561156 ( .a(n_9436), .b(n_8295), .o(n_8296) );
no02f80 g561157 ( .a(n_8858), .b(n_7700), .o(n_7701) );
no02f80 g561158 ( .a(n_7698), .b(n_7697), .o(n_7699) );
na02f80 g561159 ( .a(n_5841), .b(n_6374), .o(n_7696) );
na02f80 g561160 ( .a(n_7694), .b(n_7693), .o(n_7695) );
na02f80 g561161 ( .a(n_7691), .b(n_7690), .o(n_7692) );
no02f80 g561162 ( .a(n_7688), .b(n_7687), .o(n_7689) );
in01f80 g561163 ( .a(n_8293), .o(n_8294) );
na02f80 g561164 ( .a(n_8936), .b(n_7686), .o(n_8293) );
no02f80 g561165 ( .a(n_6879), .b(n_6878), .o(n_6880) );
na02f80 g561166 ( .a(n_6876), .b(n_6875), .o(n_6877) );
no02f80 g561167 ( .a(n_7684), .b(n_7683), .o(n_7685) );
no02f80 g561168 ( .a(n_6873), .b(n_6872), .o(n_6874) );
no02f80 g561169 ( .a(n_9053), .b(n_7681), .o(n_7682) );
no02f80 g561170 ( .a(n_6870), .b(n_6869), .o(n_6871) );
na02f80 g561171 ( .a(n_8859), .b(n_7679), .o(n_7680) );
no02f80 g561172 ( .a(n_8927), .b(n_7677), .o(n_7678) );
na02f80 g561173 ( .a(n_8927), .b(n_7675), .o(n_7676) );
no02f80 g561174 ( .a(n_7673), .b(n_7672), .o(n_7674) );
no02f80 g561175 ( .a(n_7670), .b(n_7669), .o(n_7671) );
na02f80 g561176 ( .a(n_5836), .b(n_6360), .o(n_7668) );
no02f80 g561177 ( .a(n_7666), .b(n_7665), .o(n_7667) );
no02f80 g561178 ( .a(n_7663), .b(n_7662), .o(n_7664) );
na02f80 g561179 ( .a(n_11097), .b(n_7660), .o(n_7661) );
na02f80 g561180 ( .a(n_8594), .b(n_7404), .o(n_7405) );
no02f80 g561181 ( .a(FE_OFN787_n_8855), .b(n_7658), .o(n_7659) );
na02f80 g561182 ( .a(n_6868), .b(n_6867), .o(n_10725) );
na02f80 g561183 ( .a(n_8011), .b(n_8010), .o(n_8012) );
na02f80 g561184 ( .a(n_7656), .b(n_7655), .o(n_7657) );
na02f80 g561185 ( .a(n_5829), .b(n_6367), .o(n_7654) );
in01f80 g561186 ( .a(n_8291), .o(n_8292) );
na02f80 g561187 ( .a(n_11557), .b(n_7653), .o(n_8291) );
no02f80 g561188 ( .a(n_9249), .b(n_10194), .o(n_6866) );
no02f80 g561189 ( .a(n_7651), .b(n_7650), .o(n_7652) );
na02f80 g561190 ( .a(n_8710), .b(n_7648), .o(n_7649) );
na02f80 g561191 ( .a(n_7646), .b(n_7645), .o(n_7647) );
na02f80 g561192 ( .a(FE_OFN708_n_8059), .b(n_6864), .o(n_6865) );
na02f80 g561193 ( .a(n_8064), .b(n_6862), .o(n_6863) );
in01f80 g561194 ( .a(n_8289), .o(n_8290) );
no03m80 g561195 ( .a(n_7589), .b(n_7590), .c(n_7591), .o(n_8289) );
in01f80 g561196 ( .a(n_7643), .o(n_9858) );
no02f80 g561197 ( .a(n_6861), .b(n_6860), .o(n_7643) );
na02f80 g561198 ( .a(n_8558), .b(n_7641), .o(n_7642) );
na02f80 g561199 ( .a(n_8072), .b(n_6858), .o(n_6859) );
no02f80 g561200 ( .a(n_8052), .b(n_6856), .o(n_6857) );
no02f80 g561201 ( .a(n_8050), .b(FE_OFN971_n_6854), .o(n_6855) );
na02f80 g561202 ( .a(FE_OFN873_n_8070), .b(n_6852), .o(n_6853) );
no02f80 g561203 ( .a(n_8791), .b(n_7639), .o(n_7640) );
oa12f80 g561204 ( .a(n_3200), .b(n_4154), .c(n_3731), .o(n_11238) );
oa12f80 g561205 ( .a(n_2830), .b(n_4649), .c(n_3776), .o(n_11232) );
oa12f80 g561206 ( .a(n_3345), .b(n_4208), .c(n_3732), .o(n_11252) );
oa12f80 g561207 ( .a(n_3336), .b(n_4648), .c(n_3393), .o(n_11214) );
oa12f80 g561208 ( .a(n_2841), .b(n_4650), .c(n_4022), .o(n_11223) );
na02f80 g561209 ( .a(n_8919), .b(n_8920), .o(n_7638) );
no02f80 g561210 ( .a(n_6850), .b(n_6849), .o(n_6851) );
no02f80 g561211 ( .a(n_6847), .b(n_6846), .o(n_6848) );
na02f80 g561212 ( .a(n_11103), .b(n_6356), .o(n_7637) );
no02f80 g561213 ( .a(n_6844), .b(n_6843), .o(n_6845) );
no02f80 g561214 ( .a(n_9179), .b(n_8287), .o(n_8288) );
no02f80 g561215 ( .a(n_6640), .b(FE_OFN548_n_10452), .o(n_7636) );
na02f80 g561216 ( .a(FE_OFN1280_n_8068), .b(n_6841), .o(n_6842) );
na02f80 g561217 ( .a(n_11094), .b(n_9582), .o(n_6840) );
no02f80 g561218 ( .a(n_6838), .b(n_6837), .o(n_6839) );
na02f80 g561219 ( .a(n_8956), .b(n_8285), .o(n_8286) );
no02f80 g561220 ( .a(n_8903), .b(n_7634), .o(n_7635) );
in01f80 g561221 ( .a(n_10419), .o(n_14533) );
no02f80 g561222 ( .a(n_7428), .b(n_7427), .o(n_10419) );
in01f80 g561223 ( .a(n_8283), .o(n_8284) );
na02f80 g561224 ( .a(n_7428), .b(n_7427), .o(n_8283) );
in01f80 g561225 ( .a(n_8282), .o(n_9846) );
na02f80 g561226 ( .a(n_7633), .b(n_7632), .o(n_8282) );
in01f80 g561227 ( .a(n_7631), .o(n_10721) );
no02f80 g561228 ( .a(n_6836), .b(n_6835), .o(n_7631) );
na02f80 g561229 ( .a(n_6834), .b(n_6833), .o(n_9848) );
no02f80 g561230 ( .a(n_6832), .b(n_6831), .o(n_9844) );
in01f80 g561231 ( .a(n_8901), .o(n_11070) );
na02f80 g561232 ( .a(n_7630), .b(n_7629), .o(n_8901) );
no02f80 g561233 ( .a(n_7625), .b(n_7624), .o(n_9466) );
in01f80 g561234 ( .a(n_8823), .o(n_8824) );
no02f80 g561235 ( .a(n_8281), .b(n_8280), .o(n_8823) );
na02f80 g561236 ( .a(n_8281), .b(n_8280), .o(n_10342) );
in01f80 g561237 ( .a(n_8278), .o(n_8279) );
na02f80 g561238 ( .a(n_7627), .b(n_7626), .o(n_8278) );
no02f80 g561239 ( .a(n_7627), .b(n_7626), .o(n_9465) );
oa12f80 g561240 ( .a(n_3804), .b(n_7191), .c(n_3807), .o(n_8610) );
in01f80 g561241 ( .a(n_8276), .o(n_8277) );
na02f80 g561242 ( .a(n_7625), .b(n_7624), .o(n_8276) );
no02f80 g561243 ( .a(n_6829), .b(n_6828), .o(n_6830) );
no02f80 g561244 ( .a(n_8573), .b(n_7622), .o(n_7623) );
no02f80 g561245 ( .a(n_7620), .b(n_7619), .o(n_7621) );
in01f80 g561246 ( .a(n_11458), .o(n_8275) );
na02f80 g561247 ( .a(n_7620), .b(n_7457), .o(n_11458) );
na02f80 g561248 ( .a(n_8017), .b(n_6704), .o(n_6705) );
ao12f80 g561249 ( .a(n_4989), .b(n_6652), .c(n_8397), .o(n_9342) );
no02f80 g561250 ( .a(n_8055), .b(n_6826), .o(n_6827) );
na02f80 g561251 ( .a(n_8031), .b(FE_OFN676_n_6824), .o(n_6825) );
in01f80 g561252 ( .a(n_8273), .o(n_8274) );
no03m80 g561253 ( .a(n_7595), .b(n_7596), .c(n_7597), .o(n_8273) );
no02f80 g561254 ( .a(n_8051), .b(FE_OFN973_n_6822), .o(n_6823) );
ao12f80 g561255 ( .a(n_6325), .b(n_4588), .c(x_in_57_14), .o(n_8196) );
no02f80 g561256 ( .a(n_8190), .b(n_6820), .o(n_6821) );
na02f80 g561257 ( .a(n_6818), .b(n_6817), .o(n_6819) );
no02f80 g561258 ( .a(n_6815), .b(n_6814), .o(n_6816) );
no02f80 g561259 ( .a(n_6812), .b(n_6811), .o(n_6813) );
in01f80 g561260 ( .a(n_8271), .o(n_8272) );
no03m80 g561261 ( .a(n_7592), .b(n_7593), .c(n_7594), .o(n_8271) );
no02f80 g561262 ( .a(n_7617), .b(FE_OFN845_n_7616), .o(n_7618) );
na02f80 g561263 ( .a(n_6809), .b(n_6808), .o(n_6810) );
no02f80 g561264 ( .a(n_6806), .b(n_6805), .o(n_6807) );
no02f80 g561265 ( .a(n_6803), .b(n_6802), .o(n_6804) );
no02f80 g561266 ( .a(n_7614), .b(n_7613), .o(n_7615) );
ao12f80 g561267 ( .a(n_3151), .b(n_5878), .c(n_4863), .o(n_6801) );
na02f80 g561268 ( .a(n_8570), .b(n_7611), .o(n_7612) );
no02f80 g561269 ( .a(n_8858), .b(n_4880), .o(n_7610) );
no02f80 g561270 ( .a(n_8859), .b(n_4864), .o(n_7609) );
in01f80 g561271 ( .a(n_8269), .o(n_8270) );
na02f80 g561272 ( .a(n_7391), .b(n_7390), .o(n_8269) );
no02f80 g561273 ( .a(n_7391), .b(n_7390), .o(n_9464) );
na02f80 g561274 ( .a(n_8768), .b(n_8569), .o(n_7608) );
no02f80 g561275 ( .a(n_7606), .b(n_7605), .o(n_7607) );
no02f80 g561276 ( .a(n_8267), .b(n_8266), .o(n_8268) );
no02f80 g561277 ( .a(n_9425), .b(n_9424), .o(n_8265) );
no02f80 g561278 ( .a(n_7603), .b(n_7602), .o(n_7604) );
no02f80 g561279 ( .a(n_9225), .b(n_8441), .o(n_6800) );
na02f80 g561280 ( .a(n_6798), .b(n_6797), .o(n_6799) );
no02f80 g561281 ( .a(n_6795), .b(n_3767), .o(n_6796) );
oa12f80 g561282 ( .a(n_7945), .b(n_5844), .c(n_5838), .o(n_6794) );
no02f80 g561283 ( .a(n_6793), .b(n_6792), .o(n_9803) );
na02f80 g561284 ( .a(n_8062), .b(n_6790), .o(n_6791) );
oa12f80 g561285 ( .a(n_4834), .b(n_5435), .c(n_2534), .o(n_6400) );
in01f80 g561286 ( .a(n_7600), .o(n_7601) );
ao12f80 g561287 ( .a(n_2290), .b(n_6789), .c(n_6788), .o(n_7600) );
oa12f80 g561288 ( .a(n_9187), .b(n_7019), .c(n_6580), .o(n_12104) );
ao12f80 g561289 ( .a(n_7599), .b(n_9540), .c(n_7598), .o(n_9178) );
ao12f80 g561290 ( .a(n_5439), .b(n_11320), .c(n_6643), .o(n_13939) );
oa12f80 g561291 ( .a(n_7597), .b(n_7596), .c(n_7595), .o(n_9558) );
oa12f80 g561292 ( .a(n_7594), .b(n_7593), .c(n_7592), .o(n_9557) );
oa12f80 g561293 ( .a(n_5864), .b(n_7958), .c(n_5863), .o(n_11627) );
oa22f80 g561294 ( .a(n_10851), .b(n_3325), .c(FE_OFN1073_n_6399), .d(n_2028), .o(n_13279) );
in01f80 g561295 ( .a(n_8802), .o(n_6787) );
oa12f80 g561296 ( .a(n_6769), .b(n_5784), .c(n_3195), .o(n_8802) );
oa12f80 g561297 ( .a(n_7591), .b(n_7590), .c(n_7589), .o(n_9554) );
oa12f80 g561298 ( .a(n_8769), .b(n_6739), .c(n_6740), .o(n_8779) );
na03f80 g561299 ( .a(n_4589), .b(n_6326), .c(n_3821), .o(n_8264) );
oa12f80 g561300 ( .a(n_4842), .b(n_7478), .c(n_7477), .o(n_9186) );
ao12f80 g561301 ( .a(n_7058), .b(n_9964), .c(n_7057), .o(n_13703) );
na02f80 g561302 ( .a(n_4917), .b(n_8747), .o(n_6786) );
no02f80 g561303 ( .a(n_5442), .b(n_4733), .o(n_13424) );
in01f80 g561304 ( .a(n_9623), .o(n_7587) );
oa22f80 g561305 ( .a(n_4735), .b(n_6785), .c(n_9072), .d(n_6784), .o(n_9623) );
in01f80 g561306 ( .a(n_8263), .o(n_14282) );
ao12f80 g561307 ( .a(n_6035), .b(n_9010), .c(n_7481), .o(n_8263) );
ao22s80 g561308 ( .a(n_4718), .b(n_6783), .c(n_3490), .d(FE_OFN801_n_6782), .o(n_11848) );
in01f80 g561309 ( .a(n_14278), .o(n_8822) );
no02f80 g561310 ( .a(n_6642), .b(n_5190), .o(n_14278) );
oa22f80 g561311 ( .a(n_6398), .b(n_2053), .c(x_in_23_12), .d(x_in_23_10), .o(n_8797) );
oa22f80 g561312 ( .a(n_6397), .b(n_2293), .c(x_in_15_12), .d(x_in_15_10), .o(n_8806) );
oa22f80 g561313 ( .a(n_6396), .b(n_2136), .c(x_in_47_12), .d(x_in_47_10), .o(n_8805) );
oa22f80 g561314 ( .a(n_6395), .b(n_2252), .c(x_in_55_12), .d(x_in_55_10), .o(n_8799) );
oa22f80 g561315 ( .a(n_6394), .b(n_2291), .c(x_in_31_12), .d(x_in_31_10), .o(n_8798) );
oa22f80 g561316 ( .a(n_6393), .b(n_2076), .c(x_in_63_12), .d(x_in_63_10), .o(n_8804) );
ao12f80 g561317 ( .a(n_6031), .b(n_9082), .c(n_7551), .o(n_14008) );
in01f80 g561318 ( .a(n_8262), .o(n_13929) );
oa22f80 g561319 ( .a(n_4968), .b(n_7540), .c(n_8982), .d(n_7541), .o(n_8262) );
oa22f80 g561320 ( .a(n_5186), .b(n_7479), .c(n_9066), .d(n_7480), .o(n_14268) );
no02f80 g561321 ( .a(n_4839), .b(n_8108), .o(n_6392) );
na02f80 g561322 ( .a(n_6467), .b(n_9088), .o(n_8261) );
no02f80 g561323 ( .a(n_5578), .b(x_in_9_13), .o(n_8705) );
in01f80 g561324 ( .a(n_14452), .o(n_8260) );
no02f80 g561325 ( .a(n_6036), .b(n_4703), .o(n_14452) );
oa22f80 g561326 ( .a(n_4356), .b(n_6747), .c(n_8674), .d(n_6748), .o(n_14792) );
oa12f80 g561327 ( .a(n_7736), .b(n_8704), .c(x_in_9_12), .o(n_7586) );
oa12f80 g561328 ( .a(n_5434), .b(n_5485), .c(n_2119), .o(n_11997) );
ao12f80 g561329 ( .a(n_5165), .b(n_7204), .c(n_8305), .o(n_10892) );
oa12f80 g561330 ( .a(n_5300), .b(n_5299), .c(n_6781), .o(n_14097) );
in01f80 g561331 ( .a(n_7584), .o(n_7585) );
oa22f80 g561332 ( .a(n_4695), .b(n_6780), .c(n_9139), .d(n_6779), .o(n_7584) );
oa12f80 g561333 ( .a(n_5710), .b(n_5862), .c(n_5848), .o(n_10712) );
in01f80 g561334 ( .a(n_7582), .o(n_7583) );
ao22s80 g561335 ( .a(n_4684), .b(n_6828), .c(n_5320), .d(n_5321), .o(n_7582) );
oa22f80 g561336 ( .a(n_5177), .b(n_7448), .c(n_9135), .d(n_7449), .o(n_11858) );
ao12f80 g561337 ( .a(n_5420), .b(n_3570), .c(n_6713), .o(n_11118) );
oa12f80 g561338 ( .a(n_6777), .b(n_6776), .c(n_6775), .o(n_6778) );
oa12f80 g561339 ( .a(n_5724), .b(n_7581), .c(n_5835), .o(n_11853) );
in01f80 g561340 ( .a(n_8258), .o(n_8259) );
ao22s80 g561341 ( .a(n_5196), .b(n_5969), .c(n_7847), .d(n_5747), .o(n_8258) );
oa22f80 g561342 ( .a(n_5171), .b(n_7552), .c(n_9132), .d(n_7553), .o(n_11940) );
oa22f80 g561343 ( .a(n_4334), .b(n_7662), .c(n_5830), .d(n_5825), .o(n_10757) );
no03m80 g561344 ( .a(n_6763), .b(n_6764), .c(n_6773), .o(n_6774) );
in01f80 g561345 ( .a(n_8256), .o(n_8257) );
oa22f80 g561346 ( .a(n_5167), .b(n_7467), .c(n_9129), .d(n_7466), .o(n_8256) );
ao12f80 g561347 ( .a(n_6008), .b(n_3651), .c(n_6749), .o(n_11160) );
in01f80 g561348 ( .a(n_7579), .o(n_7580) );
oa22f80 g561349 ( .a(n_4678), .b(n_6743), .c(n_8722), .d(n_6744), .o(n_7579) );
in01f80 g561350 ( .a(n_7577), .o(n_7578) );
ao12f80 g561351 ( .a(n_4966), .b(n_5669), .c(x_in_17_3), .o(n_7577) );
oa22f80 g561352 ( .a(n_5160), .b(n_7502), .c(n_9123), .d(n_7503), .o(n_11776) );
in01f80 g561353 ( .a(n_8254), .o(n_8255) );
oa12f80 g561354 ( .a(n_6006), .b(n_8734), .c(n_6709), .o(n_8254) );
oa12f80 g561355 ( .a(n_6630), .b(n_8731), .c(n_6715), .o(n_11123) );
ao22s80 g561356 ( .a(n_4675), .b(n_6772), .c(n_4028), .d(FE_OFN803_n_6771), .o(n_13105) );
in01f80 g561357 ( .a(n_8252), .o(n_8253) );
oa22f80 g561358 ( .a(n_5069), .b(n_6728), .c(n_8719), .d(n_6727), .o(n_8252) );
ao12f80 g561359 ( .a(n_5412), .b(n_5345), .c(n_5346), .o(n_10735) );
in01f80 g561360 ( .a(n_7573), .o(n_9601) );
oa22f80 g561361 ( .a(n_4580), .b(n_6770), .c(FE_OFN1089_n_8985), .d(n_6769), .o(n_7573) );
oa12f80 g561362 ( .a(n_5997), .b(n_5295), .c(n_5296), .o(n_9809) );
in01f80 g561363 ( .a(n_8820), .o(n_8821) );
oa12f80 g561364 ( .a(n_6627), .b(n_8728), .c(FE_OFN692_n_6708), .o(n_8820) );
ao12f80 g561365 ( .a(n_5410), .b(n_8297), .c(x_in_37_5), .o(n_11436) );
in01f80 g561366 ( .a(FE_OFN1085_n_14427), .o(n_7572) );
oa22f80 g561367 ( .a(n_4653), .b(n_6768), .c(FE_OFN1274_n_8977), .d(n_6767), .o(n_14427) );
oa22f80 g561368 ( .a(n_4147), .b(n_7672), .c(n_5837), .d(n_5900), .o(n_12432) );
oa12f80 g561369 ( .a(n_6045), .b(n_8092), .c(n_8522), .o(n_13444) );
ao22s80 g561370 ( .a(n_5145), .b(n_7435), .c(n_7571), .d(x_in_21_2), .o(n_13909) );
ao12f80 g561371 ( .a(n_6012), .b(n_9338), .c(n_6724), .o(n_13895) );
oa22f80 g561372 ( .a(n_4925), .b(n_7442), .c(n_8971), .d(n_7443), .o(n_14273) );
ao12f80 g561373 ( .a(n_6009), .b(n_4938), .c(n_7445), .o(n_13864) );
in01f80 g561374 ( .a(n_7569), .o(n_7570) );
ao22s80 g561375 ( .a(n_4181), .b(n_6766), .c(n_3681), .d(x_in_37_11), .o(n_7569) );
oa22f80 g561376 ( .a(n_3377), .b(n_7147), .c(n_5674), .d(n_5866), .o(n_13210) );
in01f80 g561377 ( .a(n_8250), .o(n_8251) );
ao22s80 g561378 ( .a(n_5139), .b(n_5867), .c(n_7602), .d(n_5868), .o(n_8250) );
in01f80 g561379 ( .a(n_14226), .o(n_7568) );
oa22f80 g561380 ( .a(n_4398), .b(n_6722), .c(FE_OFN1091_n_8621), .d(n_6723), .o(n_14226) );
oa12f80 g561381 ( .a(n_6043), .b(n_8142), .c(n_8929), .o(n_13403) );
no02f80 g561382 ( .a(n_5486), .b(n_4402), .o(n_8757) );
oa22f80 g561383 ( .a(n_4658), .b(n_10224), .c(n_8546), .d(n_6984), .o(n_12673) );
in01f80 g561384 ( .a(n_8818), .o(n_8819) );
oa12f80 g561385 ( .a(n_6639), .b(n_6573), .c(n_5137), .o(n_8818) );
oa22f80 g561386 ( .a(n_3426), .b(n_6391), .c(n_6390), .d(n_8696), .o(n_8193) );
ao12f80 g561387 ( .a(n_7489), .b(n_5783), .c(n_7490), .o(n_9886) );
ao12f80 g561388 ( .a(n_6776), .b(n_6777), .c(n_5134), .o(n_7567) );
ao12f80 g561389 ( .a(n_5397), .b(n_5384), .c(n_5383), .o(n_8788) );
in01f80 g561390 ( .a(n_8816), .o(n_8817) );
ao22s80 g561391 ( .a(n_5791), .b(n_5892), .c(n_6475), .d(n_2391), .o(n_8816) );
in01f80 g561392 ( .a(n_8248), .o(n_8249) );
oa22f80 g561393 ( .a(n_5141), .b(n_7557), .c(n_7556), .d(n_6746), .o(n_8248) );
oa12f80 g561394 ( .a(n_6773), .b(n_6764), .c(n_6763), .o(n_6765) );
in01f80 g561395 ( .a(n_8814), .o(n_8815) );
oa22f80 g561396 ( .a(n_5796), .b(n_7518), .c(n_7519), .d(n_10477), .o(n_8814) );
ao12f80 g561397 ( .a(n_5948), .b(n_3917), .c(x_in_53_2), .o(n_7566) );
oa12f80 g561398 ( .a(n_4328), .b(n_4826), .c(n_4327), .o(n_8800) );
in01f80 g561399 ( .a(n_9639), .o(n_8247) );
ao12f80 g561400 ( .a(n_6132), .b(n_6131), .c(n_6373), .o(n_9639) );
in01f80 g561401 ( .a(n_7564), .o(n_7565) );
oa12f80 g561402 ( .a(n_5610), .b(n_5769), .c(x_in_61_13), .o(n_7564) );
oa22f80 g561403 ( .a(n_5092), .b(n_6769), .c(n_6770), .d(n_4579), .o(n_8986) );
oa12f80 g561404 ( .a(n_4380), .b(n_6389), .c(n_4740), .o(n_8158) );
in01f80 g561405 ( .a(n_7563), .o(n_9192) );
oa12f80 g561406 ( .a(n_5504), .b(n_5503), .c(x_in_59_3), .o(n_7563) );
in01f80 g561407 ( .a(n_10404), .o(n_8246) );
ao12f80 g561408 ( .a(n_6208), .b(n_6207), .c(n_6437), .o(n_10404) );
oa12f80 g561409 ( .a(n_5625), .b(n_5624), .c(x_in_59_13), .o(n_8683) );
ao12f80 g561410 ( .a(n_5463), .b(n_5784), .c(n_9088), .o(n_9335) );
in01f80 g561411 ( .a(n_9611), .o(n_7562) );
oa12f80 g561412 ( .a(n_5636), .b(n_5635), .c(n_5916), .o(n_9611) );
ao12f80 g561413 ( .a(n_4856), .b(n_6388), .c(n_5695), .o(n_8153) );
ao22s80 g561414 ( .a(n_5148), .b(n_6366), .c(n_8086), .d(n_4196), .o(n_13393) );
oa12f80 g561415 ( .a(n_6048), .b(n_8089), .c(n_6387), .o(n_13859) );
in01f80 g561416 ( .a(n_9607), .o(n_9609) );
oa22f80 g561417 ( .a(n_4417), .b(n_6760), .c(n_4418), .d(n_9604), .o(n_9607) );
ao12f80 g561418 ( .a(n_6655), .b(n_6654), .c(n_6653), .o(n_9521) );
in01f80 g561419 ( .a(n_9576), .o(n_7561) );
oa22f80 g561420 ( .a(n_4796), .b(n_8482), .c(n_5496), .d(x_in_59_11), .o(n_9576) );
oa12f80 g561421 ( .a(n_4865), .b(n_6047), .c(n_6387), .o(n_8090) );
oa12f80 g561422 ( .a(n_5518), .b(n_5517), .c(x_in_25_4), .o(n_10314) );
in01f80 g561423 ( .a(n_10425), .o(n_8245) );
ao12f80 g561424 ( .a(n_6066), .b(n_6065), .c(n_6064), .o(n_10425) );
ao22s80 g561425 ( .a(n_6308), .b(n_7560), .c(n_7559), .d(n_6307), .o(n_9075) );
in01f80 g561426 ( .a(n_9593), .o(n_7558) );
oa12f80 g561427 ( .a(n_5552), .b(n_5551), .c(x_in_11_6), .o(n_9593) );
ao22s80 g561428 ( .a(n_7557), .b(n_5140), .c(n_5078), .d(n_7556), .o(n_9107) );
ao22s80 g561429 ( .a(n_4912), .b(n_6386), .c(n_6385), .d(n_4911), .o(n_8104) );
in01f80 g561430 ( .a(n_6758), .o(n_6759) );
oa22f80 g561431 ( .a(n_6384), .b(n_6383), .c(n_4001), .d(n_6382), .o(n_6758) );
ao12f80 g561432 ( .a(n_5609), .b(n_5608), .c(x_in_43_8), .o(n_6757) );
in01f80 g561433 ( .a(n_9269), .o(n_6756) );
oa12f80 g561434 ( .a(n_4849), .b(n_4848), .c(x_in_61_14), .o(n_9269) );
ao12f80 g561435 ( .a(n_4838), .b(n_6381), .c(n_5567), .o(n_8148) );
ao22s80 g561436 ( .a(n_7555), .b(n_3832), .c(n_5081), .d(n_7554), .o(n_9089) );
in01f80 g561437 ( .a(n_9271), .o(n_6755) );
ao22s80 g561438 ( .a(n_5041), .b(n_6380), .c(n_3799), .d(x_in_3_11), .o(n_9271) );
ao12f80 g561439 ( .a(n_4889), .b(n_6379), .c(n_5633), .o(n_8155) );
oa22f80 g561440 ( .a(n_4987), .b(n_7553), .c(n_7552), .d(n_5170), .o(n_9133) );
oa22f80 g561441 ( .a(n_5665), .b(n_6779), .c(n_6780), .d(n_4694), .o(n_9140) );
oa12f80 g561442 ( .a(n_6196), .b(n_7019), .c(n_7385), .o(n_9188) );
in01f80 g561443 ( .a(n_9260), .o(n_6754) );
ao22s80 g561444 ( .a(n_5502), .b(x_in_27_13), .c(n_3583), .d(n_7229), .o(n_9260) );
oa12f80 g561445 ( .a(n_5522), .b(n_5521), .c(x_in_19_5), .o(n_8659) );
ao22s80 g561446 ( .a(n_4631), .b(n_6733), .c(FE_OFN646_n_6732), .d(n_2417), .o(n_8628) );
in01f80 g561447 ( .a(n_8171), .o(n_9278) );
oa22f80 g561448 ( .a(n_4879), .b(n_6380), .c(n_3800), .d(x_in_3_11), .o(n_8171) );
in01f80 g561449 ( .a(n_9674), .o(n_10538) );
oa12f80 g561450 ( .a(n_6186), .b(n_6185), .c(n_6184), .o(n_9674) );
in01f80 g561451 ( .a(n_9653), .o(n_9109) );
oa12f80 g561452 ( .a(n_5462), .b(n_5461), .c(n_5460), .o(n_9653) );
in01f80 g561453 ( .a(n_10527), .o(n_9452) );
oa12f80 g561454 ( .a(n_6199), .b(n_6198), .c(FE_OFN1262_n_6197), .o(n_10527) );
ao12f80 g561455 ( .a(n_6277), .b(n_6276), .c(n_7551), .o(n_9083) );
ao12f80 g561456 ( .a(n_5529), .b(n_5528), .c(x_in_3_8), .o(n_9580) );
in01f80 g561457 ( .a(n_9328), .o(n_7550) );
oa12f80 g561458 ( .a(n_5644), .b(n_5643), .c(n_5642), .o(n_9328) );
in01f80 g561459 ( .a(n_10530), .o(n_8244) );
ao12f80 g561460 ( .a(n_6192), .b(n_6191), .c(n_6190), .o(n_10530) );
in01f80 g561461 ( .a(n_7548), .o(n_7549) );
oa22f80 g561462 ( .a(n_4478), .b(x_in_31_12), .c(n_6394), .d(n_6753), .o(n_7548) );
oa12f80 g561463 ( .a(n_5560), .b(n_5559), .c(n_5558), .o(n_9301) );
in01f80 g561464 ( .a(n_10542), .o(n_10532) );
oa12f80 g561465 ( .a(n_6171), .b(n_6170), .c(n_6169), .o(n_10542) );
in01f80 g561466 ( .a(n_10397), .o(n_9507) );
oa12f80 g561467 ( .a(n_6163), .b(n_6162), .c(n_6161), .o(n_10397) );
oa22f80 g561468 ( .a(n_3745), .b(FE_OFN239_n_4162), .c(n_1636), .d(FE_OFN1119_rst), .o(n_6752) );
in01f80 g561469 ( .a(n_10504), .o(n_8243) );
oa12f80 g561470 ( .a(n_6189), .b(n_6188), .c(n_6187), .o(n_10504) );
in01f80 g561471 ( .a(n_9341), .o(n_7547) );
ao12f80 g561472 ( .a(n_5533), .b(n_5532), .c(x_in_59_6), .o(n_9341) );
in01f80 g561473 ( .a(n_9025), .o(n_10417) );
oa12f80 g561474 ( .a(n_5715), .b(n_5714), .c(n_5713), .o(n_9025) );
in01f80 g561475 ( .a(n_7545), .o(n_7546) );
oa12f80 g561476 ( .a(n_5444), .b(n_6751), .c(n_6750), .o(n_7545) );
ao12f80 g561477 ( .a(n_5467), .b(n_6007), .c(n_6749), .o(n_8726) );
in01f80 g561478 ( .a(n_9677), .o(n_7544) );
oa12f80 g561479 ( .a(n_5584), .b(n_5583), .c(x_in_59_13), .o(n_9677) );
oa22f80 g561480 ( .a(n_4537), .b(n_6748), .c(n_6747), .d(n_4355), .o(n_8675) );
in01f80 g561481 ( .a(n_9320), .o(n_7543) );
ao12f80 g561482 ( .a(n_5550), .b(n_5549), .c(x_in_11_7), .o(n_9320) );
in01f80 g561483 ( .a(n_9655), .o(n_7542) );
ao12f80 g561484 ( .a(n_5613), .b(n_5612), .c(n_5611), .o(n_9655) );
oa22f80 g561485 ( .a(n_4591), .b(n_6746), .c(n_5626), .d(x_in_3_13), .o(n_8656) );
oa22f80 g561486 ( .a(n_5085), .b(n_7541), .c(n_7540), .d(n_4967), .o(n_8983) );
in01f80 g561487 ( .a(n_10546), .o(n_9518) );
oa12f80 g561488 ( .a(n_6180), .b(n_6179), .c(FE_OFN1260_n_6178), .o(n_10546) );
oa22f80 g561489 ( .a(n_5090), .b(n_6784), .c(n_6785), .d(n_4734), .o(n_9073) );
in01f80 g561490 ( .a(n_10543), .o(n_9462) );
oa12f80 g561491 ( .a(n_6069), .b(n_6068), .c(n_6067), .o(n_10543) );
ao22s80 g561492 ( .a(n_4988), .b(FE_OFN803_n_6771), .c(n_6772), .d(n_4674), .o(n_9121) );
in01f80 g561493 ( .a(n_9164), .o(n_10420) );
oa12f80 g561494 ( .a(n_6177), .b(n_6176), .c(n_6175), .o(n_9164) );
in01f80 g561495 ( .a(n_9784), .o(n_10559) );
oa12f80 g561496 ( .a(n_6202), .b(n_6201), .c(n_6200), .o(n_9784) );
in01f80 g561497 ( .a(n_9219), .o(n_6745) );
ao22s80 g561498 ( .a(n_5065), .b(x_in_27_10), .c(n_3801), .d(n_7417), .o(n_9219) );
oa22f80 g561499 ( .a(n_6783), .b(n_4717), .c(n_5071), .d(FE_OFN801_n_6782), .o(n_9147) );
oa22f80 g561500 ( .a(n_4858), .b(n_6378), .c(n_6377), .d(n_4857), .o(n_8137) );
oa22f80 g561501 ( .a(n_4802), .b(n_6744), .c(n_6743), .d(n_4677), .o(n_8723) );
ao12f80 g561502 ( .a(n_4741), .b(n_4331), .c(n_6389), .o(n_14003) );
ao12f80 g561503 ( .a(n_4975), .b(n_4974), .c(x_in_27_7), .o(n_6742) );
in01f80 g561504 ( .a(n_9080), .o(n_10515) );
oa12f80 g561505 ( .a(n_5765), .b(n_5764), .c(n_5763), .o(n_9080) );
in01f80 g561506 ( .a(n_10395), .o(n_9455) );
oa12f80 g561507 ( .a(n_6028), .b(n_6027), .c(n_6026), .o(n_10395) );
in01f80 g561508 ( .a(n_10551), .o(n_9515) );
oa12f80 g561509 ( .a(n_6144), .b(n_6143), .c(n_6142), .o(n_10551) );
in01f80 g561510 ( .a(n_9290), .o(n_7539) );
ao12f80 g561511 ( .a(n_4996), .b(n_5437), .c(x_in_35_13), .o(n_9290) );
in01f80 g561512 ( .a(n_7537), .o(n_7538) );
oa22f80 g561513 ( .a(n_4477), .b(x_in_23_12), .c(n_6398), .d(n_7323), .o(n_7537) );
in01f80 g561514 ( .a(n_10388), .o(n_10386) );
oa12f80 g561515 ( .a(n_6440), .b(n_6439), .c(n_6438), .o(n_10388) );
oa12f80 g561516 ( .a(n_4827), .b(n_5827), .c(x_in_53_1), .o(n_10754) );
oa22f80 g561517 ( .a(n_3743), .b(FE_OFN230_n_4162), .c(n_694), .d(FE_OFN331_n_4860), .o(n_7536) );
in01f80 g561518 ( .a(n_7534), .o(n_7535) );
ao12f80 g561519 ( .a(n_5458), .b(n_5457), .c(n_5456), .o(n_7534) );
in01f80 g561520 ( .a(n_9300), .o(n_7533) );
ao12f80 g561521 ( .a(n_5237), .b(n_5663), .c(x_in_35_10), .o(n_9300) );
in01f80 g561522 ( .a(n_9669), .o(n_7532) );
oa12f80 g561523 ( .a(n_5566), .b(n_5565), .c(x_in_35_9), .o(n_9669) );
in01f80 g561524 ( .a(n_9665), .o(n_7531) );
oa12f80 g561525 ( .a(n_5588), .b(n_5587), .c(x_in_35_8), .o(n_9665) );
in01f80 g561526 ( .a(n_7529), .o(n_7530) );
oa22f80 g561527 ( .a(n_4505), .b(x_in_15_12), .c(n_6397), .d(n_7338), .o(n_7529) );
na02f80 g561528 ( .a(n_7951), .b(n_3867), .o(n_7528) );
in01f80 g561529 ( .a(n_9315), .o(n_7527) );
ao12f80 g561530 ( .a(n_5607), .b(n_5606), .c(x_in_35_7), .o(n_9315) );
in01f80 g561531 ( .a(n_9663), .o(n_7526) );
ao12f80 g561532 ( .a(n_5523), .b(n_5659), .c(x_in_35_6), .o(n_9663) );
ao12f80 g561533 ( .a(n_5508), .b(n_5507), .c(x_in_35_5), .o(n_8669) );
in01f80 g561534 ( .a(n_10505), .o(n_9500) );
oa12f80 g561535 ( .a(n_6097), .b(n_6096), .c(n_6095), .o(n_10505) );
ao22s80 g561536 ( .a(n_3769), .b(n_6376), .c(n_6375), .d(n_6374), .o(n_8121) );
in01f80 g561537 ( .a(n_10508), .o(n_9488) );
oa12f80 g561538 ( .a(n_6159), .b(n_6158), .c(FE_OFN875_n_6157), .o(n_10508) );
in01f80 g561539 ( .a(n_10502), .o(n_9497) );
oa12f80 g561540 ( .a(n_6156), .b(n_6155), .c(FE_OFN871_n_6154), .o(n_10502) );
in01f80 g561541 ( .a(n_10498), .o(n_9494) );
oa12f80 g561542 ( .a(n_6153), .b(n_6152), .c(FE_OFN867_n_6151), .o(n_10498) );
in01f80 g561543 ( .a(n_10493), .o(n_8242) );
ao12f80 g561544 ( .a(n_6150), .b(n_6149), .c(n_6148), .o(n_10493) );
in01f80 g561545 ( .a(n_10490), .o(n_8241) );
oa12f80 g561546 ( .a(n_6147), .b(n_6146), .c(n_6145), .o(n_10490) );
in01f80 g561547 ( .a(n_9168), .o(n_10488) );
oa12f80 g561548 ( .a(n_6174), .b(n_6173), .c(n_6172), .o(n_9168) );
in01f80 g561549 ( .a(n_8239), .o(n_8240) );
ao12f80 g561550 ( .a(n_5779), .b(n_5778), .c(n_5777), .o(n_8239) );
ao12f80 g561551 ( .a(n_5632), .b(n_6447), .c(x_in_35_13), .o(n_8665) );
in01f80 g561552 ( .a(n_7524), .o(n_7525) );
oa22f80 g561553 ( .a(n_4667), .b(x_in_47_12), .c(n_6396), .d(n_7247), .o(n_7524) );
ao12f80 g561554 ( .a(n_5709), .b(n_5708), .c(FE_OFN765_n_5707), .o(n_13350) );
in01f80 g561555 ( .a(n_9288), .o(n_7523) );
oa12f80 g561556 ( .a(n_5580), .b(n_5579), .c(x_in_35_13), .o(n_9288) );
in01f80 g561557 ( .a(n_9284), .o(n_6741) );
ao12f80 g561558 ( .a(n_4851), .b(n_4850), .c(x_in_61_2), .o(n_9284) );
ao22s80 g561559 ( .a(n_6288), .b(x_in_7_13), .c(n_4569), .d(n_7285), .o(n_8633) );
in01f80 g561560 ( .a(n_9656), .o(n_7522) );
ao12f80 g561561 ( .a(n_5000), .b(n_4999), .c(n_4998), .o(n_9656) );
in01f80 g561562 ( .a(n_9657), .o(n_7521) );
ao12f80 g561563 ( .a(n_5491), .b(n_5490), .c(n_5489), .o(n_9657) );
in01f80 g561564 ( .a(n_9652), .o(n_7520) );
ao12f80 g561565 ( .a(n_5618), .b(n_5617), .c(n_5616), .o(n_9652) );
in01f80 g561566 ( .a(n_8992), .o(n_10514) );
oa12f80 g561567 ( .a(n_6051), .b(n_6050), .c(n_6049), .o(n_8992) );
in01f80 g561568 ( .a(n_9650), .o(n_9114) );
oa12f80 g561569 ( .a(n_5466), .b(n_5465), .c(n_5464), .o(n_9650) );
oa22f80 g561570 ( .a(n_4527), .b(n_6740), .c(n_6739), .d(n_3017), .o(n_8770) );
in01f80 g561571 ( .a(n_9648), .o(n_9647) );
oa12f80 g561572 ( .a(n_5470), .b(n_5469), .c(n_5468), .o(n_9648) );
ao12f80 g561573 ( .a(n_5455), .b(n_5454), .c(n_5453), .o(n_9337) );
oa22f80 g561574 ( .a(n_6371), .b(n_2034), .c(n_5390), .d(x_in_35_1), .o(n_10751) );
oa12f80 g561575 ( .a(n_5648), .b(n_6371), .c(n_5832), .o(n_9318) );
in01f80 g561576 ( .a(n_9614), .o(n_9613) );
oa12f80 g561577 ( .a(n_5687), .b(n_5686), .c(n_5685), .o(n_9614) );
in01f80 g561578 ( .a(n_10479), .o(n_8238) );
oa12f80 g561579 ( .a(n_6232), .b(n_6231), .c(n_6230), .o(n_10479) );
in01f80 g561580 ( .a(n_10474), .o(n_8237) );
ao12f80 g561581 ( .a(n_6141), .b(n_6140), .c(n_6139), .o(n_10474) );
ao12f80 g561582 ( .a(n_6279), .b(n_6278), .c(x_in_59_14), .o(n_23238) );
in01f80 g561583 ( .a(n_8235), .o(n_8236) );
oa22f80 g561584 ( .a(n_5072), .b(n_7519), .c(n_7518), .d(n_5795), .o(n_8235) );
in01f80 g561585 ( .a(n_10478), .o(n_8234) );
ao12f80 g561586 ( .a(n_6287), .b(n_6286), .c(n_6285), .o(n_10478) );
in01f80 g561587 ( .a(n_9642), .o(n_7517) );
ao12f80 g561588 ( .a(n_5495), .b(n_5682), .c(x_in_19_12), .o(n_9642) );
in01f80 g561589 ( .a(n_9644), .o(n_7516) );
ao12f80 g561590 ( .a(n_5343), .b(n_5557), .c(x_in_19_13), .o(n_9644) );
ao12f80 g561591 ( .a(n_5623), .b(n_5622), .c(FE_OFN458_n_5621), .o(n_6736) );
in01f80 g561592 ( .a(n_10461), .o(n_8233) );
ao12f80 g561593 ( .a(n_6138), .b(n_6137), .c(n_6136), .o(n_10461) );
in01f80 g561594 ( .a(n_9640), .o(n_7515) );
ao22s80 g561595 ( .a(n_5487), .b(x_in_19_11), .c(n_4400), .d(n_7765), .o(n_9640) );
in01f80 g561596 ( .a(n_10471), .o(n_9478) );
oa12f80 g561597 ( .a(n_6135), .b(n_6134), .c(n_6133), .o(n_10471) );
in01f80 g561598 ( .a(n_9636), .o(n_7514) );
ao12f80 g561599 ( .a(n_5539), .b(n_5664), .c(x_in_19_10), .o(n_9636) );
in01f80 g561600 ( .a(n_10476), .o(n_9485) );
oa12f80 g561601 ( .a(n_6091), .b(n_6090), .c(FE_OFN1222_n_6089), .o(n_10476) );
in01f80 g561602 ( .a(n_10468), .o(n_8232) );
oa12f80 g561603 ( .a(n_6446), .b(n_6445), .c(FE_OFN706_n_6444), .o(n_10468) );
in01f80 g561604 ( .a(n_9634), .o(n_7513) );
ao12f80 g561605 ( .a(n_5254), .b(n_5538), .c(x_in_19_9), .o(n_9634) );
in01f80 g561606 ( .a(n_10466), .o(n_8231) );
ao12f80 g561607 ( .a(n_6077), .b(n_6076), .c(n_6075), .o(n_10466) );
in01f80 g561608 ( .a(n_10463), .o(n_8230) );
oa12f80 g561609 ( .a(n_5726), .b(n_5725), .c(n_6017), .o(n_10463) );
in01f80 g561610 ( .a(n_9632), .o(n_7512) );
ao12f80 g561611 ( .a(n_5534), .b(n_5555), .c(x_in_19_8), .o(n_9632) );
in01f80 g561612 ( .a(n_10459), .o(n_8229) );
ao12f80 g561613 ( .a(n_6093), .b(n_6092), .c(n_6315), .o(n_10459) );
ao12f80 g561614 ( .a(n_5735), .b(n_5734), .c(n_6641), .o(n_9008) );
in01f80 g561615 ( .a(n_10457), .o(n_8228) );
oa12f80 g561616 ( .a(n_6130), .b(n_6129), .c(n_6128), .o(n_10457) );
in01f80 g561617 ( .a(n_9158), .o(n_10454) );
oa12f80 g561618 ( .a(n_6195), .b(n_6194), .c(n_6193), .o(n_9158) );
in01f80 g561619 ( .a(n_9267), .o(n_7511) );
ao12f80 g561620 ( .a(n_5536), .b(n_5535), .c(x_in_19_6), .o(n_9267) );
oa12f80 g561621 ( .a(n_6319), .b(n_6318), .c(n_6317), .o(n_9045) );
oa12f80 g561622 ( .a(n_6074), .b(n_6073), .c(FE_OFN550_n_6072), .o(n_10447) );
ao12f80 g561623 ( .a(n_6060), .b(n_6059), .c(n_6058), .o(n_10446) );
in01f80 g561624 ( .a(n_7509), .o(n_7510) );
ao12f80 g561625 ( .a(n_5511), .b(n_5510), .c(x_in_3_5), .o(n_7509) );
in01f80 g561626 ( .a(n_9262), .o(n_6735) );
ao22s80 g561627 ( .a(n_5488), .b(n_7765), .c(n_3728), .d(x_in_19_11), .o(n_9262) );
in01f80 g561628 ( .a(n_9649), .o(n_7508) );
ao12f80 g561629 ( .a(n_5480), .b(n_5479), .c(n_5478), .o(n_9649) );
in01f80 g561630 ( .a(n_9853), .o(n_8227) );
oa12f80 g561631 ( .a(n_6124), .b(n_6123), .c(n_6122), .o(n_9853) );
in01f80 g561632 ( .a(n_10354), .o(n_9474) );
oa12f80 g561633 ( .a(n_6121), .b(n_6120), .c(n_6119), .o(n_10354) );
ao12f80 g561634 ( .a(n_5527), .b(n_5667), .c(x_in_3_10), .o(n_9583) );
in01f80 g561635 ( .a(n_10445), .o(n_9491) );
oa12f80 g561636 ( .a(n_6118), .b(n_6117), .c(FE_OFN1278_n_6116), .o(n_10445) );
in01f80 g561637 ( .a(n_10443), .o(n_9471) );
oa12f80 g561638 ( .a(n_6106), .b(n_6105), .c(n_6104), .o(n_10443) );
in01f80 g561639 ( .a(n_10369), .o(n_9524) );
oa12f80 g561640 ( .a(n_6115), .b(n_6114), .c(n_6113), .o(n_10369) );
in01f80 g561641 ( .a(n_10368), .o(n_8226) );
oa12f80 g561642 ( .a(n_6112), .b(n_6111), .c(n_6110), .o(n_10368) );
in01f80 g561643 ( .a(n_10438), .o(n_8225) );
ao12f80 g561644 ( .a(n_6109), .b(n_6108), .c(n_6107), .o(n_10438) );
in01f80 g561645 ( .a(n_10436), .o(n_8224) );
oa12f80 g561646 ( .a(n_6103), .b(n_6102), .c(n_6101), .o(n_10436) );
in01f80 g561647 ( .a(n_9275), .o(n_6734) );
ao22s80 g561648 ( .a(n_5493), .b(x_in_27_11), .c(n_4083), .d(n_8513), .o(n_9275) );
in01f80 g561649 ( .a(n_9161), .o(n_10433) );
oa12f80 g561650 ( .a(n_6100), .b(n_6099), .c(n_6098), .o(n_9161) );
in01f80 g561651 ( .a(n_7506), .o(n_7507) );
ao12f80 g561652 ( .a(n_5449), .b(n_5448), .c(n_5447), .o(n_7506) );
in01f80 g561653 ( .a(n_10401), .o(n_8223) );
oa12f80 g561654 ( .a(n_6206), .b(n_6205), .c(n_6204), .o(n_10401) );
in01f80 g561655 ( .a(n_7504), .o(n_7505) );
oa22f80 g561656 ( .a(n_4874), .b(x_in_63_12), .c(n_6393), .d(n_8206), .o(n_7504) );
oa22f80 g561657 ( .a(n_4947), .b(n_7503), .c(n_7502), .d(n_5159), .o(n_9124) );
in01f80 g561658 ( .a(n_7500), .o(n_7501) );
ao12f80 g561659 ( .a(n_5671), .b(n_5670), .c(x_in_43_5), .o(n_7500) );
in01f80 g561660 ( .a(n_10432), .o(n_10427) );
oa22f80 g561661 ( .a(n_4985), .b(n_7499), .c(n_4986), .d(n_7498), .o(n_10432) );
ao12f80 g561662 ( .a(n_6127), .b(n_6126), .c(n_6125), .o(n_10449) );
in01f80 g561663 ( .a(n_9330), .o(n_7497) );
oa12f80 g561664 ( .a(n_5647), .b(n_5646), .c(n_5645), .o(n_9330) );
oa12f80 g561665 ( .a(n_4837), .b(n_4836), .c(n_4835), .o(n_10729) );
ao22s80 g561666 ( .a(n_4002), .b(n_6369), .c(n_6368), .d(n_6367), .o(n_8127) );
ao12f80 g561667 ( .a(n_4866), .b(n_6366), .c(n_5431), .o(n_8087) );
oa22f80 g561668 ( .a(n_4190), .b(n_6390), .c(n_6391), .d(n_3425), .o(n_8697) );
oa12f80 g561669 ( .a(n_5594), .b(n_5593), .c(n_5592), .o(n_8619) );
in01f80 g561670 ( .a(n_7495), .o(n_7496) );
ao12f80 g561671 ( .a(n_5452), .b(n_5451), .c(n_5450), .o(n_7495) );
oa22f80 g561672 ( .a(n_6733), .b(n_4630), .c(n_4156), .d(FE_OFN646_n_6732), .o(n_8694) );
ao22s80 g561673 ( .a(n_5597), .b(n_6731), .c(n_6730), .d(n_5596), .o(n_8651) );
in01f80 g561674 ( .a(n_9793), .o(n_8222) );
ao12f80 g561675 ( .a(n_6353), .b(n_6429), .c(x_in_51_9), .o(n_9793) );
in01f80 g561676 ( .a(n_9621), .o(n_7494) );
oa12f80 g561677 ( .a(n_5575), .b(n_5574), .c(x_in_51_7), .o(n_9621) );
in01f80 g561678 ( .a(n_9787), .o(n_8221) );
ao12f80 g561679 ( .a(n_5737), .b(n_5736), .c(x_in_59_9), .o(n_9787) );
oa12f80 g561680 ( .a(n_5641), .b(n_5640), .c(n_5639), .o(n_9311) );
in01f80 g561681 ( .a(n_9247), .o(n_6729) );
ao22s80 g561682 ( .a(n_5684), .b(n_8420), .c(n_3730), .d(x_in_51_11), .o(n_9247) );
ao22s80 g561683 ( .a(n_6728), .b(n_5068), .c(n_4399), .d(n_6727), .o(n_8720) );
oa22f80 g561684 ( .a(n_3740), .b(FE_OFN309_n_3069), .c(n_1076), .d(FE_OFN129_n_27449), .o(n_7493) );
in01f80 g561685 ( .a(n_9294), .o(n_7492) );
ao22s80 g561686 ( .a(n_6402), .b(x_in_35_11), .c(n_4158), .d(n_8524), .o(n_9294) );
ao12f80 g561687 ( .a(n_5637), .b(n_6311), .c(x_in_51_13), .o(n_8648) );
ao12f80 g561688 ( .a(n_5676), .b(n_5675), .c(x_in_3_12), .o(n_9689) );
ao12f80 g561689 ( .a(n_5602), .b(n_5601), .c(x_in_51_13), .o(n_9837) );
in01f80 g561690 ( .a(n_9616), .o(n_7491) );
oa22f80 g561691 ( .a(n_3842), .b(n_6959), .c(n_6958), .d(n_3843), .o(n_9616) );
oa22f80 g561692 ( .a(n_5120), .b(n_7490), .c(n_7489), .d(n_3001), .o(n_9092) );
in01f80 g561693 ( .a(n_9296), .o(n_7488) );
oa22f80 g561694 ( .a(n_6271), .b(n_6726), .c(n_4510), .d(x_in_9_13), .o(n_9296) );
oa12f80 g561695 ( .a(n_5673), .b(n_5672), .c(x_in_59_5), .o(n_8615) );
in01f80 g561696 ( .a(n_7486), .o(n_7487) );
ao12f80 g561697 ( .a(n_4907), .b(n_4906), .c(FE_OFN1258_n_4905), .o(n_7486) );
ao22s80 g561698 ( .a(n_5662), .b(n_2105), .c(n_4932), .d(x_in_51_3), .o(n_9834) );
in01f80 g561699 ( .a(n_8812), .o(n_8813) );
ao22s80 g561700 ( .a(n_5773), .b(n_5855), .c(n_8608), .d(n_5856), .o(n_8812) );
oa22f80 g561701 ( .a(n_5662), .b(n_5980), .c(n_3874), .d(n_10817), .o(n_10714) );
in01f80 g561702 ( .a(n_10411), .o(n_8220) );
ao12f80 g561703 ( .a(n_6221), .b(n_6220), .c(n_6219), .o(n_10411) );
ao22s80 g561704 ( .a(n_6725), .b(x_in_9_13), .c(n_4681), .d(n_6726), .o(n_9208) );
in01f80 g561705 ( .a(n_10414), .o(n_10393) );
oa12f80 g561706 ( .a(n_6218), .b(n_6217), .c(n_6216), .o(n_10414) );
in01f80 g561707 ( .a(n_10407), .o(n_8219) );
oa12f80 g561708 ( .a(n_6211), .b(n_6210), .c(n_6209), .o(n_10407) );
oa22f80 g561709 ( .a(n_3483), .b(FE_OFN260_n_4280), .c(n_1057), .d(FE_OFN355_n_4860), .o(n_7485) );
in01f80 g561710 ( .a(n_8686), .o(n_7484) );
oa12f80 g561711 ( .a(n_5484), .b(n_5483), .c(n_5482), .o(n_8686) );
in01f80 g561712 ( .a(n_10391), .o(n_8218) );
oa12f80 g561713 ( .a(n_5719), .b(n_5718), .c(n_5913), .o(n_10391) );
ao12f80 g561714 ( .a(n_5553), .b(n_6011), .c(n_6724), .o(n_8699) );
in01f80 g561715 ( .a(n_8169), .o(n_9215) );
oa22f80 g561716 ( .a(n_3785), .b(n_6746), .c(n_5096), .d(x_in_3_13), .o(n_8169) );
in01f80 g561717 ( .a(n_9606), .o(n_7483) );
ao12f80 g561718 ( .a(n_5564), .b(n_5563), .c(x_in_41_15), .o(n_9606) );
oa12f80 g561719 ( .a(n_6088), .b(n_6087), .c(n_6086), .o(n_10702) );
in01f80 g561720 ( .a(n_9292), .o(n_7482) );
ao12f80 g561721 ( .a(n_5582), .b(n_5581), .c(x_in_59_12), .o(n_9292) );
in01f80 g561722 ( .a(n_10556), .o(n_10511) );
oa12f80 g561723 ( .a(n_6168), .b(n_6167), .c(FE_OFN578_n_6424), .o(n_10556) );
in01f80 g561724 ( .a(n_10350), .o(n_9459) );
oa12f80 g561725 ( .a(n_6215), .b(n_6214), .c(n_6213), .o(n_10350) );
oa22f80 g561726 ( .a(n_4535), .b(n_6723), .c(n_6722), .d(n_4397), .o(n_8622) );
oa22f80 g561727 ( .a(n_4854), .b(n_8598), .c(n_6365), .d(n_4853), .o(n_8151) );
ao12f80 g561728 ( .a(n_6283), .b(n_6282), .c(n_7481), .o(n_9011) );
ao12f80 g561729 ( .a(n_4982), .b(n_5516), .c(x_in_3_6), .o(n_9685) );
oa12f80 g561730 ( .a(n_4831), .b(n_5703), .c(x_in_25_1), .o(n_10679) );
oa22f80 g561731 ( .a(n_5080), .b(n_7480), .c(n_7479), .d(n_5185), .o(n_9067) );
ao12f80 g561732 ( .a(n_5697), .b(n_5702), .c(x_in_7_6), .o(n_6721) );
oa22f80 g561733 ( .a(n_6364), .b(n_2098), .c(n_3786), .d(n_6363), .o(n_8109) );
ao22s80 g561734 ( .a(n_4736), .b(FE_OFN674_n_6720), .c(n_6719), .d(n_2929), .o(n_8748) );
in01f80 g561735 ( .a(n_10524), .o(n_9503) );
oa12f80 g561736 ( .a(n_6085), .b(n_6084), .c(n_6083), .o(n_10524) );
ao22s80 g561737 ( .a(n_7478), .b(n_2736), .c(n_5093), .d(n_7477), .o(n_9127) );
in01f80 g561738 ( .a(n_9310), .o(n_7476) );
ao12f80 g561739 ( .a(n_5562), .b(n_5561), .c(x_in_11_12), .o(n_9310) );
in01f80 g561740 ( .a(n_9781), .o(n_8217) );
ao22s80 g561741 ( .a(n_5103), .b(n_7475), .c(n_5102), .d(n_7474), .o(n_9781) );
in01f80 g561742 ( .a(n_9333), .o(n_7473) );
ao12f80 g561743 ( .a(n_5570), .b(n_5569), .c(x_in_11_13), .o(n_9333) );
in01f80 g561744 ( .a(n_9237), .o(n_6718) );
ao22s80 g561745 ( .a(n_5301), .b(x_in_11_11), .c(n_3805), .d(n_7818), .o(n_9237) );
in01f80 g561746 ( .a(n_9326), .o(n_7472) );
ao12f80 g561747 ( .a(n_5544), .b(n_5661), .c(x_in_11_10), .o(n_9326) );
in01f80 g561748 ( .a(n_7470), .o(n_7471) );
oa22f80 g561749 ( .a(n_6717), .b(n_5571), .c(n_5572), .d(n_6716), .o(n_7470) );
in01f80 g561750 ( .a(n_9324), .o(n_7469) );
ao12f80 g561751 ( .a(n_5545), .b(n_5660), .c(x_in_11_9), .o(n_9324) );
in01f80 g561752 ( .a(n_9322), .o(n_7468) );
ao12f80 g561753 ( .a(n_5547), .b(n_5546), .c(x_in_11_8), .o(n_9322) );
oa12f80 g561754 ( .a(n_5474), .b(n_6629), .c(n_6715), .o(n_8732) );
in01f80 g561755 ( .a(n_9230), .o(n_6714) );
ao22s80 g561756 ( .a(n_5445), .b(x_in_43_12), .c(n_4072), .d(n_7263), .o(n_9230) );
ao22s80 g561757 ( .a(n_7467), .b(n_5166), .c(n_4994), .d(n_7466), .o(n_9130) );
oa12f80 g561758 ( .a(n_5543), .b(n_5542), .c(x_in_11_5), .o(n_8640) );
ao22s80 g561759 ( .a(n_3997), .b(n_6362), .c(n_6361), .d(n_6360), .o(n_8160) );
in01f80 g561760 ( .a(n_10536), .o(n_9510) );
oa12f80 g561761 ( .a(n_6080), .b(n_6079), .c(n_6078), .o(n_10536) );
oa22f80 g561762 ( .a(n_3446), .b(FE_OFN306_n_3069), .c(n_1063), .d(FE_OFN64_n_27012), .o(n_7465) );
oa12f80 g561763 ( .a(n_5472), .b(n_5471), .c(n_6713), .o(n_8738) );
in01f80 g561764 ( .a(n_9234), .o(n_6710) );
ao22s80 g561765 ( .a(n_5514), .b(n_7818), .c(n_3808), .d(x_in_11_11), .o(n_9234) );
oa12f80 g561766 ( .a(n_5473), .b(n_6005), .c(n_6709), .o(n_8735) );
oa12f80 g561767 ( .a(n_5477), .b(n_6626), .c(FE_OFN692_n_6708), .o(n_8729) );
oa22f80 g561768 ( .a(n_6789), .b(n_3266), .c(n_5073), .d(n_6788), .o(n_9172) );
oa12f80 g561769 ( .a(n_4983), .b(n_5428), .c(n_6707), .o(n_8702) );
oa12f80 g561770 ( .a(n_5651), .b(n_5650), .c(x_in_11_13), .o(n_8637) );
in01f80 g561771 ( .a(n_7463), .o(n_7464) );
oa12f80 g561772 ( .a(n_5429), .b(n_6707), .c(n_8701), .o(n_7463) );
in01f80 g561773 ( .a(n_7461), .o(n_7462) );
oa22f80 g561774 ( .a(n_4519), .b(x_in_55_12), .c(n_6395), .d(n_7278), .o(n_7461) );
in01f80 g561775 ( .a(n_9064), .o(n_10554) );
oa12f80 g561776 ( .a(n_6166), .b(n_6165), .c(n_6164), .o(n_9064) );
in01f80 g561777 ( .a(n_9250), .o(n_6706) );
ao22s80 g561778 ( .a(n_5509), .b(x_in_43_10), .c(n_3787), .d(n_6496), .o(n_9250) );
oa12f80 g561779 ( .a(n_5620), .b(n_5619), .c(x_in_5_8), .o(n_8792) );
in01f80 g561780 ( .a(n_9232), .o(n_6703) );
ao22s80 g561781 ( .a(n_5548), .b(x_in_43_13), .c(n_4058), .d(n_7274), .o(n_9232) );
in01f80 g561782 ( .a(n_9239), .o(n_6702) );
ao22s80 g561783 ( .a(n_5494), .b(x_in_43_11), .c(n_3798), .d(n_8443), .o(n_9239) );
in01f80 g561784 ( .a(n_9306), .o(n_7460) );
ao22s80 g561785 ( .a(n_4893), .b(x_in_43_9), .c(n_5500), .d(n_7268), .o(n_9306) );
ao12f80 g561786 ( .a(n_5481), .b(n_6476), .c(n_6475), .o(n_9177) );
in01f80 g561787 ( .a(n_9313), .o(n_7459) );
ao12f80 g561788 ( .a(n_5506), .b(n_5505), .c(x_in_43_8), .o(n_9313) );
in01f80 g561789 ( .a(n_9304), .o(n_7458) );
ao12f80 g561790 ( .a(n_5513), .b(n_5520), .c(x_in_43_7), .o(n_9304) );
in01f80 g561791 ( .a(n_9590), .o(n_9002) );
oa12f80 g561792 ( .a(n_5499), .b(n_5498), .c(x_in_43_6), .o(n_9590) );
ao22s80 g561793 ( .a(n_6474), .b(n_6473), .c(n_4530), .d(n_6472), .o(n_8740) );
oa12f80 g561794 ( .a(n_5541), .b(n_5540), .c(FE_OFN1184_n_6701), .o(n_8691) );
oa12f80 g561795 ( .a(n_5414), .b(FE_OFN1184_n_6701), .c(n_8690), .o(n_8782) );
in01f80 g561796 ( .a(n_9228), .o(n_6700) );
ao22s80 g561797 ( .a(n_5492), .b(n_8443), .c(n_3802), .d(x_in_43_11), .o(n_9228) );
in01f80 g561798 ( .a(n_10521), .o(n_8216) );
oa12f80 g561799 ( .a(n_6063), .b(n_6062), .c(n_6061), .o(n_10521) );
oa22f80 g561800 ( .a(n_4586), .b(n_7274), .c(n_5340), .d(x_in_43_13), .o(n_8672) );
in01f80 g561801 ( .a(n_9244), .o(n_6699) );
oa22f80 g561802 ( .a(n_3852), .b(n_8541), .c(n_5693), .d(n_6359), .o(n_9244) );
oa22f80 g561803 ( .a(n_6303), .b(n_7456), .c(n_6304), .d(n_7455), .o(n_9077) );
in01f80 g561804 ( .a(n_8112), .o(n_9241) );
oa22f80 g561805 ( .a(n_3128), .b(n_5717), .c(n_5716), .d(x_in_37_0), .o(n_8112) );
ao22s80 g561806 ( .a(n_6668), .b(n_7454), .c(n_7453), .d(n_6667), .o(n_8996) );
in01f80 g561807 ( .a(n_6697), .o(n_6698) );
oa22f80 g561808 ( .a(n_6358), .b(n_3380), .c(n_6357), .d(n_6356), .o(n_6697) );
ao12f80 g561809 ( .a(n_6235), .b(n_6234), .c(n_6478), .o(n_9097) );
oa12f80 g561810 ( .a(n_5475), .b(n_6476), .c(n_5889), .o(n_8775) );
in01f80 g561811 ( .a(n_11410), .o(n_9389) );
oa12f80 g561812 ( .a(n_7421), .b(n_7420), .c(n_7419), .o(n_11410) );
in01f80 g561813 ( .a(n_8688), .o(n_9587) );
oa12f80 g561814 ( .a(n_5531), .b(n_5530), .c(x_in_3_7), .o(n_8688) );
in01f80 g561815 ( .a(n_9217), .o(n_6696) );
oa22f80 g561816 ( .a(n_3795), .b(n_7289), .c(n_5152), .d(x_in_27_9), .o(n_9217) );
in01f80 g561817 ( .a(FE_OFN1206_n_9308), .o(n_7452) );
ao22s80 g561818 ( .a(n_6272), .b(x_in_27_8), .c(n_4546), .d(n_7287), .o(n_9308) );
in01f80 g561819 ( .a(n_9317), .o(n_7451) );
ao12f80 g561820 ( .a(n_5497), .b(n_5681), .c(x_in_27_7), .o(n_9317) );
in01f80 g561821 ( .a(n_9597), .o(n_8989) );
oa12f80 g561822 ( .a(n_5512), .b(n_5678), .c(x_in_27_6), .o(n_9597) );
in01f80 g561823 ( .a(n_8214), .o(n_8215) );
oa12f80 g561824 ( .a(n_6300), .b(n_6299), .c(x_in_27_5), .o(n_8214) );
in01f80 g561825 ( .a(n_8715), .o(n_9686) );
oa12f80 g561826 ( .a(n_5526), .b(n_5525), .c(x_in_3_9), .o(n_8715) );
ao12f80 g561827 ( .a(n_6674), .b(n_6532), .c(n_4168), .o(n_8213) );
in01f80 g561828 ( .a(n_9671), .o(n_7450) );
oa12f80 g561829 ( .a(n_5577), .b(n_5576), .c(x_in_35_12), .o(n_9671) );
in01f80 g561830 ( .a(n_9221), .o(n_6695) );
ao22s80 g561831 ( .a(n_5100), .b(x_in_27_12), .c(n_3791), .d(n_7402), .o(n_9221) );
in01f80 g561832 ( .a(n_9223), .o(n_6694) );
ao22s80 g561833 ( .a(n_5683), .b(n_8513), .c(n_3837), .d(x_in_27_11), .o(n_9223) );
in01f80 g561834 ( .a(n_9055), .o(n_10429) );
oa12f80 g561835 ( .a(n_6057), .b(n_6056), .c(n_6055), .o(n_9055) );
oa22f80 g561836 ( .a(n_5084), .b(n_6767), .c(n_6768), .d(n_4651), .o(n_8978) );
oa22f80 g561837 ( .a(n_5001), .b(n_7449), .c(n_7448), .d(n_5176), .o(n_9136) );
oa22f80 g561838 ( .a(n_4587), .b(n_7229), .c(n_5614), .d(x_in_27_13), .o(n_8625) );
oa22f80 g561839 ( .a(n_4844), .b(n_6355), .c(n_6354), .d(n_4843), .o(n_8163) );
in01f80 g561840 ( .a(n_9679), .o(n_10549) );
oa12f80 g561841 ( .a(n_5722), .b(n_5721), .c(FE_OFN991_n_5720), .o(n_9679) );
ao22s80 g561842 ( .a(n_7599), .b(n_5385), .c(n_5760), .d(n_7598), .o(n_9541) );
oa12f80 g561843 ( .a(n_6224), .b(n_6223), .c(n_7445), .o(n_8975) );
in01f80 g561844 ( .a(n_10540), .o(n_10518) );
oa12f80 g561845 ( .a(n_6183), .b(n_6182), .c(n_6181), .o(n_10540) );
oa22f80 g561846 ( .a(n_3738), .b(FE_OFN249_n_4162), .c(n_1574), .d(FE_OFN76_n_27012), .o(n_7444) );
oa22f80 g561847 ( .a(n_4935), .b(n_7443), .c(n_7442), .d(n_4923), .o(n_8972) );
in01f80 g561848 ( .a(n_10496), .o(n_8212) );
oa12f80 g561849 ( .a(n_6054), .b(n_6053), .c(n_6052), .o(n_10496) );
oa12f80 g561850 ( .a(n_5586), .b(n_5585), .c(x_in_59_10), .o(n_8643) );
oa12f80 g561851 ( .a(n_6314), .b(n_6313), .c(n_7144), .o(n_9863) );
ao22s80 g561852 ( .a(n_4407), .b(n_4088), .c(n_4406), .d(n_5717), .o(n_11440) );
in01f80 g561853 ( .a(n_7440), .o(n_7441) );
oa12f80 g561854 ( .a(n_5590), .b(n_5589), .c(n_6643), .o(n_7440) );
oa12f80 g561855 ( .a(n_5604), .b(n_5603), .c(n_6693), .o(n_10615) );
oa12f80 g561856 ( .a(n_5056), .b(n_5694), .c(x_in_1_4), .o(n_8793) );
oa22f80 g561857 ( .a(n_3759), .b(FE_OFN256_n_4280), .c(n_1562), .d(n_29617), .o(n_6692) );
oa22f80 g561858 ( .a(n_5022), .b(FE_OFN256_n_4280), .c(n_555), .d(FE_OFN1108_rst), .o(n_7439) );
oa22f80 g561859 ( .a(FE_OFN827_n_3772), .b(n_29046), .c(n_411), .d(FE_OFN326_n_4860), .o(n_7416) );
oa22f80 g561860 ( .a(n_3748), .b(FE_OFN187_n_29496), .c(n_1600), .d(FE_OFN15_n_29068), .o(n_6691) );
oa22f80 g561861 ( .a(n_7218), .b(FE_OFN303_n_3069), .c(n_1485), .d(n_27709), .o(n_7438) );
oa22f80 g561862 ( .a(n_6297), .b(FE_OFN309_n_3069), .c(n_682), .d(FE_OFN69_n_27012), .o(n_7437) );
ao22s80 g561863 ( .a(n_6295), .b(n_6689), .c(n_6530), .d(n_4389), .o(n_6690) );
ao22s80 g561864 ( .a(n_6293), .b(n_6687), .c(n_6528), .d(n_6013), .o(n_6688) );
ao22s80 g561865 ( .a(n_6294), .b(n_6711), .c(n_4921), .d(n_4469), .o(n_6712) );
ao22s80 g561866 ( .a(n_5711), .b(n_6685), .c(n_6524), .d(n_4224), .o(n_6686) );
ao22s80 g561867 ( .a(n_5712), .b(n_6683), .c(n_6526), .d(n_4548), .o(n_6684) );
ao22s80 g561868 ( .a(n_6291), .b(n_6483), .c(n_6522), .d(n_6015), .o(n_6682) );
in01f80 g561869 ( .a(n_9703), .o(n_8211) );
ao22s80 g561870 ( .a(n_7217), .b(x_in_45_13), .c(n_5094), .d(n_7216), .o(n_9703) );
in01f80 g561871 ( .a(n_9254), .o(n_6681) );
ao22s80 g561872 ( .a(n_5668), .b(x_in_51_11), .c(n_4039), .d(n_8420), .o(n_9254) );
oa22f80 g561873 ( .a(n_6042), .b(n_8929), .c(n_3836), .d(x_in_61_4), .o(n_8143) );
ao22s80 g561874 ( .a(n_4729), .b(x_in_33_11), .c(n_6680), .d(n_12178), .o(n_8743) );
oa22f80 g561875 ( .a(n_6044), .b(n_8522), .c(n_3375), .d(x_in_7_4), .o(n_8093) );
in01f80 g561876 ( .a(n_9298), .o(n_7436) );
ao22s80 g561877 ( .a(n_4536), .b(n_8482), .c(n_5746), .d(x_in_59_11), .o(n_9298) );
ao22s80 g561878 ( .a(n_3846), .b(x_in_33_12), .c(n_5440), .d(n_12635), .o(n_8115) );
in01f80 g561879 ( .a(n_9660), .o(n_7644) );
oa22f80 g561880 ( .a(n_5741), .b(x_in_35_11), .c(n_4387), .d(n_8524), .o(n_9660) );
in01f80 g561881 ( .a(n_8209), .o(n_8210) );
oa22f80 g561882 ( .a(n_7435), .b(n_7434), .c(n_5097), .d(x_in_21_2), .o(n_8209) );
ao22s80 g561883 ( .a(n_3826), .b(x_in_33_6), .c(n_6352), .d(n_12172), .o(n_8174) );
in01f80 g561884 ( .a(n_9252), .o(n_6679) );
ao22s80 g561885 ( .a(n_4995), .b(x_in_51_10), .c(n_3851), .d(n_5283), .o(n_9252) );
in01f80 g561886 ( .a(n_9245), .o(n_7040) );
oa22f80 g561887 ( .a(n_3850), .b(n_6351), .c(n_5638), .d(x_in_51_8), .o(n_9245) );
ao22s80 g561888 ( .a(n_5652), .b(x_in_51_6), .c(n_3865), .d(n_6350), .o(n_8479) );
ao22s80 g561889 ( .a(n_3812), .b(x_in_33_10), .c(n_6349), .d(n_12634), .o(n_8183) );
ao22s80 g561890 ( .a(n_4054), .b(x_in_33_9), .c(n_6348), .d(n_8884), .o(n_8745) );
ao22s80 g561891 ( .a(n_3519), .b(x_in_33_8), .c(n_6347), .d(n_12175), .o(n_8180) );
ao22s80 g561892 ( .a(n_3813), .b(x_in_33_7), .c(n_6346), .d(n_8885), .o(n_8177) );
ao22s80 g561893 ( .a(n_6345), .b(n_5653), .c(n_6344), .d(n_5654), .o(n_8101) );
ao22s80 g561894 ( .a(n_4543), .b(x_in_33_4), .c(n_7201), .d(n_5281), .o(n_8751) );
in01f80 g561895 ( .a(n_9256), .o(n_6678) );
ao22s80 g561896 ( .a(n_5067), .b(x_in_51_12), .c(n_3484), .d(n_6420), .o(n_9256) );
in01f80 g561897 ( .a(n_9619), .o(n_7433) );
ao12f80 g561898 ( .a(n_4764), .b(n_10948), .c(n_5925), .o(n_9619) );
in01f80 g561899 ( .a(n_9213), .o(n_7202) );
ao22s80 g561900 ( .a(n_5692), .b(x_in_59_8), .c(n_3995), .d(n_5691), .o(n_9213) );
in01f80 g561901 ( .a(n_9264), .o(n_6677) );
ao22s80 g561902 ( .a(n_4961), .b(x_in_19_7), .c(n_3735), .d(n_5940), .o(n_9264) );
in01f80 g561903 ( .a(n_9259), .o(n_6676) );
oa22f80 g561904 ( .a(n_3892), .b(n_5689), .c(n_5690), .d(x_in_51_13), .o(n_9259) );
in01f80 g561905 ( .a(n_7431), .o(n_7432) );
ao22s80 g561906 ( .a(n_4303), .b(x_in_13_12), .c(n_4304), .d(n_5926), .o(n_7431) );
ao22s80 g561907 ( .a(n_3816), .b(x_in_33_5), .c(n_6343), .d(n_11297), .o(n_8186) );
in01f80 g561908 ( .a(n_9281), .o(n_6675) );
ao22s80 g561909 ( .a(n_5591), .b(x_in_59_7), .c(n_3733), .d(n_5699), .o(n_9281) );
oa22f80 g561910 ( .a(n_6342), .b(n_3369), .c(n_6341), .d(n_3856), .o(n_8097) );
ao22s80 g561911 ( .a(n_6340), .b(n_5656), .c(n_6339), .d(n_5657), .o(n_8629) );
oa22f80 g561912 ( .a(n_6450), .b(n_3840), .c(n_6449), .d(n_3857), .o(n_8129) );
oa22f80 g561913 ( .a(n_6338), .b(n_6337), .c(n_6336), .d(n_3906), .o(n_8099) );
ao22s80 g561914 ( .a(n_7430), .b(n_7209), .c(n_7429), .d(n_7208), .o(n_8998) );
ao22s80 g561915 ( .a(n_6335), .b(n_3877), .c(n_6334), .d(n_6333), .o(n_8095) );
ao22s80 g561916 ( .a(n_5183), .b(n_7793), .c(n_5852), .d(n_7653), .o(n_9117) );
oa22f80 g561917 ( .a(n_4830), .b(n_3074), .c(n_3858), .d(n_4018), .o(n_8801) );
no02f80 g561918 ( .a(n_6366), .b(n_5431), .o(n_4866) );
na02f80 g561919 ( .a(n_6047), .b(n_6387), .o(n_4865) );
na02f80 g561920 ( .a(n_6389), .b(n_4740), .o(n_4380) );
na02f80 g561921 ( .a(n_5657), .b(n_5656), .o(n_5658) );
no02f80 g561922 ( .a(n_6673), .b(x_in_39_6), .o(n_6674) );
na02f80 g561923 ( .a(n_5654), .b(n_5653), .o(n_5655) );
na02f80 g561924 ( .a(n_12281), .b(n_14115), .o(n_8387) );
na02f80 g561925 ( .a(n_5202), .b(n_6671), .o(n_6672) );
in01f80 g561926 ( .a(n_6332), .o(n_10316) );
no02f80 g561927 ( .a(n_5067), .b(n_6420), .o(n_6332) );
in01f80 g561928 ( .a(n_6331), .o(n_11367) );
no02f80 g561929 ( .a(n_5652), .b(n_6350), .o(n_6331) );
no02f80 g561930 ( .a(n_6449), .b(n_6450), .o(n_4864) );
no02f80 g561931 ( .a(n_10983), .b(n_13232), .o(n_7169) );
na02f80 g561932 ( .a(n_5106), .b(n_6038), .o(n_6670) );
no02f80 g561933 ( .a(n_3171), .b(n_4601), .o(n_6417) );
oa12f80 g561934 ( .a(n_5105), .b(n_6330), .c(n_1995), .o(n_13306) );
na02f80 g561935 ( .a(n_5650), .b(x_in_11_13), .o(n_5651) );
na02f80 g561936 ( .a(n_5649), .b(x_in_4_2), .o(n_7972) );
in01f80 g561937 ( .a(n_6328), .o(n_6329) );
no02f80 g561938 ( .a(n_5649), .b(x_in_4_2), .o(n_6328) );
oa12f80 g561939 ( .a(n_4863), .b(n_4862), .c(n_1981), .o(n_10975) );
no02f80 g561940 ( .a(n_6341), .b(n_6342), .o(n_4880) );
na02f80 g561941 ( .a(n_7209), .b(n_7208), .o(n_7210) );
na02f80 g561942 ( .a(n_5694), .b(x_in_1_4), .o(n_5056) );
na02f80 g561943 ( .a(n_6371), .b(n_5832), .o(n_5648) );
na02f80 g561944 ( .a(n_5646), .b(n_5645), .o(n_5647) );
na02f80 g561945 ( .a(n_4949), .b(x_in_0_2), .o(n_7976) );
in01f80 g561946 ( .a(n_6432), .o(n_6433) );
no02f80 g561947 ( .a(n_4949), .b(x_in_0_2), .o(n_6432) );
no02f80 g561948 ( .a(n_4861), .b(n_9034), .o(n_7953) );
na02f80 g561949 ( .a(n_5643), .b(n_5642), .o(n_5644) );
na02f80 g561950 ( .a(n_5640), .b(n_5639), .o(n_5641) );
no02f80 g561951 ( .a(n_11609), .b(n_5101), .o(n_7929) );
in01f80 g561952 ( .a(n_6327), .o(n_10311) );
no02f80 g561953 ( .a(n_4995), .b(n_5283), .o(n_6327) );
in01f80 g561954 ( .a(n_6436), .o(n_12111) );
no02f80 g561955 ( .a(n_5638), .b(n_6351), .o(n_6436) );
na02f80 g561956 ( .a(n_4826), .b(n_4327), .o(n_4328) );
na02f80 g561957 ( .a(n_8195), .b(n_6325), .o(n_6326) );
na02f80 g561958 ( .a(n_5686), .b(n_5685), .o(n_5687) );
in01f80 g561959 ( .a(n_6323), .o(n_6324) );
na02f80 g561960 ( .a(n_4769), .b(n_5688), .o(n_6323) );
in01f80 g561961 ( .a(n_6322), .o(n_10308) );
no02f80 g561962 ( .a(n_5690), .b(n_5689), .o(n_6322) );
no02f80 g561963 ( .a(n_6311), .b(x_in_51_13), .o(n_5637) );
na02f80 g561964 ( .a(n_4680), .b(n_5006), .o(n_8385) );
in01f80 g561965 ( .a(n_6321), .o(n_7909) );
na02f80 g561966 ( .a(n_5694), .b(n_247), .o(n_6321) );
in01f80 g561967 ( .a(n_5921), .o(n_10305) );
no02f80 g561968 ( .a(n_5668), .b(n_8420), .o(n_5921) );
in01f80 g561969 ( .a(n_6320), .o(n_12107) );
no02f80 g561970 ( .a(n_5692), .b(n_5691), .o(n_6320) );
na02f80 g561971 ( .a(n_5635), .b(n_5916), .o(n_5636) );
no02f80 g561972 ( .a(n_5778), .b(n_5777), .o(n_5779) );
na02f80 g561973 ( .a(n_6318), .b(n_6317), .o(n_6319) );
in01f80 g561974 ( .a(n_6316), .o(n_8478) );
no02f80 g561975 ( .a(n_5693), .b(n_8541), .o(n_6316) );
na02f80 g561976 ( .a(n_4009), .b(n_5695), .o(n_5696) );
in01f80 g561977 ( .a(n_8391), .o(n_7426) );
na02f80 g561978 ( .a(n_6673), .b(n_6500), .o(n_8391) );
na02f80 g561979 ( .a(n_4010), .b(n_5633), .o(n_5634) );
no02f80 g561980 ( .a(n_5702), .b(x_in_7_6), .o(n_5697) );
no02f80 g561981 ( .a(n_6447), .b(x_in_35_13), .o(n_5632) );
no02f80 g561982 ( .a(n_4858), .b(n_4857), .o(n_4859) );
no02f80 g561983 ( .a(n_6388), .b(n_5695), .o(n_4856) );
no02f80 g561984 ( .a(n_6379), .b(n_5633), .o(n_4889) );
na02f80 g561985 ( .a(n_7889), .b(n_10894), .o(n_5631) );
no02f80 g561986 ( .a(n_7889), .b(n_10894), .o(n_5630) );
na02f80 g561987 ( .a(n_5650), .b(n_8636), .o(n_4993) );
no02f80 g561988 ( .a(n_7891), .b(n_10889), .o(n_5629) );
na02f80 g561989 ( .a(n_7891), .b(n_10889), .o(n_5628) );
no02f80 g561990 ( .a(n_4854), .b(n_4853), .o(n_4855) );
na02f80 g561991 ( .a(n_5626), .b(n_8655), .o(n_5627) );
na02f80 g561992 ( .a(n_6313), .b(n_7144), .o(n_6314) );
na02f80 g561993 ( .a(n_6311), .b(n_4840), .o(n_6312) );
na02f80 g561994 ( .a(n_6441), .b(n_3149), .o(n_6442) );
na02f80 g561995 ( .a(n_5624), .b(x_in_59_13), .o(n_5625) );
no02f80 g561996 ( .a(n_4999), .b(n_4998), .o(n_5000) );
in01f80 g561997 ( .a(n_7422), .o(n_7423) );
no02f80 g561998 ( .a(n_5114), .b(n_7215), .o(n_7422) );
no02f80 g561999 ( .a(n_4850), .b(x_in_61_2), .o(n_4851) );
na02f80 g562000 ( .a(n_4848), .b(x_in_61_14), .o(n_4849) );
in01f80 g562001 ( .a(n_6468), .o(n_6469) );
na02f80 g562002 ( .a(n_6443), .b(n_3148), .o(n_6468) );
no02f80 g562003 ( .a(n_5622), .b(FE_OFN458_n_5621), .o(n_5623) );
na02f80 g562004 ( .a(n_6308), .b(n_6307), .o(n_6309) );
na02f80 g562005 ( .a(n_5619), .b(x_in_5_8), .o(n_5620) );
no02f80 g562006 ( .a(n_5617), .b(n_5616), .o(n_5618) );
na02f80 g562007 ( .a(n_5614), .b(n_8624), .o(n_5615) );
no02f80 g562008 ( .a(n_5612), .b(n_5611), .o(n_5613) );
na02f80 g562009 ( .a(n_5340), .b(n_8671), .o(n_5341) );
na02f80 g562010 ( .a(n_6447), .b(n_4381), .o(n_6448) );
na02f80 g562011 ( .a(n_5769), .b(x_in_61_13), .o(n_5610) );
no02f80 g562012 ( .a(n_4974), .b(x_in_27_7), .o(n_4975) );
in01f80 g562013 ( .a(n_9409), .o(n_8840) );
no02f80 g562014 ( .a(n_7217), .b(n_7216), .o(n_9409) );
no02f80 g562015 ( .a(n_5608), .b(x_in_43_8), .o(n_5609) );
in01f80 g562016 ( .a(n_6511), .o(n_6306) );
na02f80 g562017 ( .a(n_5702), .b(n_5968), .o(n_6511) );
no02f80 g562018 ( .a(n_5606), .b(x_in_35_7), .o(n_5607) );
in01f80 g562019 ( .a(n_8461), .o(n_8463) );
no02f80 g562020 ( .a(n_32742), .b(n_2938), .o(n_8461) );
no02f80 g562021 ( .a(n_6304), .b(n_6303), .o(n_6305) );
ao12f80 g562022 ( .a(n_3199), .b(n_5325), .c(x_in_51_11), .o(n_8476) );
in01f80 g562023 ( .a(n_6301), .o(n_6302) );
no02f80 g562024 ( .a(n_3395), .b(n_5605), .o(n_6301) );
na02f80 g562025 ( .a(n_6299), .b(x_in_27_5), .o(n_6300) );
na02f80 g562026 ( .a(n_5603), .b(n_6693), .o(n_5604) );
no02f80 g562027 ( .a(n_5601), .b(x_in_51_13), .o(n_5602) );
no02f80 g562028 ( .a(n_5708), .b(FE_OFN765_n_5707), .o(n_5709) );
in01f80 g562029 ( .a(n_10869), .o(n_5600) );
na02f80 g562030 ( .a(n_4850), .b(n_4143), .o(n_10869) );
ao12f80 g562031 ( .a(n_2695), .b(n_4927), .c(x_in_51_9), .o(n_8471) );
no02f80 g562032 ( .a(n_6297), .b(n_6296), .o(n_6298) );
in01f80 g562033 ( .a(n_7220), .o(n_8843) );
no02f80 g562034 ( .a(n_6451), .b(n_6296), .o(n_7220) );
na02f80 g562035 ( .a(n_3243), .b(n_3342), .o(n_8192) );
na02f80 g562036 ( .a(n_4848), .b(n_4847), .o(n_11335) );
na02f80 g562037 ( .a(n_6668), .b(n_6667), .o(n_6669) );
in01f80 g562038 ( .a(n_8434), .o(n_6666) );
no02f80 g562039 ( .a(n_6295), .b(x_in_23_6), .o(n_8434) );
in01f80 g562040 ( .a(n_8436), .o(n_6665) );
no02f80 g562041 ( .a(n_5711), .b(x_in_55_6), .o(n_8436) );
in01f80 g562042 ( .a(n_8426), .o(n_6664) );
no02f80 g562043 ( .a(n_6294), .b(x_in_63_6), .o(n_8426) );
in01f80 g562044 ( .a(n_8432), .o(n_6663) );
no02f80 g562045 ( .a(n_6293), .b(x_in_15_6), .o(n_8432) );
na02f80 g562046 ( .a(n_19015), .b(n_4585), .o(n_6292) );
na02f80 g562047 ( .a(n_5597), .b(n_5596), .o(n_5598) );
in01f80 g562048 ( .a(n_8810), .o(n_7199) );
na02f80 g562049 ( .a(n_3190), .b(n_4846), .o(n_8810) );
na02f80 g562050 ( .a(n_2770), .b(n_4846), .o(n_9185) );
in01f80 g562051 ( .a(n_8430), .o(n_6662) );
no02f80 g562052 ( .a(n_5712), .b(x_in_47_6), .o(n_8430) );
in01f80 g562053 ( .a(n_8428), .o(n_6661) );
no02f80 g562054 ( .a(n_6291), .b(x_in_31_6), .o(n_8428) );
na02f80 g562055 ( .a(n_5624), .b(n_8682), .o(n_5595) );
in01f80 g562056 ( .a(n_8474), .o(n_6290) );
no02f80 g562057 ( .a(n_32736), .b(n_3314), .o(n_8474) );
na02f80 g562058 ( .a(n_7420), .b(n_7419), .o(n_7421) );
no02f80 g562059 ( .a(n_5437), .b(x_in_35_13), .o(n_4996) );
na02f80 g562060 ( .a(n_6288), .b(n_4878), .o(n_6289) );
ao12f80 g562061 ( .a(n_3212), .b(n_4936), .c(x_in_51_7), .o(n_8466) );
no02f80 g562062 ( .a(n_6286), .b(n_6285), .o(n_6287) );
na02f80 g562063 ( .a(n_6719), .b(FE_OFN674_n_6720), .o(n_4917) );
na02f80 g562064 ( .a(n_5593), .b(n_5592), .o(n_5594) );
in01f80 g562065 ( .a(n_5731), .o(n_11343) );
no02f80 g562066 ( .a(n_4961), .b(n_5940), .o(n_5731) );
in01f80 g562067 ( .a(n_6284), .o(n_10302) );
no02f80 g562068 ( .a(n_5591), .b(n_5699), .o(n_6284) );
na02f80 g562069 ( .a(n_2833), .b(n_4151), .o(n_8781) );
na02f80 g562070 ( .a(n_4912), .b(n_4911), .o(n_4913) );
no02f80 g562071 ( .a(n_6660), .b(x_in_38_1), .o(n_8944) );
na02f80 g562072 ( .a(n_6660), .b(x_in_38_1), .o(n_8945) );
in01f80 g562073 ( .a(n_6658), .o(n_6659) );
na02f80 g562074 ( .a(n_13246), .b(n_8438), .o(n_6658) );
in01f80 g562075 ( .a(n_6656), .o(n_6657) );
no02f80 g562076 ( .a(n_13246), .b(n_8438), .o(n_6656) );
no02f80 g562077 ( .a(n_6461), .b(n_4029), .o(n_13490) );
na02f80 g562078 ( .a(n_5589), .b(n_6643), .o(n_5590) );
no02f80 g562079 ( .a(n_4844), .b(n_4843), .o(n_4845) );
no02f80 g562080 ( .a(n_6282), .b(n_7481), .o(n_6283) );
no02f80 g562081 ( .a(n_5736), .b(x_in_59_9), .o(n_5737) );
na02f80 g562082 ( .a(n_5587), .b(x_in_35_8), .o(n_5588) );
na02f80 g562083 ( .a(n_6030), .b(x_in_3_4), .o(n_10909) );
in01f80 g562084 ( .a(n_7112), .o(n_6281) );
na02f80 g562085 ( .a(n_4974), .b(n_5680), .o(n_7112) );
na02f80 g562086 ( .a(n_5585), .b(x_in_59_10), .o(n_5586) );
na02f80 g562087 ( .a(n_5583), .b(x_in_59_13), .o(n_5584) );
in01f80 g562088 ( .a(n_7105), .o(n_6280) );
na02f80 g562089 ( .a(n_5619), .b(n_5291), .o(n_7105) );
no02f80 g562090 ( .a(n_6278), .b(x_in_59_14), .o(n_6279) );
no02f80 g562091 ( .a(n_5734), .b(n_6641), .o(n_5735) );
na02f80 g562092 ( .a(n_6014), .b(x_in_3_8), .o(n_10905) );
no02f80 g562093 ( .a(n_5581), .b(x_in_59_12), .o(n_5582) );
ao12f80 g562094 ( .a(n_3198), .b(n_4841), .c(x_in_51_12), .o(n_8512) );
no02f80 g562095 ( .a(n_5663), .b(x_in_35_10), .o(n_5237) );
no02f80 g562096 ( .a(n_6276), .b(n_7551), .o(n_6277) );
in01f80 g562097 ( .a(n_7930), .o(n_8845) );
na02f80 g562098 ( .a(n_5741), .b(n_8524), .o(n_7930) );
in01f80 g562099 ( .a(n_7095), .o(n_5744) );
na02f80 g562100 ( .a(n_5608), .b(n_5501), .o(n_7095) );
na02f80 g562101 ( .a(n_6010), .b(x_in_3_6), .o(n_10900) );
no02f80 g562102 ( .a(n_6364), .b(n_6363), .o(n_4839) );
in01f80 g562103 ( .a(n_7880), .o(n_8849) );
na02f80 g562104 ( .a(n_5746), .b(n_8482), .o(n_7880) );
na02f80 g562105 ( .a(n_5579), .b(x_in_35_13), .o(n_5580) );
no02f80 g562106 ( .a(n_6725), .b(n_9207), .o(n_5578) );
no02f80 g562107 ( .a(n_6654), .b(n_6653), .o(n_6655) );
na02f80 g562108 ( .a(n_7555), .b(n_7554), .o(n_6467) );
na02f80 g562109 ( .a(n_5576), .b(x_in_35_12), .o(n_5577) );
no02f80 g562110 ( .a(n_5516), .b(x_in_3_6), .o(n_4982) );
na02f80 g562111 ( .a(n_5769), .b(n_9334), .o(n_5770) );
na02f80 g562112 ( .a(n_5428), .b(n_6707), .o(n_4983) );
in01f80 g562113 ( .a(n_11245), .o(n_6275) );
no02f80 g562114 ( .a(n_5606), .b(n_4942), .o(n_11245) );
na02f80 g562115 ( .a(n_5574), .b(x_in_51_7), .o(n_5575) );
na02f80 g562116 ( .a(n_3194), .b(n_3052), .o(n_8778) );
na02f80 g562117 ( .a(n_5572), .b(n_5571), .o(n_5573) );
na02f80 g562118 ( .a(n_6652), .b(n_4990), .o(n_8398) );
in01f80 g562119 ( .a(n_6274), .o(n_10296) );
no02f80 g562120 ( .a(n_5535), .b(n_5326), .o(n_6274) );
no02f80 g562121 ( .a(n_5569), .b(x_in_11_13), .o(n_5570) );
in01f80 g562122 ( .a(n_6273), .o(n_10293) );
no02f80 g562123 ( .a(n_5569), .b(n_2681), .o(n_6273) );
na02f80 g562124 ( .a(n_6001), .b(x_in_3_10), .o(n_10875) );
na02f80 g562125 ( .a(n_3817), .b(n_5567), .o(n_5568) );
in01f80 g562126 ( .a(n_10576), .o(n_6618) );
no02f80 g562127 ( .a(n_6272), .b(n_7287), .o(n_10576) );
no02f80 g562128 ( .a(n_6381), .b(n_5567), .o(n_4838) );
na02f80 g562129 ( .a(n_5565), .b(x_in_35_9), .o(n_5566) );
na02f80 g562130 ( .a(n_4836), .b(n_4835), .o(n_4837) );
no02f80 g562131 ( .a(n_5563), .b(x_in_41_15), .o(n_5564) );
no02f80 g562132 ( .a(n_6429), .b(x_in_51_9), .o(n_6353) );
in01f80 g562133 ( .a(n_11206), .o(n_6041) );
no02f80 g562134 ( .a(n_5437), .b(n_5245), .o(n_11206) );
na02f80 g562135 ( .a(n_6271), .b(x_in_9_13), .o(n_7736) );
no02f80 g562136 ( .a(n_5561), .b(x_in_11_12), .o(n_5562) );
in01f80 g562137 ( .a(n_6270), .o(n_11323) );
no02f80 g562138 ( .a(n_5561), .b(n_5025), .o(n_6270) );
na02f80 g562139 ( .a(n_5559), .b(n_5558), .o(n_5560) );
in01f80 g562140 ( .a(n_6160), .o(n_10288) );
no02f80 g562141 ( .a(n_5557), .b(n_5556), .o(n_6160) );
in01f80 g562142 ( .a(n_6269), .o(n_11317) );
no02f80 g562143 ( .a(n_5555), .b(n_5554), .o(n_6269) );
in01f80 g562144 ( .a(n_6268), .o(n_11209) );
no02f80 g562145 ( .a(n_5583), .b(n_2635), .o(n_6268) );
no02f80 g562146 ( .a(n_5538), .b(x_in_19_9), .o(n_5254) );
no02f80 g562147 ( .a(n_6011), .b(n_6724), .o(n_5553) );
na02f80 g562148 ( .a(n_5551), .b(x_in_11_6), .o(n_5552) );
in01f80 g562149 ( .a(n_6267), .o(n_10279) );
no02f80 g562150 ( .a(n_5502), .b(n_7229), .o(n_6267) );
no02f80 g562151 ( .a(n_5549), .b(x_in_11_7), .o(n_5550) );
in01f80 g562152 ( .a(n_6310), .o(n_10282) );
no02f80 g562153 ( .a(n_5548), .b(n_7274), .o(n_6310) );
no02f80 g562154 ( .a(n_5546), .b(x_in_11_8), .o(n_5547) );
no02f80 g562155 ( .a(n_5660), .b(x_in_11_9), .o(n_5545) );
in01f80 g562156 ( .a(n_6266), .o(n_10285) );
no02f80 g562157 ( .a(n_5661), .b(n_3229), .o(n_6266) );
in01f80 g562158 ( .a(n_6265), .o(n_11311) );
no02f80 g562159 ( .a(n_5660), .b(n_5310), .o(n_6265) );
in01f80 g562160 ( .a(n_6264), .o(n_11314) );
no02f80 g562161 ( .a(n_5546), .b(n_5352), .o(n_6264) );
in01f80 g562162 ( .a(n_6263), .o(n_11308) );
no02f80 g562163 ( .a(n_5549), .b(n_5089), .o(n_6263) );
in01f80 g562164 ( .a(n_6262), .o(n_11305) );
no02f80 g562165 ( .a(n_5551), .b(n_5309), .o(n_6262) );
no02f80 g562166 ( .a(n_5661), .b(x_in_11_10), .o(n_5544) );
no02f80 g562167 ( .a(n_6651), .b(n_5786), .o(n_19669) );
no02f80 g562168 ( .a(n_5557), .b(x_in_19_13), .o(n_5343) );
na02f80 g562169 ( .a(n_5542), .b(x_in_11_5), .o(n_5543) );
na02f80 g562170 ( .a(n_5540), .b(FE_OFN1184_n_6701), .o(n_5541) );
no02f80 g562171 ( .a(n_5664), .b(x_in_19_10), .o(n_5539) );
in01f80 g562172 ( .a(n_11182), .o(n_6370) );
no02f80 g562173 ( .a(n_5587), .b(n_4939), .o(n_11182) );
na02f80 g562174 ( .a(n_10765), .b(n_7835), .o(n_6261) );
no02f80 g562175 ( .a(n_10765), .b(n_7835), .o(n_6260) );
in01f80 g562176 ( .a(n_6259), .o(n_11189) );
no02f80 g562177 ( .a(n_5663), .b(n_2652), .o(n_6259) );
in01f80 g562178 ( .a(n_6258), .o(n_11285) );
no02f80 g562179 ( .a(n_5664), .b(n_3020), .o(n_6258) );
in01f80 g562180 ( .a(n_6257), .o(n_11255) );
no02f80 g562181 ( .a(n_5538), .b(n_5537), .o(n_6257) );
no02f80 g562182 ( .a(n_5535), .b(x_in_19_6), .o(n_5536) );
in01f80 g562183 ( .a(n_6256), .o(n_10276) );
no02f80 g562184 ( .a(n_5445), .b(n_7263), .o(n_6256) );
no02f80 g562185 ( .a(n_5555), .b(x_in_19_8), .o(n_5534) );
no02f80 g562186 ( .a(n_5670), .b(x_in_43_5), .o(n_5671) );
in01f80 g562187 ( .a(n_6255), .o(n_10273) );
no02f80 g562188 ( .a(n_5100), .b(n_7402), .o(n_6255) );
in01f80 g562189 ( .a(n_11176), .o(n_6254) );
no02f80 g562190 ( .a(n_5585), .b(n_2668), .o(n_11176) );
na02f80 g562191 ( .a(n_4805), .b(x_in_59_9), .o(n_11094) );
no02f80 g562192 ( .a(n_5532), .b(x_in_59_6), .o(n_5533) );
na02f80 g562193 ( .a(n_5530), .b(x_in_3_7), .o(n_5531) );
no02f80 g562194 ( .a(n_5528), .b(x_in_3_8), .o(n_5529) );
in01f80 g562195 ( .a(n_6253), .o(n_10264) );
no02f80 g562196 ( .a(n_5667), .b(n_5666), .o(n_6253) );
in01f80 g562197 ( .a(n_11192), .o(n_6650) );
no02f80 g562198 ( .a(n_6402), .b(n_8524), .o(n_11192) );
no02f80 g562199 ( .a(n_5667), .b(x_in_3_10), .o(n_5527) );
na02f80 g562200 ( .a(n_5525), .b(x_in_3_9), .o(n_5526) );
na02f80 g562201 ( .a(n_3783), .b(x_in_3_7), .o(n_11282) );
in01f80 g562202 ( .a(n_6252), .o(n_11291) );
no02f80 g562203 ( .a(n_5528), .b(n_5524), .o(n_6252) );
na02f80 g562204 ( .a(n_5672), .b(x_in_59_5), .o(n_5673) );
no02f80 g562205 ( .a(n_4873), .b(x_in_25_4), .o(n_9956) );
in01f80 g562206 ( .a(n_6251), .o(n_11288) );
no02f80 g562207 ( .a(n_5659), .b(n_5369), .o(n_6251) );
no02f80 g562208 ( .a(n_5659), .b(x_in_35_6), .o(n_5523) );
na02f80 g562209 ( .a(n_5521), .b(x_in_19_5), .o(n_5522) );
in01f80 g562210 ( .a(n_6250), .o(n_11294) );
no02f80 g562211 ( .a(n_5520), .b(n_5519), .o(n_6250) );
in01f80 g562212 ( .a(n_6426), .o(n_11220) );
no02f80 g562213 ( .a(n_5565), .b(n_5098), .o(n_6426) );
na02f80 g562214 ( .a(n_5517), .b(x_in_25_4), .o(n_5518) );
in01f80 g562215 ( .a(n_6249), .o(n_11378) );
no02f80 g562216 ( .a(n_5516), .b(n_5515), .o(n_6249) );
in01f80 g562217 ( .a(n_6419), .o(n_11279) );
no02f80 g562218 ( .a(n_5301), .b(n_7818), .o(n_6419) );
no02f80 g562219 ( .a(n_5675), .b(x_in_3_12), .o(n_5676) );
in01f80 g562220 ( .a(n_7003), .o(n_8450) );
no02f80 g562221 ( .a(n_5514), .b(x_in_11_11), .o(n_7003) );
in01f80 g562222 ( .a(n_6248), .o(n_10267) );
no02f80 g562223 ( .a(n_5532), .b(n_5275), .o(n_6248) );
no02f80 g562224 ( .a(n_5520), .b(x_in_43_7), .o(n_5513) );
in01f80 g562225 ( .a(n_6247), .o(n_11276) );
no02f80 g562226 ( .a(n_5678), .b(n_5677), .o(n_6247) );
na02f80 g562227 ( .a(n_5678), .b(x_in_27_6), .o(n_5512) );
na02f80 g562228 ( .a(n_3750), .b(x_in_3_9), .o(n_11273) );
in01f80 g562229 ( .a(n_6246), .o(n_10270) );
no02f80 g562230 ( .a(n_5675), .b(n_5247), .o(n_6246) );
in01f80 g562231 ( .a(n_6245), .o(n_11097) );
no02f80 g562232 ( .a(n_5581), .b(n_4992), .o(n_6245) );
in01f80 g562233 ( .a(n_6421), .o(n_11267) );
no02f80 g562234 ( .a(n_5498), .b(n_5327), .o(n_6421) );
no02f80 g562235 ( .a(n_5510), .b(x_in_3_5), .o(n_5511) );
in01f80 g562236 ( .a(n_6244), .o(n_10261) );
no02f80 g562237 ( .a(n_5509), .b(n_6496), .o(n_6244) );
no02f80 g562238 ( .a(n_5507), .b(x_in_35_5), .o(n_5508) );
in01f80 g562239 ( .a(n_6243), .o(n_10255) );
no02f80 g562240 ( .a(n_5152), .b(n_7289), .o(n_6243) );
no02f80 g562241 ( .a(n_5505), .b(x_in_43_8), .o(n_5506) );
na02f80 g562242 ( .a(n_5503), .b(x_in_59_3), .o(n_5504) );
in01f80 g562243 ( .a(n_6242), .o(n_10258) );
no02f80 g562244 ( .a(n_5065), .b(n_7417), .o(n_6242) );
na02f80 g562245 ( .a(n_4215), .b(x_in_35_13), .o(n_9868) );
in01f80 g562246 ( .a(n_6241), .o(n_11270) );
no02f80 g562247 ( .a(n_5505), .b(n_5501), .o(n_6241) );
in01f80 g562248 ( .a(n_6240), .o(n_11179) );
no02f80 g562249 ( .a(n_5576), .b(n_5032), .o(n_6240) );
in01f80 g562250 ( .a(n_10239), .o(n_6239) );
na02f80 g562251 ( .a(n_5500), .b(x_in_43_9), .o(n_10239) );
na02f80 g562252 ( .a(n_5498), .b(x_in_43_6), .o(n_5499) );
in01f80 g562253 ( .a(n_6238), .o(n_11264) );
no02f80 g562254 ( .a(n_5681), .b(n_5680), .o(n_6238) );
no02f80 g562255 ( .a(n_5681), .b(x_in_27_7), .o(n_5497) );
in01f80 g562256 ( .a(n_11186), .o(n_6237) );
no02f80 g562257 ( .a(n_5496), .b(n_8482), .o(n_11186) );
in01f80 g562258 ( .a(n_10228), .o(n_6236) );
no02f80 g562259 ( .a(n_5574), .b(n_5331), .o(n_10228) );
na02f80 g562260 ( .a(n_7204), .b(n_5164), .o(n_9396) );
no02f80 g562261 ( .a(n_6234), .b(n_6478), .o(n_6235) );
no02f80 g562262 ( .a(n_5682), .b(x_in_19_12), .o(n_5495) );
in01f80 g562263 ( .a(n_6233), .o(n_11258) );
no02f80 g562264 ( .a(n_5682), .b(n_5244), .o(n_6233) );
in01f80 g562265 ( .a(n_6971), .o(n_8505) );
no02f80 g562266 ( .a(n_5683), .b(x_in_27_11), .o(n_6971) );
na02f80 g562267 ( .a(n_6231), .b(n_6230), .o(n_6232) );
in01f80 g562268 ( .a(n_6229), .o(n_10247) );
no02f80 g562269 ( .a(n_5494), .b(n_8443), .o(n_6229) );
in01f80 g562270 ( .a(n_6228), .o(n_10250) );
no02f80 g562271 ( .a(n_5493), .b(n_8513), .o(n_6228) );
in01f80 g562272 ( .a(n_6465), .o(n_8446) );
no02f80 g562273 ( .a(n_5492), .b(x_in_43_11), .o(n_6465) );
no02f80 g562274 ( .a(n_5490), .b(n_5489), .o(n_5491) );
in01f80 g562275 ( .a(n_6649), .o(n_10231) );
no02f80 g562276 ( .a(n_6429), .b(n_5332), .o(n_6649) );
in01f80 g562277 ( .a(n_8520), .o(n_7724) );
no02f80 g562278 ( .a(n_5684), .b(x_in_51_11), .o(n_8520) );
in01f80 g562279 ( .a(n_6227), .o(n_10244) );
no02f80 g562280 ( .a(n_5096), .b(n_6746), .o(n_6227) );
in01f80 g562281 ( .a(n_7414), .o(n_7415) );
na02f80 g562282 ( .a(n_5179), .b(x_in_17_4), .o(n_7414) );
na02f80 g562283 ( .a(n_4879), .b(x_in_3_11), .o(n_11682) );
na02f80 g562284 ( .a(n_6225), .b(n_5988), .o(n_6226) );
in01f80 g562285 ( .a(n_6964), .o(n_8507) );
no02f80 g562286 ( .a(n_5041), .b(x_in_3_11), .o(n_6964) );
na02f80 g562287 ( .a(n_6223), .b(n_7445), .o(n_6224) );
in01f80 g562288 ( .a(n_6948), .o(n_8487) );
no02f80 g562289 ( .a(n_5488), .b(x_in_19_11), .o(n_6948) );
in01f80 g562290 ( .a(n_6222), .o(n_11235) );
no02f80 g562291 ( .a(n_5487), .b(n_7765), .o(n_6222) );
no02f80 g562292 ( .a(n_5433), .b(n_5485), .o(n_5486) );
na02f80 g562293 ( .a(n_5238), .b(x_in_17_13), .o(n_7207) );
no02f80 g562294 ( .a(n_6648), .b(n_5128), .o(n_17495) );
na02f80 g562295 ( .a(n_5483), .b(n_5482), .o(n_5484) );
no02f80 g562296 ( .a(n_6220), .b(n_6219), .o(n_6221) );
na02f80 g562297 ( .a(n_6217), .b(n_6216), .o(n_6218) );
no02f80 g562298 ( .a(n_6476), .b(n_6475), .o(n_5481) );
na02f80 g562299 ( .a(n_6647), .b(n_4962), .o(n_8395) );
na02f80 g562300 ( .a(n_6646), .b(n_5793), .o(n_16639) );
no02f80 g562301 ( .a(n_4971), .b(n_4032), .o(n_9096) );
no02f80 g562302 ( .a(n_5479), .b(n_5478), .o(n_5480) );
na02f80 g562303 ( .a(n_6626), .b(FE_OFN692_n_6708), .o(n_5477) );
na02f80 g562304 ( .a(n_6476), .b(n_5476), .o(n_13226) );
na02f80 g562305 ( .a(n_6476), .b(n_5889), .o(n_5475) );
na02f80 g562306 ( .a(n_6629), .b(n_6715), .o(n_5474) );
na02f80 g562307 ( .a(n_6005), .b(n_6709), .o(n_5473) );
ao12f80 g562308 ( .a(n_4818), .b(n_4364), .c(n_3087), .o(n_9881) );
na02f80 g562309 ( .a(n_6214), .b(n_6213), .o(n_6215) );
no02f80 g562310 ( .a(n_4404), .b(n_7581), .o(n_6212) );
na02f80 g562311 ( .a(n_6210), .b(n_6209), .o(n_6211) );
na02f80 g562312 ( .a(n_5471), .b(n_6713), .o(n_5472) );
no02f80 g562313 ( .a(n_6207), .b(n_6437), .o(n_6208) );
na02f80 g562314 ( .a(n_5469), .b(n_5468), .o(n_5470) );
no02f80 g562315 ( .a(n_6007), .b(n_6749), .o(n_5467) );
na02f80 g562316 ( .a(n_5465), .b(n_5464), .o(n_5466) );
no02f80 g562317 ( .a(n_5784), .b(n_9088), .o(n_5463) );
na02f80 g562318 ( .a(n_6205), .b(n_6204), .o(n_6206) );
na02f80 g562319 ( .a(n_4612), .b(n_6203), .o(n_7954) );
na02f80 g562320 ( .a(n_6201), .b(n_6200), .o(n_6202) );
na02f80 g562321 ( .a(n_5461), .b(n_5460), .o(n_5462) );
oa12f80 g562322 ( .a(n_5992), .b(n_5993), .c(n_3089), .o(n_11508) );
ao12f80 g562323 ( .a(n_5990), .b(n_5991), .c(n_3086), .o(n_10787) );
oa12f80 g562324 ( .a(n_5459), .b(n_4817), .c(n_3280), .o(n_9345) );
ao22s80 g562325 ( .a(n_5380), .b(n_3219), .c(n_7156), .d(n_5430), .o(n_10177) );
na02f80 g562326 ( .a(n_6198), .b(FE_OFN1262_n_6197), .o(n_6199) );
ao12f80 g562327 ( .a(n_5994), .b(n_5995), .c(n_3088), .o(n_9343) );
oa12f80 g562328 ( .a(n_10073), .b(n_6296), .c(x_in_13_3), .o(n_7988) );
no02f80 g562329 ( .a(n_5457), .b(n_5456), .o(n_5458) );
oa12f80 g562330 ( .a(n_9385), .b(n_4787), .c(x_in_31_4), .o(n_7979) );
na02f80 g562331 ( .a(n_7019), .b(n_7385), .o(n_6196) );
na02f80 g562332 ( .a(n_6194), .b(n_6193), .o(n_6195) );
no02f80 g562333 ( .a(n_6191), .b(n_6190), .o(n_6192) );
oa12f80 g562334 ( .a(n_10103), .b(n_4788), .c(x_in_55_4), .o(n_7981) );
oa12f80 g562335 ( .a(n_10105), .b(n_4785), .c(x_in_15_4), .o(n_7992) );
ao12f80 g562336 ( .a(n_8408), .b(n_5212), .c(n_5211), .o(n_8407) );
na02f80 g562337 ( .a(n_6188), .b(n_6187), .o(n_6189) );
oa12f80 g562338 ( .a(n_4365), .b(n_3889), .c(n_3085), .o(n_11495) );
na02f80 g562339 ( .a(n_6185), .b(n_6184), .o(n_6186) );
na02f80 g562340 ( .a(n_6182), .b(n_6181), .o(n_6183) );
na02f80 g562341 ( .a(n_6179), .b(FE_OFN1260_n_6178), .o(n_6180) );
na02f80 g562342 ( .a(n_6176), .b(n_6175), .o(n_6177) );
ao22s80 g562343 ( .a(n_5335), .b(n_3167), .c(n_6504), .d(n_5336), .o(n_10175) );
na02f80 g562344 ( .a(n_6173), .b(n_6172), .o(n_6174) );
ao12f80 g562345 ( .a(n_14491), .b(n_4765), .c(n_4828), .o(n_9180) );
na02f80 g562346 ( .a(n_6170), .b(n_6169), .o(n_6171) );
oa12f80 g562347 ( .a(n_10107), .b(n_4790), .c(x_in_23_4), .o(n_7996) );
oa12f80 g562348 ( .a(n_6070), .b(n_858), .c(n_25680), .o(n_7413) );
na02f80 g562349 ( .a(n_6167), .b(FE_OFN578_n_6424), .o(n_6168) );
na02f80 g562350 ( .a(n_6165), .b(n_6164), .o(n_6166) );
na02f80 g562351 ( .a(n_6162), .b(n_6161), .o(n_6163) );
in01f80 g562352 ( .a(n_6644), .o(n_6645) );
ao12f80 g562353 ( .a(n_3362), .b(n_3236), .c(n_5923), .o(n_6644) );
ao12f80 g562354 ( .a(n_8416), .b(n_6563), .c(n_5023), .o(n_8413) );
na02f80 g562355 ( .a(n_6027), .b(n_6026), .o(n_6028) );
na02f80 g562356 ( .a(n_6439), .b(n_6438), .o(n_6440) );
oa12f80 g562357 ( .a(n_10101), .b(n_4789), .c(x_in_47_4), .o(n_7990) );
na02f80 g562358 ( .a(n_6158), .b(FE_OFN875_n_6157), .o(n_6159) );
na02f80 g562359 ( .a(n_6155), .b(FE_OFN871_n_6154), .o(n_6156) );
na02f80 g562360 ( .a(n_6152), .b(FE_OFN867_n_6151), .o(n_6153) );
no02f80 g562361 ( .a(n_6149), .b(n_6148), .o(n_6150) );
na02f80 g562362 ( .a(n_6146), .b(n_6145), .o(n_6147) );
ao22s80 g562363 ( .a(n_5364), .b(n_3168), .c(n_7159), .d(n_5365), .o(n_11082) );
na02f80 g562364 ( .a(n_6143), .b(n_6142), .o(n_6144) );
no02f80 g562365 ( .a(n_5454), .b(n_5453), .o(n_5455) );
na02f80 g562366 ( .a(n_5764), .b(n_5763), .o(n_5765) );
no02f80 g562367 ( .a(n_6140), .b(n_6139), .o(n_6141) );
no02f80 g562368 ( .a(n_6137), .b(n_6136), .o(n_6138) );
na02f80 g562369 ( .a(n_6134), .b(n_6133), .o(n_6135) );
na02f80 g562370 ( .a(n_6445), .b(FE_OFN706_n_6444), .o(n_6446) );
na02f80 g562371 ( .a(n_5725), .b(n_6017), .o(n_5726) );
no02f80 g562372 ( .a(n_6131), .b(n_6373), .o(n_6132) );
na02f80 g562373 ( .a(n_6129), .b(n_6128), .o(n_6130) );
no02f80 g562374 ( .a(n_6126), .b(n_6125), .o(n_6127) );
ao22s80 g562375 ( .a(n_5372), .b(n_3166), .c(n_7153), .d(n_5373), .o(n_12127) );
na02f80 g562376 ( .a(n_6123), .b(n_6122), .o(n_6124) );
oa12f80 g562377 ( .a(n_10097), .b(n_4786), .c(x_in_63_4), .o(n_7986) );
na02f80 g562378 ( .a(n_6120), .b(n_6119), .o(n_6121) );
na02f80 g562379 ( .a(n_6117), .b(FE_OFN1278_n_6116), .o(n_6118) );
na02f80 g562380 ( .a(n_6114), .b(n_6113), .o(n_6115) );
na02f80 g562381 ( .a(n_6111), .b(n_6110), .o(n_6112) );
no02f80 g562382 ( .a(n_6108), .b(n_6107), .o(n_6109) );
na02f80 g562383 ( .a(n_6105), .b(n_6104), .o(n_6106) );
na02f80 g562384 ( .a(n_6102), .b(n_6101), .o(n_6103) );
na02f80 g562385 ( .a(n_6099), .b(n_6098), .o(n_6100) );
no02f80 g562386 ( .a(n_5451), .b(n_5450), .o(n_5452) );
oa12f80 g562387 ( .a(n_7221), .b(n_223), .c(FE_OFN76_n_27012), .o(n_7412) );
no02f80 g562388 ( .a(n_7218), .b(n_6081), .o(n_7219) );
na02f80 g562389 ( .a(n_6096), .b(n_6095), .o(n_6097) );
ao12f80 g562390 ( .a(n_4861), .b(n_3646), .c(x_in_13_3), .o(n_8842) );
ao22s80 g562391 ( .a(n_5350), .b(n_3163), .c(n_7150), .d(n_5351), .o(n_10169) );
na02f80 g562392 ( .a(n_4353), .b(n_5729), .o(n_14582) );
no02f80 g562393 ( .a(n_6092), .b(n_6315), .o(n_6093) );
ao22s80 g562394 ( .a(n_4945), .b(n_3161), .c(n_7162), .d(n_4946), .o(n_10171) );
oa12f80 g562395 ( .a(n_10059), .b(n_4891), .c(x_in_45_4), .o(n_7994) );
in01f80 g562396 ( .a(n_11579), .o(n_7983) );
ao12f80 g562397 ( .a(n_7958), .b(n_4020), .c(n_7195), .o(n_11579) );
ao12f80 g562398 ( .a(n_8412), .b(n_5218), .c(n_5217), .o(n_8411) );
ao12f80 g562399 ( .a(n_8410), .b(n_6571), .c(n_5219), .o(n_8409) );
ao12f80 g562400 ( .a(n_8406), .b(n_6577), .c(n_5221), .o(n_8401) );
no02f80 g562401 ( .a(n_5448), .b(n_5447), .o(n_5449) );
oa12f80 g562402 ( .a(n_7964), .b(n_5864), .c(x_in_9_1), .o(n_5710) );
na02f80 g562403 ( .a(n_6090), .b(FE_OFN1222_n_6089), .o(n_6091) );
oa12f80 g562404 ( .a(n_9422), .b(n_4895), .c(n_4894), .o(n_7866) );
oa12f80 g562405 ( .a(n_4833), .b(n_4832), .c(x_in_41_0), .o(n_4834) );
na02f80 g562406 ( .a(n_6087), .b(n_6086), .o(n_6088) );
ao12f80 g562407 ( .a(n_5191), .b(n_5250), .c(n_5446), .o(n_8394) );
na02f80 g562408 ( .a(n_6084), .b(n_6083), .o(n_6085) );
no02f80 g562409 ( .a(n_6082), .b(n_6081), .o(n_7620) );
na02f80 g562410 ( .a(n_6079), .b(n_6078), .o(n_6080) );
no02f80 g562411 ( .a(n_6076), .b(n_6075), .o(n_6077) );
na02f80 g562412 ( .a(n_6073), .b(FE_OFN550_n_6072), .o(n_6074) );
na02f80 g562413 ( .a(n_5714), .b(n_5713), .o(n_5715) );
oa12f80 g562414 ( .a(n_6070), .b(n_868), .c(FE_OFN1106_rst), .o(n_6071) );
na02f80 g562415 ( .a(n_5718), .b(n_5913), .o(n_5719) );
na02f80 g562416 ( .a(n_5721), .b(FE_OFN991_n_5720), .o(n_5722) );
na02f80 g562417 ( .a(n_6068), .b(n_6067), .o(n_6069) );
no02f80 g562418 ( .a(n_6065), .b(n_6064), .o(n_6066) );
na02f80 g562419 ( .a(n_6062), .b(n_6061), .o(n_6063) );
oa12f80 g562420 ( .a(n_7221), .b(n_1535), .c(FE_OFN127_n_27449), .o(n_7222) );
oa12f80 g562421 ( .a(n_7973), .b(n_8477), .c(n_5723), .o(n_5724) );
no02f80 g562422 ( .a(n_6059), .b(n_6058), .o(n_6060) );
na02f80 g562423 ( .a(n_6056), .b(n_6055), .o(n_6057) );
na02f80 g562424 ( .a(n_6053), .b(n_6052), .o(n_6054) );
na02f80 g562425 ( .a(n_6050), .b(n_6049), .o(n_6051) );
no02f80 g562426 ( .a(n_4906), .b(FE_OFN1258_n_4905), .o(n_4907) );
oa12f80 g562427 ( .a(n_4830), .b(n_289), .c(x_in_25_3), .o(n_4831) );
na03f80 g562428 ( .a(n_4592), .b(n_4828), .c(x_in_29_0), .o(n_4829) );
oa12f80 g562429 ( .a(n_7961), .b(n_5844), .c(n_5443), .o(n_5444) );
oa12f80 g562430 ( .a(n_6047), .b(n_5840), .c(n_3447), .o(n_6048) );
oa22f80 g562431 ( .a(n_3635), .b(n_4280), .c(n_1513), .d(FE_OFN105_n_27449), .o(n_7411) );
oa12f80 g562432 ( .a(n_7225), .b(n_1022), .c(FE_OFN1181_rst), .o(n_6046) );
oa12f80 g562433 ( .a(n_7409), .b(n_669), .c(FE_OFN60_n_27012), .o(n_7410) );
oa12f80 g562434 ( .a(n_7409), .b(n_1293), .c(FE_OFN193_n_28928), .o(n_7408) );
oa22f80 g562435 ( .a(n_3633), .b(n_29046), .c(n_546), .d(n_27449), .o(n_7224) );
oa12f80 g562436 ( .a(n_7225), .b(n_180), .c(FE_OFN134_n_27449), .o(n_7226) );
oa12f80 g562437 ( .a(n_4826), .b(n_4825), .c(x_in_53_3), .o(n_4827) );
ao12f80 g562438 ( .a(n_7129), .b(n_6576), .c(n_5207), .o(n_8415) );
ao12f80 g562439 ( .a(n_5593), .b(n_8618), .c(n_4732), .o(n_5442) );
oa12f80 g562440 ( .a(n_5440), .b(n_8114), .c(x_in_33_12), .o(n_5441) );
ao12f80 g562441 ( .a(n_5589), .b(n_12606), .c(n_2629), .o(n_5439) );
oa12f80 g562442 ( .a(n_10920), .b(n_2935), .c(x_in_49_2), .o(n_5438) );
oa12f80 g562443 ( .a(x_in_49_1), .b(n_3510), .c(x_in_49_0), .o(n_4824) );
oa12f80 g562444 ( .a(n_4175), .b(n_5308), .c(x_in_57_10), .o(n_13288) );
oa12f80 g562445 ( .a(n_6044), .b(n_5847), .c(x_in_7_4), .o(n_6045) );
oa12f80 g562446 ( .a(n_6042), .b(n_5828), .c(x_in_61_4), .o(n_6043) );
oa12f80 g562447 ( .a(n_7166), .b(n_5328), .c(x_in_13_1), .o(n_10099) );
oa22f80 g562448 ( .a(n_3066), .b(x_in_33_1), .c(n_5319), .d(x_in_33_0), .o(n_7945) );
na03f80 g562449 ( .a(n_5277), .b(n_3605), .c(x_in_25_1), .o(n_6040) );
in01f80 g562450 ( .a(n_9602), .o(n_8440) );
oa12f80 g562451 ( .a(n_5426), .b(n_5425), .c(x_in_21_15), .o(n_9602) );
oa22f80 g562452 ( .a(n_3275), .b(n_6216), .c(n_4346), .d(n_4345), .o(n_12344) );
in01f80 g562454 ( .a(n_10151), .o(n_6037) );
oa12f80 g562455 ( .a(n_5446), .b(n_5436), .c(n_5435), .o(n_10151) );
ao22s80 g562456 ( .a(n_4820), .b(n_2150), .c(x_in_33_1), .d(x_in_33_0), .o(n_9831) );
oa12f80 g562457 ( .a(n_4685), .b(n_3566), .c(n_5848), .o(n_7196) );
ao22s80 g562458 ( .a(n_4061), .b(n_6213), .c(n_4483), .d(n_4482), .o(n_11832) );
ao12f80 g562459 ( .a(n_5091), .b(n_4702), .c(n_6653), .o(n_6036) );
no02f80 g562460 ( .a(n_6282), .b(n_4723), .o(n_6035) );
oa22f80 g562461 ( .a(n_3112), .b(x_in_57_1), .c(n_5267), .d(x_in_57_0), .o(n_8025) );
ao12f80 g562462 ( .a(n_8414), .b(n_5210), .c(n_5209), .o(n_8417) );
ao12f80 g562463 ( .a(n_4581), .b(n_4432), .c(n_4433), .o(n_11844) );
ao12f80 g562464 ( .a(n_4584), .b(n_4436), .c(n_4437), .o(n_11838) );
ao12f80 g562465 ( .a(n_3262), .b(FE_OFN1250_n_5334), .c(x_in_51_13), .o(n_9440) );
ao22s80 g562466 ( .a(n_2846), .b(n_6139), .c(n_4455), .d(n_4453), .o(n_12367) );
ao12f80 g562467 ( .a(n_4810), .b(n_4446), .c(n_4447), .o(n_11850) );
oa22f80 g562468 ( .a(n_3080), .b(FE_OFN550_n_6072), .c(n_3878), .d(n_4479), .o(n_11900) );
ao12f80 g562469 ( .a(n_4973), .b(n_5189), .c(n_6641), .o(n_6642) );
ao12f80 g562470 ( .a(n_4576), .b(n_4421), .c(n_4422), .o(n_7617) );
ao22s80 g562471 ( .a(n_3693), .b(n_6373), .c(n_6372), .d(n_4480), .o(n_11915) );
ao22s80 g562472 ( .a(n_3512), .b(n_6058), .c(n_5265), .d(n_4475), .o(n_11896) );
in01f80 g562473 ( .a(n_6033), .o(n_6034) );
oa22f80 g562474 ( .a(n_2862), .b(n_5057), .c(n_7088), .d(x_in_25_6), .o(n_6033) );
in01f80 g562475 ( .a(n_6640), .o(n_11903) );
oa12f80 g562476 ( .a(n_4171), .b(n_6032), .c(n_4166), .o(n_6640) );
oa22f80 g562477 ( .a(n_3142), .b(n_6061), .c(n_4504), .d(n_4503), .o(n_12368) );
ao12f80 g562478 ( .a(n_4572), .b(n_4797), .c(n_4798), .o(n_11863) );
oa22f80 g562479 ( .a(n_3283), .b(n_6145), .c(n_4488), .d(n_4487), .o(n_11949) );
oa22f80 g562480 ( .a(n_3137), .b(n_6128), .c(n_4442), .d(n_4441), .o(n_11912) );
oa22f80 g562481 ( .a(n_3286), .b(n_6101), .c(n_4465), .d(n_4464), .o(n_11879) );
oa22f80 g562482 ( .a(n_2840), .b(n_6142), .c(n_4507), .d(n_4506), .o(n_12318) );
no02f80 g562483 ( .a(n_6276), .b(n_3540), .o(n_6031) );
ao12f80 g562484 ( .a(n_3071), .b(n_3751), .c(x_in_41_14), .o(n_7914) );
oa22f80 g562485 ( .a(n_3133), .b(n_5315), .c(n_7082), .d(x_in_25_7), .o(n_9825) );
ao12f80 g562486 ( .a(n_5381), .b(n_4823), .c(n_4822), .o(n_11333) );
ao22s80 g562487 ( .a(n_2706), .b(n_6136), .c(n_5263), .d(n_4456), .o(n_11930) );
oa12f80 g562488 ( .a(n_5433), .b(n_2956), .c(n_8756), .o(n_5434) );
oa12f80 g562489 ( .a(n_6030), .b(n_5930), .c(x_in_3_2), .o(n_9684) );
ao12f80 g562490 ( .a(n_9982), .b(n_3542), .c(x_in_5_3), .o(n_7175) );
oa12f80 g562491 ( .a(n_2878), .b(n_5123), .c(x_in_59_4), .o(n_7933) );
ao12f80 g562492 ( .a(n_4870), .b(n_5299), .c(n_6781), .o(n_5300) );
oa22f80 g562493 ( .a(n_3688), .b(n_6122), .c(n_4474), .d(n_4473), .o(n_11893) );
in01f80 g562494 ( .a(n_10684), .o(n_6422) );
oa22f80 g562495 ( .a(n_2722), .b(n_5318), .c(n_7079), .d(x_in_25_12), .o(n_10684) );
in01f80 g562496 ( .a(n_9813), .o(n_6029) );
oa22f80 g562497 ( .a(n_3130), .b(n_5316), .c(n_7073), .d(x_in_25_8), .o(n_9813) );
ao12f80 g562498 ( .a(n_2295), .b(n_4821), .c(n_2568), .o(n_9827) );
in01f80 g562499 ( .a(n_10689), .o(n_6423) );
oa22f80 g562500 ( .a(n_2744), .b(n_4909), .c(n_7067), .d(x_in_25_10), .o(n_10689) );
in01f80 g562501 ( .a(FE_OFN1276_n_12754), .o(n_6025) );
oa22f80 g562502 ( .a(n_2761), .b(FE_OFN1278_n_6116), .c(n_4472), .d(n_4471), .o(n_12754) );
in01f80 g562503 ( .a(FE_OFN572_n_12800), .o(n_7203) );
oa22f80 g562504 ( .a(n_4131), .b(FE_OFN578_n_6424), .c(n_4370), .d(n_4369), .o(n_12800) );
in01f80 g562505 ( .a(n_12787), .o(n_6024) );
oa22f80 g562506 ( .a(n_3296), .b(FE_OFN875_n_6157), .c(n_4532), .d(n_4531), .o(n_12787) );
oa22f80 g562507 ( .a(n_2778), .b(n_5285), .c(n_7064), .d(x_in_25_11), .o(n_9829) );
ao12f80 g562508 ( .a(n_3854), .b(n_4928), .c(n_4890), .o(n_11870) );
ao12f80 g562509 ( .a(n_4568), .b(n_4582), .c(n_4583), .o(n_11946) );
ao12f80 g562510 ( .a(n_4565), .b(n_4258), .c(n_4259), .o(n_11909) );
oa22f80 g562511 ( .a(n_2816), .b(n_6133), .c(n_4885), .d(n_4883), .o(n_12373) );
ao12f80 g562512 ( .a(n_4564), .b(n_6023), .c(n_4427), .o(n_11985) );
oa22f80 g562513 ( .a(n_2694), .b(n_6095), .c(n_4499), .d(n_4497), .o(n_11964) );
ao12f80 g562514 ( .a(n_4563), .b(n_6022), .c(n_4512), .o(n_12012) );
oa22f80 g562515 ( .a(n_3123), .b(n_6119), .c(n_4524), .d(n_4522), .o(n_12369) );
oa12f80 g562516 ( .a(n_7020), .b(n_3911), .c(x_in_57_4), .o(n_7165) );
ao22s80 g562517 ( .a(n_3671), .b(n_6064), .c(n_6021), .d(n_4145), .o(n_12033) );
oa12f80 g562518 ( .a(n_4476), .b(n_3646), .c(n_2224), .o(n_7113) );
ao12f80 g562519 ( .a(n_4560), .b(n_4461), .c(n_4462), .o(n_11876) );
ao12f80 g562520 ( .a(n_4559), .b(n_4450), .c(n_4451), .o(n_11994) );
ao22s80 g562521 ( .a(n_4095), .b(n_6190), .c(n_4521), .d(n_4520), .o(n_12042) );
oa22f80 g562522 ( .a(n_3288), .b(n_6438), .c(n_2444), .d(n_4457), .o(n_11968) );
oa22f80 g562523 ( .a(n_3374), .b(n_6078), .c(n_4444), .d(n_4443), .o(n_12030) );
oa22f80 g562524 ( .a(n_4136), .b(FE_OFN871_n_6154), .c(n_4496), .d(n_4495), .o(n_11961) );
oa22f80 g562525 ( .a(n_3469), .b(FE_OFN706_n_6444), .c(n_4459), .d(n_4458), .o(n_11927) );
oa22f80 g562526 ( .a(n_3452), .b(n_6104), .c(n_4199), .d(n_4198), .o(n_12372) );
oa22f80 g562527 ( .a(n_3667), .b(FE_OFN1262_n_6197), .c(n_4430), .d(n_4429), .o(n_12007) );
ao12f80 g562528 ( .a(n_4558), .b(n_4373), .c(n_4374), .o(n_11982) );
ao12f80 g562529 ( .a(n_4557), .b(n_4515), .c(n_4516), .o(n_11976) );
oa22f80 g562530 ( .a(n_3340), .b(n_6110), .c(n_4467), .d(n_4466), .o(n_12370) );
oa22f80 g562531 ( .a(n_3121), .b(n_6187), .c(n_4414), .d(n_4413), .o(n_12022) );
oa22f80 g562532 ( .a(n_3329), .b(FE_OFN1260_n_6178), .c(n_4501), .d(n_4500), .o(n_12351) );
oa22f80 g562533 ( .a(n_4092), .b(n_6204), .c(n_4186), .d(n_4185), .o(n_11866) );
oa12f80 g562534 ( .a(n_6512), .b(n_6521), .c(x_in_35_3), .o(n_8838) );
in01f80 g562535 ( .a(n_12811), .o(n_6020) );
oa22f80 g562536 ( .a(n_3302), .b(n_6169), .c(n_4310), .d(n_4309), .o(n_12811) );
in01f80 g562537 ( .a(FE_OFN987_n_12804), .o(n_6019) );
oa22f80 g562538 ( .a(n_3308), .b(n_6181), .c(n_4509), .d(n_4508), .o(n_12804) );
in01f80 g562539 ( .a(FE_OFN1216_n_12761), .o(n_6018) );
oa22f80 g562540 ( .a(n_3116), .b(FE_OFN1222_n_6089), .c(n_4485), .d(n_4484), .o(n_12761) );
oa12f80 g562541 ( .a(n_5432), .b(n_3604), .c(x_in_33_5), .o(n_8185) );
oa22f80 g562542 ( .a(n_3674), .b(n_6052), .c(n_4412), .d(n_4411), .o(n_11955) );
oa22f80 g562543 ( .a(n_3422), .b(n_6017), .c(n_4440), .d(n_4439), .o(n_11921) );
ao12f80 g562544 ( .a(n_4556), .b(n_4492), .c(n_4493), .o(n_11973) );
oa22f80 g562545 ( .a(n_3118), .b(n_6067), .c(n_2425), .d(n_4408), .o(n_12001) );
oa22f80 g562546 ( .a(n_3297), .b(n_6026), .c(n_2524), .d(n_4486), .o(n_11814) );
ao22s80 g562547 ( .a(n_3433), .b(n_6107), .c(n_4218), .d(n_4217), .o(n_11882) );
ao22s80 g562548 ( .a(n_4045), .b(x_in_19_13), .c(x_in_19_14), .d(x_in_19_12), .o(n_6016) );
ao22s80 g562549 ( .a(n_3461), .b(n_6148), .c(n_4490), .d(n_4489), .o(n_11952) );
ao22s80 g562550 ( .a(n_3664), .b(n_6315), .c(n_4210), .d(n_4209), .o(n_11918) );
na02f80 g562551 ( .a(n_5138), .b(n_8360), .o(n_6639) );
oa22f80 g562552 ( .a(n_2867), .b(FE_OFN867_n_6151), .c(n_4549), .d(n_4547), .o(n_11958) );
ao22s80 g562553 ( .a(n_4112), .b(n_6075), .c(n_6015), .d(n_4425), .o(n_11924) );
oa12f80 g562554 ( .a(n_6014), .b(n_5732), .c(x_in_3_6), .o(n_9584) );
ao12f80 g562555 ( .a(n_4809), .b(n_4807), .c(x_in_1_1), .o(n_7206) );
ao12f80 g562556 ( .a(n_4241), .b(n_6013), .c(n_4502), .o(n_11979) );
oa22f80 g562557 ( .a(n_3111), .b(n_6161), .c(n_4390), .d(n_4388), .o(n_12025) );
oa22f80 g562558 ( .a(n_2882), .b(n_6113), .c(n_4470), .d(n_4468), .o(n_12371) );
oa22f80 g562559 ( .a(n_2887), .b(n_6083), .c(n_4225), .d(n_4223), .o(n_12004) );
ao12f80 g562560 ( .a(n_6011), .b(n_3631), .c(n_2555), .o(n_6012) );
ao12f80 g562561 ( .a(x_in_61_3), .b(n_4197), .c(n_5431), .o(n_10902) );
in01f80 g562562 ( .a(n_6637), .o(n_6638) );
ao12f80 g562563 ( .a(n_8358), .b(n_6216), .c(n_4659), .o(n_6637) );
ao22s80 g562564 ( .a(n_3569), .b(n_5294), .c(n_6952), .d(x_in_5_6), .o(n_9807) );
oa12f80 g562565 ( .a(n_6010), .b(n_5874), .c(x_in_3_4), .o(n_9581) );
ao22s80 g562566 ( .a(n_5456), .b(n_2687), .c(n_3749), .d(x_in_15_2), .o(n_12016) );
ao22s80 g562567 ( .a(n_5447), .b(n_2572), .c(n_3764), .d(x_in_63_2), .o(n_11873) );
oa12f80 g562568 ( .a(n_3823), .b(n_3761), .c(n_5430), .o(n_12019) );
ao22s80 g562569 ( .a(FE_OFN1258_n_4905), .b(n_2566), .c(n_4065), .d(x_in_55_2), .o(n_11991) );
na02f80 g562570 ( .a(n_5428), .b(n_3884), .o(n_5429) );
oa12f80 g562571 ( .a(n_9932), .b(n_5322), .c(n_3387), .o(n_7171) );
ao12f80 g562572 ( .a(n_3819), .b(n_2147), .c(x_in_47_2), .o(n_11943) );
ao12f80 g562573 ( .a(n_3492), .b(n_2205), .c(x_in_31_2), .o(n_11906) );
oa12f80 g562574 ( .a(n_5427), .b(n_3896), .c(x_in_33_4), .o(n_8750) );
oa12f80 g562575 ( .a(x_in_17_2), .b(n_5853), .c(n_3723), .o(n_11339) );
oa12f80 g562576 ( .a(n_5426), .b(n_5425), .c(n_5872), .o(n_7772) );
oa12f80 g562577 ( .a(n_6636), .b(n_4969), .c(x_in_33_9), .o(n_8966) );
oa12f80 g562578 ( .a(n_5424), .b(n_3359), .c(x_in_33_6), .o(n_8173) );
oa12f80 g562579 ( .a(n_5423), .b(n_3636), .c(x_in_33_10), .o(n_8182) );
oa12f80 g562580 ( .a(n_5064), .b(n_3891), .c(x_in_33_8), .o(n_8179) );
oa12f80 g562581 ( .a(n_5422), .b(n_3403), .c(x_in_33_7), .o(n_8176) );
oa12f80 g562582 ( .a(n_5421), .b(FE_OFN933_n_4950), .c(x_in_51_9), .o(n_7176) );
ao22s80 g562583 ( .a(n_4819), .b(n_2640), .c(n_2769), .d(x_in_25_11), .o(n_6415) );
oa12f80 g562584 ( .a(n_5759), .b(n_12697), .c(x_in_33_11), .o(n_8742) );
ao12f80 g562585 ( .a(n_5471), .b(n_8737), .c(n_2994), .o(n_5420) );
ao12f80 g562586 ( .a(n_3770), .b(n_5489), .c(n_5418), .o(n_5419) );
ao12f80 g562587 ( .a(n_6223), .b(FE_OFN1087_n_8974), .c(n_3576), .o(n_6009) );
oa12f80 g562588 ( .a(n_3244), .b(n_2854), .c(n_5306), .o(n_9819) );
in01f80 g562589 ( .a(n_6634), .o(n_6635) );
ao22s80 g562590 ( .a(n_3561), .b(n_5276), .c(n_6912), .d(x_in_57_13), .o(n_6634) );
in01f80 g562591 ( .a(n_6632), .o(n_6633) );
ao22s80 g562592 ( .a(n_3416), .b(n_5288), .c(n_6923), .d(x_in_5_13), .o(n_6632) );
ao12f80 g562593 ( .a(n_6007), .b(n_8725), .c(n_2995), .o(n_6008) );
in01f80 g562594 ( .a(n_6631), .o(n_8905) );
ao22s80 g562595 ( .a(n_4100), .b(n_7498), .c(n_4957), .d(n_4231), .o(n_6631) );
oa12f80 g562596 ( .a(n_2710), .b(n_2852), .c(n_5036), .o(n_9860) );
na02f80 g562597 ( .a(n_6005), .b(n_4682), .o(n_6006) );
na02f80 g562598 ( .a(n_6629), .b(n_5169), .o(n_6630) );
in01f80 g562599 ( .a(FE_OFN1232_n_12068), .o(n_6004) );
ao22s80 g562600 ( .a(n_5645), .b(n_2569), .c(n_4955), .d(x_in_41_10), .o(n_12068) );
ao22s80 g562601 ( .a(n_5417), .b(n_2631), .c(n_5416), .d(x_in_49_1), .o(n_12940) );
oa12f80 g562602 ( .a(n_6628), .b(n_6958), .c(x_in_51_11), .o(n_8392) );
na02f80 g562603 ( .a(n_6626), .b(n_5043), .o(n_6627) );
ao12f80 g562604 ( .a(n_4542), .b(n_7693), .c(x_in_21_13), .o(n_10646) );
no02f80 g562605 ( .a(n_6849), .b(n_3915), .o(n_4966) );
ao12f80 g562606 ( .a(n_6929), .b(n_4868), .c(x_in_17_5), .o(n_9980) );
in01f80 g562607 ( .a(n_6624), .o(n_6625) );
ao22s80 g562608 ( .a(n_4036), .b(n_5389), .c(n_6895), .d(x_in_5_10), .o(n_6624) );
in01f80 g562609 ( .a(n_11134), .o(n_6623) );
oa12f80 g562610 ( .a(n_4366), .b(n_3868), .c(n_5381), .o(n_11134) );
ao12f80 g562611 ( .a(n_5178), .b(n_5853), .c(n_4687), .o(n_8581) );
oa12f80 g562612 ( .a(n_4539), .b(n_7710), .c(n_5977), .o(n_10640) );
ao12f80 g562613 ( .a(n_4552), .b(n_5902), .c(x_in_33_4), .o(n_10687) );
in01f80 g562614 ( .a(n_8488), .o(n_5739) );
oa12f80 g562615 ( .a(n_3754), .b(n_2086), .c(n_5415), .o(n_8488) );
oa12f80 g562616 ( .a(n_2702), .b(n_3264), .c(n_5305), .o(n_9850) );
ao22s80 g562617 ( .a(n_4056), .b(n_5361), .c(n_6889), .d(x_in_57_7), .o(n_9817) );
oa22f80 g562618 ( .a(n_3335), .b(n_5903), .c(n_2462), .d(n_5869), .o(n_10633) );
in01f80 g562619 ( .a(n_6621), .o(n_6622) );
ao22s80 g562620 ( .a(n_3391), .b(n_5289), .c(n_6802), .d(x_in_5_12), .o(n_6621) );
na02f80 g562621 ( .a(n_5540), .b(n_3835), .o(n_5414) );
in01f80 g562622 ( .a(n_6002), .o(n_6003) );
ao22s80 g562623 ( .a(n_2807), .b(n_5885), .c(n_7658), .d(x_in_37_12), .o(n_6002) );
in01f80 g562624 ( .a(n_6619), .o(n_6620) );
ao22s80 g562625 ( .a(n_4064), .b(n_5303), .c(n_6881), .d(x_in_57_12), .o(n_6619) );
ao22s80 g562626 ( .a(n_5642), .b(n_2314), .c(n_5395), .d(x_in_41_8), .o(n_11302) );
ao22s80 g562627 ( .a(n_3093), .b(n_5292), .c(n_2483), .d(x_in_5_8), .o(n_9805) );
oa12f80 g562628 ( .a(n_6001), .b(n_5956), .c(x_in_3_8), .o(n_9690) );
ao22s80 g562629 ( .a(n_3246), .b(n_5298), .c(n_2501), .d(x_in_57_9), .o(n_9815) );
ao12f80 g562630 ( .a(n_6837), .b(n_5347), .c(n_5344), .o(n_5412) );
in01f80 g562631 ( .a(n_6616), .o(n_6617) );
oa12f80 g562632 ( .a(n_4750), .b(n_7700), .c(n_5745), .o(n_6616) );
oa12f80 g562633 ( .a(n_2997), .b(n_5756), .c(n_5905), .o(n_10845) );
in01f80 g562634 ( .a(n_6614), .o(n_6615) );
oa22f80 g562635 ( .a(n_3367), .b(n_5392), .c(n_6907), .d(n_6000), .o(n_6614) );
in01f80 g562636 ( .a(n_5998), .o(n_5999) );
oa12f80 g562637 ( .a(n_7697), .b(n_5958), .c(n_5757), .o(n_5998) );
oa12f80 g562638 ( .a(n_6808), .b(n_5297), .c(x_in_5_5), .o(n_5997) );
in01f80 g562639 ( .a(n_6612), .o(n_6613) );
ao22s80 g562640 ( .a(n_3410), .b(n_5304), .c(n_6814), .d(x_in_57_10), .o(n_6612) );
oa12f80 g562641 ( .a(n_3305), .b(n_5959), .c(n_6380), .o(n_9952) );
oa12f80 g562642 ( .a(n_4538), .b(n_2106), .c(n_5986), .o(n_11841) );
in01f80 g562643 ( .a(n_6610), .o(n_6611) );
oa12f80 g562644 ( .a(n_4590), .b(n_7679), .c(n_5962), .o(n_6610) );
ao22s80 g562645 ( .a(n_3319), .b(n_5411), .c(n_2426), .d(x_in_37_7), .o(n_10644) );
ao22s80 g562646 ( .a(n_3888), .b(n_5901), .c(n_3037), .d(x_in_21_9), .o(n_10631) );
ao12f80 g562647 ( .a(n_7605), .b(n_8295), .c(n_5742), .o(n_5410) );
in01f80 g562648 ( .a(n_6608), .o(n_6609) );
ao12f80 g562649 ( .a(n_4799), .b(n_7681), .c(x_in_37_8), .o(n_6608) );
in01f80 g562650 ( .a(n_5766), .o(n_5767) );
oa22f80 g562651 ( .a(n_3091), .b(n_5409), .c(n_5408), .d(n_4180), .o(n_5766) );
in01f80 g562652 ( .a(n_6606), .o(n_6607) );
ao22s80 g562653 ( .a(n_3594), .b(n_5270), .c(n_7076), .d(n_5271), .o(n_6606) );
ao12f80 g562654 ( .a(n_4818), .b(n_4817), .c(n_6405), .o(n_6410) );
in01f80 g562655 ( .a(n_6604), .o(n_6605) );
ao22s80 g562656 ( .a(n_3640), .b(n_5314), .c(n_6811), .d(x_in_57_11), .o(n_6604) );
in01f80 g562657 ( .a(n_6602), .o(n_6603) );
ao22s80 g562658 ( .a(n_3844), .b(n_5755), .c(n_7613), .d(x_in_5_11), .o(n_6602) );
ao12f80 g562659 ( .a(n_6898), .b(n_4869), .c(x_in_17_7), .o(n_9935) );
in01f80 g562660 ( .a(n_6600), .o(n_6601) );
ao22s80 g562661 ( .a(n_4081), .b(n_5290), .c(n_6805), .d(x_in_5_11), .o(n_6600) );
oa22f80 g562662 ( .a(n_4071), .b(n_5887), .c(n_7687), .d(n_5860), .o(n_10629) );
ao22s80 g562663 ( .a(n_7419), .b(n_2615), .c(n_5407), .d(x_in_41_12), .o(n_11229) );
oa12f80 g562664 ( .a(n_5088), .b(n_7683), .c(n_5872), .o(n_9800) );
oa22f80 g562665 ( .a(n_3645), .b(n_5740), .c(n_2898), .d(n_5884), .o(n_11434) );
in01f80 g562666 ( .a(n_5996), .o(n_8341) );
oa12f80 g562667 ( .a(n_5459), .b(n_5995), .c(n_6409), .o(n_5996) );
ao12f80 g562668 ( .a(n_5994), .b(n_5993), .c(n_3263), .o(n_7791) );
ao12f80 g562669 ( .a(n_4791), .b(n_2791), .c(x_in_21_7), .o(n_10627) );
no03m80 g562670 ( .a(n_3150), .b(n_4833), .c(x_in_41_1), .o(n_5406) );
ao12f80 g562671 ( .a(n_6878), .b(n_4816), .c(x_in_17_9), .o(n_9921) );
in01f80 g562672 ( .a(n_5404), .o(n_5405) );
oa12f80 g562673 ( .a(x_in_17_10), .b(n_4815), .c(n_5360), .o(n_5404) );
ao12f80 g562674 ( .a(n_4597), .b(n_3211), .c(x_in_21_11), .o(n_10636) );
oa12f80 g562675 ( .a(n_5992), .b(n_5991), .c(n_7790), .o(n_7782) );
ao22s80 g562676 ( .a(n_5482), .b(n_2634), .c(n_3757), .d(x_in_41_4), .o(n_11091) );
ao12f80 g562677 ( .a(n_5990), .b(n_5978), .c(n_7781), .o(n_7777) );
ao12f80 g562678 ( .a(n_6872), .b(n_4871), .c(x_in_17_11), .o(n_9903) );
oa22f80 g562679 ( .a(n_3092), .b(n_5989), .c(n_7707), .d(n_5914), .o(n_10625) );
oa22f80 g562680 ( .a(n_3914), .b(n_6200), .c(n_4403), .d(n_5988), .o(n_10746) );
oa12f80 g562681 ( .a(n_3031), .b(n_5727), .c(n_5963), .o(n_10823) );
ao12f80 g562682 ( .a(n_4814), .b(n_4813), .c(x_in_5_5), .o(n_7205) );
ao22s80 g562683 ( .a(n_3942), .b(n_5280), .c(n_2801), .d(n_6746), .o(n_12010) );
ao12f80 g562684 ( .a(n_5362), .b(n_4812), .c(x_in_17_4), .o(n_9871) );
in01f80 g562685 ( .a(n_6598), .o(n_6599) );
ao12f80 g562686 ( .a(n_4541), .b(n_7855), .c(n_5987), .o(n_6598) );
in01f80 g562687 ( .a(n_5402), .o(n_5403) );
oa12f80 g562688 ( .a(x_in_17_8), .b(n_4811), .c(n_5362), .o(n_5402) );
na02f80 g562689 ( .a(n_3890), .b(n_4033), .o(n_6956) );
oa12f80 g562690 ( .a(n_4365), .b(n_4364), .c(n_3323), .o(n_6406) );
in01f80 g562691 ( .a(n_6596), .o(n_6597) );
ao22s80 g562692 ( .a(n_3587), .b(n_5356), .c(n_6843), .d(n_10477), .o(n_6596) );
ao12f80 g562693 ( .a(n_8892), .b(n_6209), .c(n_4220), .o(n_7764) );
ao12f80 g562694 ( .a(n_8896), .b(n_4959), .c(n_4958), .o(n_8359) );
ao22s80 g562695 ( .a(n_3434), .b(n_5366), .c(n_6945), .d(n_5986), .o(n_10707) );
in01f80 g562696 ( .a(n_5984), .o(n_5985) );
oa12f80 g562697 ( .a(n_4632), .b(FE_OFN1234_n_4979), .c(n_5401), .o(n_5984) );
in01f80 g562698 ( .a(n_6594), .o(n_6595) );
ao22s80 g562699 ( .a(n_3652), .b(n_5284), .c(n_7051), .d(n_5293), .o(n_6594) );
oa22f80 g562700 ( .a(n_3316), .b(FE_OFN1202_n_5312), .c(n_4804), .d(x_in_27_4), .o(n_11690) );
in01f80 g562701 ( .a(n_6592), .o(n_6593) );
ao22s80 g562702 ( .a(n_3977), .b(n_5386), .c(n_7054), .d(n_5387), .o(n_6592) );
in01f80 g562703 ( .a(n_5400), .o(n_9098) );
ao12f80 g562704 ( .a(n_4814), .b(n_4872), .c(n_4813), .o(n_5400) );
in01f80 g562705 ( .a(n_5399), .o(n_9101) );
ao12f80 g562706 ( .a(n_4809), .b(n_4808), .c(n_4807), .o(n_5399) );
in01f80 g562707 ( .a(n_6590), .o(n_6591) );
ao12f80 g562708 ( .a(n_4806), .b(n_7754), .c(n_5939), .o(n_6590) );
oa12f80 g562709 ( .a(n_26869), .b(n_3462), .c(n_4903), .o(n_5398) );
oa12f80 g562710 ( .a(n_9426), .b(n_4646), .c(n_4645), .o(n_7918) );
no02f80 g562711 ( .a(n_3882), .b(n_6884), .o(n_5397) );
in01f80 g562712 ( .a(n_32735), .o(n_5983) );
in01f80 g562714 ( .a(n_5981), .o(n_11137) );
ao22s80 g562715 ( .a(n_5916), .b(n_2585), .c(n_5395), .d(x_in_41_5), .o(n_5981) );
oa22f80 g562716 ( .a(n_3103), .b(n_6760), .c(n_3752), .d(n_11409), .o(n_11131) );
in01f80 g562717 ( .a(n_5393), .o(n_5394) );
oa12f80 g562718 ( .a(n_4594), .b(n_6966), .c(n_4593), .o(n_5393) );
in01f80 g562719 ( .a(n_6588), .o(n_6589) );
ao22s80 g562720 ( .a(n_3639), .b(n_5980), .c(n_7757), .d(n_5979), .o(n_6588) );
ao22s80 g562721 ( .a(n_3139), .b(n_5338), .c(n_5339), .d(n_7138), .o(n_7634) );
oa22f80 g562722 ( .a(n_2637), .b(n_4916), .c(n_2046), .d(n_5095), .o(n_12829) );
ao22s80 g562723 ( .a(n_5453), .b(n_2561), .c(n_4068), .d(x_in_17_2), .o(n_11154) );
oa22f80 g562724 ( .a(n_3179), .b(n_5978), .c(n_2090), .d(n_4386), .o(n_10742) );
oa22f80 g562725 ( .a(n_6477), .b(n_7212), .c(n_7211), .d(n_5805), .o(n_9348) );
ao12f80 g562726 ( .a(n_3489), .b(n_4991), .c(n_4121), .o(n_26276) );
in01f80 g562727 ( .a(n_12692), .o(n_13093) );
oa22f80 g562728 ( .a(n_2962), .b(x_in_61_14), .c(n_2963), .d(n_4847), .o(n_12692) );
in01f80 g562729 ( .a(n_10142), .o(n_10144) );
oa12f80 g562730 ( .a(n_3625), .b(n_3624), .c(x_in_53_14), .o(n_10142) );
in01f80 g562731 ( .a(n_9687), .o(n_6587) );
ao22s80 g562732 ( .a(n_5957), .b(n_5963), .c(n_5958), .d(x_in_3_5), .o(n_9687) );
in01f80 g562733 ( .a(n_8526), .o(n_7761) );
oa12f80 g562734 ( .a(n_3790), .b(n_5391), .c(x_in_61_12), .o(n_8526) );
in01f80 g562735 ( .a(n_6585), .o(n_6586) );
oa12f80 g562736 ( .a(n_4693), .b(n_5232), .c(n_4692), .o(n_6585) );
oa22f80 g562737 ( .a(n_5753), .b(x_in_21_12), .c(n_5752), .d(n_5977), .o(n_7711) );
ao12f80 g562738 ( .a(n_5214), .b(n_5891), .c(n_5213), .o(n_8267) );
in01f80 g562739 ( .a(n_5975), .o(n_5976) );
ao12f80 g562740 ( .a(n_3960), .b(n_3959), .c(x_in_43_1), .o(n_5975) );
oa12f80 g562741 ( .a(n_3458), .b(n_3457), .c(x_in_59_1), .o(n_8614) );
oa22f80 g562742 ( .a(n_2990), .b(n_6000), .c(n_5392), .d(x_in_5_9), .o(n_6908) );
oa12f80 g562743 ( .a(n_3886), .b(n_5391), .c(n_3885), .o(n_12822) );
oa22f80 g562744 ( .a(n_5969), .b(n_5195), .c(n_5748), .d(n_5747), .o(n_7848) );
in01f80 g562745 ( .a(n_6470), .o(n_6471) );
oa12f80 g562746 ( .a(n_4214), .b(n_6437), .c(n_4213), .o(n_6470) );
in01f80 g562747 ( .a(n_6502), .o(n_9786) );
oa12f80 g562748 ( .a(n_3825), .b(n_3824), .c(x_in_59_5), .o(n_6502) );
ao12f80 g562749 ( .a(n_4252), .b(n_4251), .c(n_4250), .o(n_7858) );
in01f80 g562750 ( .a(n_6979), .o(n_9231) );
oa22f80 g562751 ( .a(n_2756), .b(x_in_43_8), .c(n_2757), .d(n_5501), .o(n_6979) );
in01f80 g562752 ( .a(n_7009), .o(n_9314) );
oa22f80 g562753 ( .a(n_5286), .b(x_in_35_3), .c(n_5287), .d(n_5390), .o(n_7009) );
in01f80 g562754 ( .a(FE_OFN482_n_13520), .o(n_5974) );
ao22s80 g562755 ( .a(n_2784), .b(n_7304), .c(n_2783), .d(x_in_7_8), .o(n_13520) );
in01f80 g562756 ( .a(FE_OFN478_n_11170), .o(n_12683) );
oa22f80 g562757 ( .a(n_2927), .b(x_in_7_4), .c(n_2928), .d(n_8522), .o(n_11170) );
oa22f80 g562758 ( .a(n_5814), .b(n_6584), .c(n_6583), .d(n_5813), .o(n_9357) );
ao22s80 g562759 ( .a(n_5674), .b(n_5868), .c(n_3376), .d(n_5866), .o(n_7148) );
ao22s80 g562760 ( .a(n_2983), .b(x_in_5_10), .c(n_5389), .d(n_5388), .o(n_6896) );
in01f80 g562761 ( .a(n_5972), .o(n_5973) );
oa12f80 g562762 ( .a(n_3931), .b(n_3930), .c(x_in_27_1), .o(n_5972) );
in01f80 g562763 ( .a(n_9577), .o(n_7705) );
oa22f80 g562764 ( .a(n_3183), .b(x_in_59_7), .c(n_3184), .d(n_5699), .o(n_9577) );
oa22f80 g562765 ( .a(n_6416), .b(n_3191), .c(n_5970), .d(x_in_49_9), .o(n_7633) );
in01f80 g562766 ( .a(n_13084), .o(n_13081) );
oa22f80 g562767 ( .a(n_2959), .b(x_in_7_14), .c(n_2960), .d(n_15590), .o(n_13084) );
ao12f80 g562768 ( .a(n_4169), .b(n_5918), .c(x_in_51_2), .o(n_8924) );
ao22s80 g562769 ( .a(n_2936), .b(n_5387), .c(n_5386), .d(x_in_11_4), .o(n_7055) );
in01f80 g562770 ( .a(n_12204), .o(n_10207) );
oa22f80 g562771 ( .a(n_5969), .b(n_5968), .c(n_5748), .d(x_in_7_6), .o(n_12204) );
in01f80 g562772 ( .a(n_11103), .o(n_9226) );
na02f80 g562773 ( .a(n_4344), .b(n_3541), .o(n_11103) );
oa12f80 g562774 ( .a(n_3585), .b(n_3584), .c(x_in_49_7), .o(n_6834) );
in01f80 g562775 ( .a(n_8020), .o(n_5967) );
oa12f80 g562776 ( .a(n_3972), .b(n_5367), .c(n_3971), .o(n_8020) );
oa22f80 g562777 ( .a(n_7598), .b(n_2507), .c(n_5385), .d(n_4000), .o(n_7097) );
in01f80 g562778 ( .a(n_8928), .o(n_8334) );
na02f80 g562779 ( .a(n_3609), .b(n_4896), .o(n_8928) );
in01f80 g562780 ( .a(n_6941), .o(n_9297) );
oa12f80 g562781 ( .a(n_3572), .b(n_3571), .c(x_in_59_14), .o(n_6941) );
in01f80 g562782 ( .a(n_5965), .o(n_5966) );
oa12f80 g562783 ( .a(n_3775), .b(n_3774), .c(n_3773), .o(n_5965) );
in01f80 g562784 ( .a(n_9437), .o(n_7400) );
no02f80 g562785 ( .a(n_4931), .b(n_4647), .o(n_9437) );
in01f80 g562786 ( .a(n_9592), .o(n_5964) );
oa12f80 g562787 ( .a(n_3937), .b(n_3936), .c(x_in_11_2), .o(n_9592) );
in01f80 g562788 ( .a(n_12147), .o(n_6582) );
ao22s80 g562789 ( .a(n_5762), .b(x_in_61_6), .c(n_5867), .d(n_5761), .o(n_12147) );
in01f80 g562790 ( .a(FE_OFN1190_n_13090), .o(n_6581) );
oa22f80 g562791 ( .a(n_8103), .b(n_7320), .c(n_3499), .d(x_in_7_9), .o(n_13090) );
oa12f80 g562792 ( .a(n_5788), .b(n_6580), .c(n_5039), .o(n_8368) );
in01f80 g562793 ( .a(n_6452), .o(n_6453) );
oa12f80 g562794 ( .a(n_4173), .b(n_4183), .c(n_4172), .o(n_6452) );
ao22s80 g562795 ( .a(n_5728), .b(n_5963), .c(n_5727), .d(x_in_3_5), .o(n_7666) );
in01f80 g562796 ( .a(n_6454), .o(n_6455) );
oa12f80 g562797 ( .a(n_4697), .b(n_4696), .c(n_5820), .o(n_6454) );
in01f80 g562798 ( .a(n_8514), .o(n_7784) );
oa22f80 g562799 ( .a(n_5278), .b(n_7402), .c(n_5279), .d(x_in_27_12), .o(n_8514) );
in01f80 g562800 ( .a(n_8597), .o(n_6579) );
oa22f80 g562801 ( .a(n_8650), .b(n_5761), .c(n_3378), .d(x_in_61_6), .o(n_8597) );
oa22f80 g562802 ( .a(n_5384), .b(n_2500), .c(n_2945), .d(n_5383), .o(n_6885) );
ao12f80 g562803 ( .a(n_4326), .b(n_5893), .c(n_4325), .o(n_7788) );
in01f80 g562804 ( .a(FE_OFN785_n_10198), .o(n_12152) );
oa22f80 g562805 ( .a(n_5163), .b(x_in_37_9), .c(n_4347), .d(n_5962), .o(n_10198) );
oa12f80 g562806 ( .a(n_4749), .b(n_4748), .c(n_5961), .o(n_10056) );
oa22f80 g562807 ( .a(n_4823), .b(n_5381), .c(n_2933), .d(x_in_41_4), .o(n_5382) );
in01f80 g562808 ( .a(n_8953), .o(n_7399) );
oa12f80 g562809 ( .a(n_5203), .b(n_5923), .c(x_in_53_12), .o(n_8953) );
oa22f80 g562810 ( .a(n_9157), .b(FE_OFN1152_n_3069), .c(n_162), .d(FE_OFN129_n_27449), .o(n_7398) );
na02f80 g562811 ( .a(n_5151), .b(n_4371), .o(n_9436) );
na02f80 g562812 ( .a(n_5063), .b(n_4528), .o(n_9419) );
ao22s80 g562813 ( .a(n_6435), .b(n_6425), .c(n_5132), .d(n_6434), .o(n_8677) );
oa22f80 g562814 ( .a(n_7396), .b(FE_OFN253_n_4280), .c(n_913), .d(FE_OFN136_n_27449), .o(n_7397) );
oa12f80 g562815 ( .a(n_4635), .b(n_4634), .c(n_5125), .o(n_7627) );
in01f80 g562816 ( .a(n_8518), .o(n_5960) );
ao22s80 g562817 ( .a(n_5375), .b(x_in_7_12), .c(n_5374), .d(n_7340), .o(n_8518) );
in01f80 g562818 ( .a(n_12637), .o(n_12613) );
oa12f80 g562819 ( .a(n_3456), .b(n_3455), .c(x_in_61_7), .o(n_12637) );
ao22s80 g562820 ( .a(n_3228), .b(n_5430), .c(n_5380), .d(x_in_23_2), .o(n_7157) );
in01f80 g562821 ( .a(n_9588), .o(n_6578) );
ao22s80 g562822 ( .a(n_5728), .b(n_5825), .c(n_5727), .d(x_in_3_3), .o(n_9588) );
in01f80 g562823 ( .a(n_8932), .o(n_8377) );
no02f80 g562824 ( .a(n_4753), .b(n_3992), .o(n_8932) );
ao22s80 g562825 ( .a(n_4627), .b(n_5378), .c(n_5377), .d(n_4626), .o(n_8167) );
oa12f80 g562826 ( .a(n_4758), .b(n_5928), .c(n_4757), .o(n_8762) );
ao12f80 g562827 ( .a(n_4726), .b(n_5850), .c(n_4725), .o(n_8791) );
oa22f80 g562828 ( .a(n_10385), .b(FE_OFN306_n_3069), .c(n_1580), .d(FE_OFN72_n_27012), .o(n_7228) );
in01f80 g562829 ( .a(n_9216), .o(n_6459) );
ao22s80 g562830 ( .a(n_5953), .b(n_5905), .c(n_5959), .d(x_in_3_9), .o(n_9216) );
in01f80 g562831 ( .a(n_7013), .o(n_9316) );
oa12f80 g562832 ( .a(n_3779), .b(n_3778), .c(x_in_27_3), .o(n_7013) );
ao12f80 g562833 ( .a(n_4561), .b(n_7815), .c(n_5931), .o(n_10148) );
oa22f80 g562834 ( .a(n_9167), .b(FE_OFN306_n_3069), .c(n_446), .d(FE_OFN357_n_4860), .o(n_7395) );
ao12f80 g562835 ( .a(n_3991), .b(n_4808), .c(x_in_0_1), .o(n_7103) );
oa12f80 g562836 ( .a(n_4671), .b(n_5922), .c(x_in_21_7), .o(n_7716) );
oa22f80 g562837 ( .a(n_5958), .b(x_in_3_7), .c(n_5957), .d(n_5757), .o(n_7698) );
in01f80 g562838 ( .a(n_6961), .o(n_9272) );
oa12f80 g562839 ( .a(n_3923), .b(n_3922), .c(x_in_3_14), .o(n_6961) );
oa22f80 g562840 ( .a(FE_OFN1250_n_5334), .b(n_5689), .c(n_5333), .d(x_in_51_13), .o(n_8511) );
oa22f80 g562841 ( .a(n_3303), .b(x_in_55_15), .c(n_3304), .d(n_5376), .o(n_8064) );
oa22f80 g562842 ( .a(n_9160), .b(FE_OFN257_n_4280), .c(n_882), .d(FE_OFN89_n_27449), .o(n_7227) );
ao22s80 g562843 ( .a(n_4624), .b(n_4920), .c(n_4919), .d(n_4623), .o(n_8145) );
ao22s80 g562844 ( .a(n_5375), .b(n_2869), .c(n_5374), .d(n_3789), .o(n_27794) );
ao22s80 g562845 ( .a(n_2692), .b(n_5373), .c(n_5372), .d(x_in_31_2), .o(n_7154) );
oa22f80 g562846 ( .a(n_5956), .b(x_in_3_10), .c(n_4124), .d(n_5666), .o(n_7646) );
in01f80 g562847 ( .a(n_11111), .o(n_12631) );
oa12f80 g562848 ( .a(n_4666), .b(n_5943), .c(x_in_21_9), .o(n_11111) );
ao12f80 g562849 ( .a(n_5035), .b(n_6577), .c(n_5034), .o(n_9116) );
ao12f80 g562850 ( .a(n_3619), .b(n_3618), .c(n_3617), .o(n_8190) );
ao12f80 g562851 ( .a(n_4161), .b(n_4160), .c(n_4159), .o(n_7745) );
in01f80 g562852 ( .a(n_6985), .o(n_5955) );
oa12f80 g562853 ( .a(n_3901), .b(n_3918), .c(x_in_53_4), .o(n_6985) );
oa22f80 g562854 ( .a(n_2909), .b(x_in_23_15), .c(n_2910), .d(n_5371), .o(n_8062) );
in01f80 g562855 ( .a(n_6915), .o(n_9291) );
oa22f80 g562856 ( .a(n_2930), .b(x_in_59_8), .c(n_2931), .d(n_5691), .o(n_6915) );
ao12f80 g562857 ( .a(n_3976), .b(n_3975), .c(n_7099), .o(n_5370) );
in01f80 g562858 ( .a(n_9672), .o(n_8312) );
oa22f80 g562859 ( .a(n_4941), .b(x_in_35_8), .c(n_4940), .d(n_4939), .o(n_9672) );
in01f80 g562860 ( .a(n_7135), .o(n_9340) );
oa12f80 g562861 ( .a(n_3574), .b(n_5269), .c(x_in_59_2), .o(n_7135) );
in01f80 g562862 ( .a(n_6917), .o(n_9293) );
oa22f80 g562863 ( .a(n_4944), .b(x_in_35_7), .c(n_4943), .d(n_4942), .o(n_6917) );
ao22s80 g562864 ( .a(n_2943), .b(n_4946), .c(n_4945), .d(x_in_15_2), .o(n_7163) );
in01f80 g562865 ( .a(n_6943), .o(n_9299) );
oa22f80 g562866 ( .a(n_5028), .b(x_in_35_6), .c(n_5027), .d(n_5369), .o(n_6943) );
in01f80 g562867 ( .a(n_9670), .o(n_7713) );
oa12f80 g562868 ( .a(n_3471), .b(n_5076), .c(x_in_35_5), .o(n_9670) );
in01f80 g562869 ( .a(n_8054), .o(n_5954) );
oa12f80 g562870 ( .a(n_3970), .b(n_3969), .c(n_3968), .o(n_8054) );
oa22f80 g562871 ( .a(n_2825), .b(x_in_15_15), .c(n_2826), .d(n_5368), .o(n_8072) );
in01f80 g562872 ( .a(n_9666), .o(n_7774) );
oa22f80 g562873 ( .a(n_2905), .b(x_in_35_4), .c(n_5367), .d(n_5987), .o(n_9666) );
ao22s80 g562874 ( .a(n_5953), .b(n_6380), .c(n_5959), .d(x_in_3_11), .o(n_7732) );
ao22s80 g562875 ( .a(n_4952), .b(n_4774), .c(n_4775), .d(n_4951), .o(n_8135) );
in01f80 g562876 ( .a(n_9662), .o(n_5951) );
ao12f80 g562877 ( .a(n_3544), .b(n_4956), .c(x_in_35_2), .o(n_9662) );
ao12f80 g562878 ( .a(n_3603), .b(n_3602), .c(x_in_35_1), .o(n_8668) );
in01f80 g562879 ( .a(n_8053), .o(n_5950) );
oa12f80 g562880 ( .a(n_3537), .b(n_3536), .c(n_3535), .o(n_8053) );
ao22s80 g562881 ( .a(n_2904), .b(n_5986), .c(n_5366), .d(x_in_45_2), .o(n_8457) );
ao12f80 g562882 ( .a(n_5162), .b(n_6576), .c(n_5161), .o(n_9423) );
in01f80 g562883 ( .a(n_8049), .o(n_5949) );
oa12f80 g562884 ( .a(n_3532), .b(n_3531), .c(n_3530), .o(n_8049) );
in01f80 g562885 ( .a(n_8919), .o(n_6575) );
no02f80 g562886 ( .a(n_4724), .b(n_3521), .o(n_8919) );
oa12f80 g562887 ( .a(n_3547), .b(n_3546), .c(n_3545), .o(n_8052) );
in01f80 g562888 ( .a(n_9279), .o(n_6574) );
ao22s80 g562889 ( .a(n_5758), .b(n_5757), .c(n_5756), .d(x_in_3_7), .o(n_9279) );
oa22f80 g562890 ( .a(n_5417), .b(n_2630), .c(n_3550), .d(n_5416), .o(n_7860) );
oa12f80 g562891 ( .a(n_3965), .b(n_3964), .c(n_3963), .o(n_8050) );
in01f80 g562892 ( .a(n_7017), .o(n_9233) );
oa22f80 g562893 ( .a(n_2920), .b(x_in_43_9), .c(n_2921), .d(n_7268), .o(n_7017) );
ao22s80 g562894 ( .a(n_2944), .b(n_5365), .c(n_5364), .d(x_in_47_2), .o(n_7160) );
in01f80 g562895 ( .a(n_8460), .o(n_8462) );
oa22f80 g562896 ( .a(n_5330), .b(n_6350), .c(n_5329), .d(x_in_51_6), .o(n_8460) );
oa22f80 g562897 ( .a(n_2711), .b(x_in_47_15), .c(n_2712), .d(n_5363), .o(n_8070) );
oa12f80 g562898 ( .a(n_5201), .b(n_5200), .c(n_5199), .o(n_10076) );
oa12f80 g562899 ( .a(n_4140), .b(n_4139), .c(n_4138), .o(n_8051) );
no03m80 g562900 ( .a(n_11201), .b(n_32729), .c(n_4825), .o(n_5948) );
ao12f80 g562901 ( .a(n_3962), .b(n_3961), .c(x_in_35_15), .o(n_8500) );
in01f80 g562902 ( .a(n_8022), .o(n_5947) );
oa12f80 g562903 ( .a(n_3956), .b(n_3955), .c(n_3954), .o(n_8022) );
in01f80 g562904 ( .a(n_8039), .o(n_8483) );
oa22f80 g562905 ( .a(n_2819), .b(n_4992), .c(n_4991), .d(x_in_59_12), .o(n_8039) );
in01f80 g562906 ( .a(n_6981), .o(n_8498) );
oa12f80 g562907 ( .a(n_3979), .b(n_5099), .c(n_3978), .o(n_6981) );
ao12f80 g562908 ( .a(n_5154), .b(n_6573), .c(n_5153), .o(n_8361) );
ao12f80 g562909 ( .a(n_4362), .b(n_4655), .c(x_in_37_3), .o(n_7894) );
oa22f80 g562910 ( .a(n_4941), .b(n_2073), .c(n_4940), .d(n_2072), .o(n_8073) );
in01f80 g562911 ( .a(n_8495), .o(n_5946) );
ao22s80 g562912 ( .a(n_4943), .b(n_2263), .c(n_4944), .d(n_2264), .o(n_8495) );
oa12f80 g562913 ( .a(n_3690), .b(n_8287), .c(x_in_17_4), .o(n_6510) );
in01f80 g562914 ( .a(n_8024), .o(n_5945) );
oa22f80 g562915 ( .a(n_5028), .b(n_2089), .c(n_5027), .d(n_2088), .o(n_8024) );
in01f80 g562916 ( .a(n_8493), .o(n_5865) );
ao12f80 g562917 ( .a(n_3559), .b(n_5076), .c(n_3558), .o(n_8493) );
in01f80 g562918 ( .a(n_8452), .o(n_7808) );
oa12f80 g562919 ( .a(n_3953), .b(n_3952), .c(x_in_7_1), .o(n_8452) );
in01f80 g562920 ( .a(n_8490), .o(n_5944) );
oa12f80 g562921 ( .a(n_3988), .b(n_4956), .c(n_3987), .o(n_8490) );
oa22f80 g562922 ( .a(n_6572), .b(n_5156), .c(n_5157), .d(x_in_35_1), .o(n_8660) );
in01f80 g562923 ( .a(n_6761), .o(n_6762) );
oa12f80 g562924 ( .a(n_4177), .b(n_4714), .c(n_4176), .o(n_6761) );
ao12f80 g562925 ( .a(n_4335), .b(n_5943), .c(x_in_21_13), .o(n_7694) );
in01f80 g562926 ( .a(n_6887), .o(n_9289) );
oa22f80 g562927 ( .a(n_2919), .b(x_in_35_9), .c(n_5099), .d(n_5098), .o(n_6887) );
ao12f80 g562928 ( .a(n_5050), .b(n_5049), .c(n_5048), .o(n_9179) );
ao22s80 g562929 ( .a(n_2951), .b(x_in_17_3), .c(n_5669), .d(n_2520), .o(n_6850) );
ao22s80 g562930 ( .a(n_3240), .b(x_in_17_5), .c(n_4868), .d(n_9646), .o(n_6930) );
ao22s80 g562931 ( .a(n_4812), .b(x_in_17_6), .c(n_3317), .d(n_5362), .o(n_6870) );
ao22s80 g562932 ( .a(n_3067), .b(x_in_17_7), .c(n_4869), .d(n_9651), .o(n_6899) );
oa12f80 g562933 ( .a(n_3528), .b(n_4820), .c(n_3527), .o(n_7194) );
ao22s80 g562934 ( .a(n_2976), .b(x_in_57_7), .c(n_5361), .d(n_4055), .o(n_6890) );
ao22s80 g562935 ( .a(n_2947), .b(x_in_17_8), .c(n_4811), .d(n_5360), .o(n_6847) );
ao22s80 g562936 ( .a(n_2774), .b(x_in_17_9), .c(n_4816), .d(n_9654), .o(n_6879) );
oa22f80 g562937 ( .a(n_4815), .b(n_5359), .c(n_3032), .d(x_in_17_10), .o(n_6902) );
ao22s80 g562938 ( .a(n_3180), .b(x_in_17_11), .c(n_4871), .d(n_5418), .o(n_6873) );
in01f80 g562939 ( .a(n_7769), .o(n_9643) );
oa22f80 g562940 ( .a(n_5858), .b(x_in_19_8), .c(n_5859), .d(n_5554), .o(n_7769) );
in01f80 g562941 ( .a(n_6936), .o(n_6427) );
oa22f80 g562942 ( .a(n_5358), .b(x_in_17_13), .c(n_5357), .d(n_10477), .o(n_6936) );
in01f80 g562943 ( .a(n_7802), .o(n_9645) );
oa22f80 g562944 ( .a(n_5936), .b(x_in_19_9), .c(n_5937), .d(n_5537), .o(n_7802) );
in01f80 g562945 ( .a(n_7823), .o(n_9641) );
oa22f80 g562946 ( .a(n_5942), .b(x_in_19_7), .c(n_5941), .d(n_5940), .o(n_7823) );
in01f80 g562947 ( .a(n_7796), .o(n_9637) );
oa22f80 g562948 ( .a(n_5876), .b(x_in_19_6), .c(n_5877), .d(n_5326), .o(n_7796) );
in01f80 g562949 ( .a(n_7850), .o(n_9635) );
oa12f80 g562950 ( .a(n_4886), .b(n_5934), .c(x_in_19_5), .o(n_7850) );
in01f80 g562951 ( .a(n_7899), .o(n_9633) );
oa22f80 g562952 ( .a(n_5933), .b(x_in_19_4), .c(n_5932), .d(n_5939), .o(n_7899) );
ao22s80 g562953 ( .a(n_5356), .b(x_in_17_13), .c(n_2946), .d(n_10477), .o(n_6844) );
oa22f80 g562954 ( .a(n_2913), .b(x_in_31_15), .c(n_2914), .d(n_5355), .o(n_8059) );
ao22s80 g562955 ( .a(n_4248), .b(n_5354), .c(n_5353), .d(n_4247), .o(n_8125) );
in01f80 g562956 ( .a(n_7041), .o(n_9263) );
oa12f80 g562957 ( .a(n_3621), .b(n_3620), .c(x_in_19_14), .o(n_7041) );
oa12f80 g562958 ( .a(n_3999), .b(n_3998), .c(n_4759), .o(n_7198) );
in01f80 g562959 ( .a(n_7005), .o(n_9309) );
oa22f80 g562960 ( .a(n_3226), .b(x_in_11_8), .c(n_3227), .d(n_5352), .o(n_7005) );
ao12f80 g562961 ( .a(n_4699), .b(n_5928), .c(n_4698), .o(n_7925) );
ao22s80 g562962 ( .a(n_2942), .b(n_5351), .c(n_5350), .d(x_in_63_2), .o(n_7151) );
oa12f80 g562963 ( .a(n_4701), .b(n_4700), .c(n_5938), .o(n_7767) );
ao22s80 g562964 ( .a(n_5937), .b(n_2511), .c(n_5936), .d(n_3781), .o(n_7833) );
oa22f80 g562965 ( .a(n_2911), .b(x_in_63_15), .c(n_2912), .d(n_5042), .o(n_8068) );
ao22s80 g562966 ( .a(n_5941), .b(n_2678), .c(n_5942), .d(n_3849), .o(n_7829) );
in01f80 g562967 ( .a(n_8046), .o(n_5935) );
ao12f80 g562968 ( .a(n_3401), .b(n_3400), .c(n_3399), .o(n_8046) );
ao12f80 g562969 ( .a(n_4665), .b(n_5934), .c(n_4664), .o(n_7825) );
ao22s80 g562970 ( .a(n_5349), .b(n_4779), .c(n_4780), .d(n_5348), .o(n_8123) );
oa22f80 g562971 ( .a(n_5933), .b(n_3838), .c(n_5932), .d(n_3415), .o(n_7821) );
ao22s80 g562972 ( .a(n_3381), .b(n_5931), .c(n_5930), .d(x_in_3_4), .o(n_7749) );
ao12f80 g562973 ( .a(n_5075), .b(n_5854), .c(n_5074), .o(n_8956) );
ao22s80 g562974 ( .a(n_5347), .b(n_5346), .c(n_5345), .d(n_5344), .o(n_6838) );
ao12f80 g562975 ( .a(n_3924), .b(n_5261), .c(n_5342), .o(n_8285) );
ao12f80 g562976 ( .a(n_4981), .b(n_6571), .c(n_4980), .o(n_9427) );
in01f80 g562977 ( .a(n_10042), .o(n_6570) );
oa12f80 g562978 ( .a(n_4754), .b(n_5824), .c(n_5929), .o(n_10042) );
in01f80 g562979 ( .a(n_8908), .o(n_6569) );
oa12f80 g562980 ( .a(n_4622), .b(n_5928), .c(n_4621), .o(n_8908) );
ao22s80 g562981 ( .a(n_3012), .b(n_5339), .c(n_5338), .d(n_3138), .o(n_7139) );
oa12f80 g562982 ( .a(n_4752), .b(n_4751), .c(x_in_1_3), .o(n_7967) );
ao22s80 g562983 ( .a(n_6750), .b(n_4317), .c(n_5443), .d(n_5337), .o(n_6704) );
in01f80 g562984 ( .a(n_8037), .o(n_5927) );
oa12f80 g562985 ( .a(n_3474), .b(n_3473), .c(n_3472), .o(n_8037) );
ao22s80 g562986 ( .a(n_3630), .b(n_5926), .c(n_5925), .d(x_in_13_12), .o(n_8903) );
oa12f80 g562987 ( .a(n_4292), .b(n_4615), .c(n_4291), .o(n_7391) );
in01f80 g562988 ( .a(n_9618), .o(n_5924) );
oa12f80 g562989 ( .a(n_3829), .b(n_3828), .c(n_3827), .o(n_9618) );
ao22s80 g562990 ( .a(n_2941), .b(n_5336), .c(n_5335), .d(x_in_55_2), .o(n_6505) );
in01f80 g562991 ( .a(n_7178), .o(n_9257) );
oa22f80 g562992 ( .a(n_4841), .b(x_in_51_8), .c(n_3347), .d(n_6351), .o(n_7178) );
in01f80 g562993 ( .a(n_9258), .o(n_7968) );
oa22f80 g562994 ( .a(FE_OFN1250_n_5334), .b(x_in_51_9), .c(n_5333), .d(n_5332), .o(n_9258) );
oa22f80 g562995 ( .a(n_5706), .b(n_4143), .c(n_5705), .d(x_in_61_2), .o(n_8545) );
in01f80 g562996 ( .a(n_7184), .o(n_9255) );
oa22f80 g562997 ( .a(n_5325), .b(x_in_51_7), .c(n_5324), .d(n_5331), .o(n_7184) );
in01f80 g562998 ( .a(n_7726), .o(n_9253) );
oa22f80 g562999 ( .a(n_4899), .b(x_in_51_6), .c(FE_OFN931_n_4898), .d(n_6350), .o(n_7726) );
in01f80 g563000 ( .a(n_7182), .o(n_9792) );
oa12f80 g563001 ( .a(n_3893), .b(n_4927), .c(x_in_51_5), .o(n_7182) );
ao22s80 g563002 ( .a(n_3496), .b(n_5988), .c(n_5923), .d(x_in_53_13), .o(n_8927) );
in01f80 g563003 ( .a(n_10188), .o(n_12165) );
oa22f80 g563004 ( .a(n_5922), .b(x_in_21_3), .c(n_3430), .d(n_6781), .o(n_10188) );
in01f80 g563005 ( .a(n_9246), .o(n_7721) );
oa22f80 g563006 ( .a(n_4901), .b(x_in_51_4), .c(FE_OFN1246_n_4900), .d(n_5979), .o(n_9246) );
in01f80 g563007 ( .a(n_9620), .o(n_7970) );
oa12f80 g563008 ( .a(n_4114), .b(n_4936), .c(x_in_51_3), .o(n_9620) );
oa22f80 g563009 ( .a(n_5330), .b(x_in_51_2), .c(n_5329), .d(n_2490), .o(n_9249) );
in01f80 g563010 ( .a(n_5919), .o(n_5920) );
ao12f80 g563011 ( .a(n_3967), .b(n_3966), .c(n_4903), .o(n_5919) );
oa22f80 g563012 ( .a(n_5808), .b(n_6508), .c(n_6507), .d(n_5807), .o(n_9350) );
ao22s80 g563013 ( .a(n_3793), .b(n_4932), .c(n_2932), .d(x_in_51_1), .o(n_7428) );
ao12f80 g563014 ( .a(n_4743), .b(n_5918), .c(n_4742), .o(n_7427) );
oa22f80 g563015 ( .a(n_5732), .b(x_in_3_8), .c(n_3575), .d(n_5524), .o(n_7656) );
oa12f80 g563016 ( .a(n_3654), .b(n_3653), .c(x_in_49_8), .o(n_6868) );
ao12f80 g563017 ( .a(n_3913), .b(n_3912), .c(x_in_49_10), .o(n_6836) );
ao12f80 g563018 ( .a(n_3727), .b(n_3726), .c(x_in_49_6), .o(n_6861) );
ao22s80 g563019 ( .a(n_3251), .b(x_in_49_5), .c(n_3250), .d(n_5095), .o(n_6793) );
ao12f80 g563020 ( .a(n_3926), .b(n_3925), .c(x_in_49_4), .o(n_6832) );
in01f80 g563021 ( .a(n_7145), .o(n_5917) );
oa12f80 g563022 ( .a(n_3614), .b(n_3613), .c(x_in_49_3), .o(n_7145) );
in01f80 g563023 ( .a(n_6993), .o(n_9276) );
oa22f80 g563024 ( .a(n_3231), .b(x_in_27_7), .c(n_3232), .d(n_5680), .o(n_6993) );
oa12f80 g563025 ( .a(n_4337), .b(n_4598), .c(n_4336), .o(n_8936) );
in01f80 g563026 ( .a(n_8421), .o(n_8425) );
oa22f80 g563027 ( .a(n_3013), .b(n_6420), .c(n_3014), .d(x_in_51_12), .o(n_8421) );
ao22s80 g563028 ( .a(n_2793), .b(x_in_13_1), .c(n_5328), .d(n_2707), .o(n_7167) );
oa12f80 g563029 ( .a(n_5206), .b(n_5205), .c(n_5204), .o(n_9354) );
oa22f80 g563030 ( .a(n_6959), .b(n_2111), .c(n_6958), .d(n_2110), .o(n_10088) );
ao12f80 g563031 ( .a(n_4014), .b(n_4916), .c(n_4013), .o(n_7062) );
oa12f80 g563032 ( .a(n_4555), .b(n_4554), .c(n_5126), .o(n_7878) );
ao12f80 g563033 ( .a(n_4324), .b(n_5916), .c(n_4323), .o(n_14988) );
in01f80 g563034 ( .a(n_6567), .o(n_6568) );
oa12f80 g563035 ( .a(n_4637), .b(n_4638), .c(n_4636), .o(n_6567) );
oa12f80 g563036 ( .a(n_4600), .b(n_4599), .c(n_5107), .o(n_8951) );
oa22f80 g563037 ( .a(n_5989), .b(x_in_21_6), .c(n_5915), .d(n_5914), .o(n_7708) );
oa12f80 g563038 ( .a(n_4607), .b(n_4606), .c(n_4605), .o(n_7625) );
in01f80 g563039 ( .a(n_6976), .o(n_8475) );
oa22f80 g563040 ( .a(n_5325), .b(n_8420), .c(n_5324), .d(x_in_51_11), .o(n_6976) );
ao12f80 g563041 ( .a(n_5110), .b(n_5109), .c(n_5108), .o(n_8281) );
in01f80 g563042 ( .a(n_8015), .o(n_6566) );
ao12f80 g563043 ( .a(n_4620), .b(n_5913), .c(n_4997), .o(n_8015) );
oa12f80 g563044 ( .a(n_4644), .b(n_4643), .c(n_4642), .o(n_8950) );
oa12f80 g563045 ( .a(n_3881), .b(n_3880), .c(n_3879), .o(n_6911) );
in01f80 g563046 ( .a(n_8083), .o(n_8467) );
oa22f80 g563047 ( .a(n_4927), .b(n_5332), .c(n_3159), .d(x_in_51_9), .o(n_8083) );
in01f80 g563048 ( .a(n_9598), .o(n_8988) );
oa12f80 g563049 ( .a(n_3941), .b(n_3940), .c(x_in_27_2), .o(n_9598) );
ao12f80 g563050 ( .a(n_3534), .b(n_3533), .c(n_7102), .o(n_5323) );
oa22f80 g563051 ( .a(n_4901), .b(n_6351), .c(FE_OFN1246_n_4900), .d(x_in_51_8), .o(n_8465) );
in01f80 g563052 ( .a(n_8542), .o(n_6565) );
oa22f80 g563053 ( .a(n_8477), .b(n_4602), .c(n_7581), .d(n_3027), .o(n_8542) );
in01f80 g563054 ( .a(n_8117), .o(n_8464) );
oa22f80 g563055 ( .a(n_4936), .b(n_5331), .c(n_3182), .d(x_in_51_7), .o(n_8117) );
in01f80 g563056 ( .a(n_8891), .o(n_6564) );
ao12f80 g563057 ( .a(n_4619), .b(n_6204), .c(n_4618), .o(n_8891) );
oa22f80 g563058 ( .a(n_5750), .b(x_in_37_9), .c(n_5749), .d(n_5962), .o(n_8859) );
in01f80 g563059 ( .a(FE_OFN484_n_12038), .o(n_5912) );
oa22f80 g563060 ( .a(n_2893), .b(x_in_7_9), .c(n_2894), .d(n_7320), .o(n_12038) );
in01f80 g563061 ( .a(n_12209), .o(n_12149) );
oa12f80 g563062 ( .a(n_3578), .b(n_3577), .c(x_in_37_14), .o(n_12209) );
in01f80 g563063 ( .a(n_5910), .o(n_5911) );
oa12f80 g563064 ( .a(n_3515), .b(n_4793), .c(n_5226), .o(n_5910) );
oa12f80 g563065 ( .a(n_4137), .b(n_5322), .c(n_4768), .o(n_7130) );
in01f80 g563066 ( .a(n_7028), .o(n_9323) );
oa12f80 g563067 ( .a(n_4085), .b(n_4084), .c(x_in_11_5), .o(n_7028) );
in01f80 g563068 ( .a(n_8458), .o(n_5909) );
oa22f80 g563069 ( .a(n_3270), .b(n_4948), .c(n_3518), .d(n_9295), .o(n_8458) );
ao22s80 g563070 ( .a(n_5908), .b(n_4782), .c(n_4783), .d(n_5907), .o(n_10761) );
in01f80 g563071 ( .a(n_25699), .o(n_24693) );
ao12f80 g563072 ( .a(n_4207), .b(n_4206), .c(n_4205), .o(n_25699) );
in01f80 g563073 ( .a(n_9617), .o(n_7810) );
oa12f80 g563074 ( .a(n_3974), .b(FE_OFN933_n_4950), .c(x_in_51_15), .o(n_9617) );
in01f80 g563075 ( .a(n_8344), .o(n_7389) );
na02f80 g563076 ( .a(n_4918), .b(n_4152), .o(n_8344) );
oa12f80 g563077 ( .a(n_9424), .b(n_4609), .c(n_4608), .o(n_7739) );
ao12f80 g563078 ( .a(n_5131), .b(n_6563), .c(n_5130), .o(n_9425) );
ao22s80 g563079 ( .a(n_4683), .b(n_5321), .c(n_5320), .d(n_5319), .o(n_6829) );
oa12f80 g563080 ( .a(n_3939), .b(n_3938), .c(x_in_9_15), .o(n_7047) );
in01f80 g563081 ( .a(n_9016), .o(n_12179) );
oa22f80 g563082 ( .a(n_5753), .b(x_in_21_8), .c(n_5752), .d(n_5860), .o(n_9016) );
ao12f80 g563083 ( .a(n_3910), .b(n_3909), .c(x_in_57_3), .o(n_7173) );
in01f80 g563084 ( .a(n_12575), .o(n_6562) );
oa22f80 g563085 ( .a(n_5706), .b(n_5839), .c(n_5705), .d(x_in_61_7), .o(n_12575) );
in01f80 g563086 ( .a(n_8510), .o(n_7845) );
oa12f80 g563087 ( .a(n_3908), .b(n_3907), .c(x_in_61_1), .o(n_8510) );
oa22f80 g563088 ( .a(n_4960), .b(n_5446), .c(n_5436), .d(n_2238), .o(n_7870) );
in01f80 g563089 ( .a(n_5906), .o(n_11140) );
ao22s80 g563090 ( .a(n_5685), .b(n_2642), .c(n_4955), .d(x_in_41_7), .o(n_5906) );
in01f80 g563091 ( .a(n_6561), .o(n_12937) );
ao22s80 g563092 ( .a(n_7475), .b(n_3648), .c(n_5407), .d(x_in_41_9), .o(n_6561) );
in01f80 g563093 ( .a(n_6995), .o(n_9305) );
oa12f80 g563094 ( .a(n_4026), .b(n_4025), .c(x_in_43_5), .o(n_6995) );
ao22s80 g563095 ( .a(n_5758), .b(n_5905), .c(n_5756), .d(x_in_3_9), .o(n_7670) );
in01f80 g563096 ( .a(n_12628), .o(n_9013) );
oa12f80 g563097 ( .a(n_4517), .b(n_5751), .c(x_in_21_7), .o(n_12628) );
ao22s80 g563098 ( .a(n_4965), .b(n_4393), .c(n_4394), .d(n_4964), .o(n_8131) );
in01f80 g563099 ( .a(n_8860), .o(n_6560) );
oa12f80 g563100 ( .a(n_4254), .b(n_5855), .c(n_4253), .o(n_8860) );
in01f80 g563101 ( .a(n_8534), .o(n_6559) );
ao12f80 g563102 ( .a(n_4235), .b(n_4629), .c(n_5904), .o(n_8534) );
in01f80 g563103 ( .a(n_6462), .o(n_6463) );
oa12f80 g563104 ( .a(n_4673), .b(n_7419), .c(n_4672), .o(n_6462) );
in01f80 g563105 ( .a(FE_OFN1200_n_10340), .o(n_12625) );
oa22f80 g563106 ( .a(n_5903), .b(x_in_21_6), .c(n_5870), .d(n_5914), .o(n_10340) );
ao22s80 g563107 ( .a(FE_OFN726_n_5240), .b(n_4984), .c(n_5241), .d(n_4800), .o(n_8753) );
in01f80 g563108 ( .a(n_8910), .o(n_5768) );
ao12f80 g563109 ( .a(n_3797), .b(FE_OFN1234_n_4979), .c(n_3796), .o(n_8910) );
ao12f80 g563110 ( .a(n_3520), .b(n_4872), .c(x_in_4_1), .o(n_7100) );
in01f80 g563111 ( .a(n_7869), .o(n_6558) );
oa12f80 g563112 ( .a(n_4728), .b(n_4727), .c(x_in_45_15), .o(n_7869) );
ao12f80 g563113 ( .a(n_3862), .b(FE_OFN845_n_7616), .c(n_4604), .o(n_8014) );
oa22f80 g563114 ( .a(n_2940), .b(x_in_25_12), .c(n_5318), .d(n_5317), .o(n_7080) );
oa12f80 g563115 ( .a(n_4012), .b(n_5215), .c(n_4011), .o(n_8017) );
oa12f80 g563116 ( .a(n_3371), .b(n_4821), .c(x_in_25_9), .o(n_7071) );
oa22f80 g563117 ( .a(n_2725), .b(x_in_25_8), .c(n_5316), .d(n_3129), .o(n_7074) );
oa22f80 g563118 ( .a(n_3028), .b(x_in_25_7), .c(n_5315), .d(n_3132), .o(n_7083) );
oa22f80 g563119 ( .a(n_2925), .b(x_in_25_6), .c(n_5057), .d(n_3771), .o(n_7089) );
ao22s80 g563120 ( .a(n_3290), .b(n_4593), .c(n_4594), .d(x_in_25_5), .o(n_6967) );
ao12f80 g563121 ( .a(n_4711), .b(n_4710), .c(n_5902), .o(n_7799) );
ao12f80 g563122 ( .a(n_3478), .b(n_5701), .c(n_5700), .o(n_8789) );
ao22s80 g563123 ( .a(n_2958), .b(x_in_57_11), .c(n_5314), .d(n_5313), .o(n_6812) );
in01f80 g563124 ( .a(n_6556), .o(n_6557) );
oa12f80 g563125 ( .a(n_4204), .b(n_5223), .c(n_4203), .o(n_6556) );
in01f80 g563126 ( .a(n_6554), .o(n_6555) );
oa22f80 g563127 ( .a(n_5774), .b(x_in_45_12), .c(n_3562), .d(n_10486), .o(n_6554) );
ao22s80 g563128 ( .a(FE_OFN1202_n_5312), .b(n_5679), .c(n_2818), .d(x_in_27_4), .o(n_7049) );
oa22f80 g563129 ( .a(n_4819), .b(n_5311), .c(n_2745), .d(x_in_25_13), .o(n_7125) );
ao12f80 g563130 ( .a(n_3861), .b(n_3860), .c(n_3859), .o(n_25405) );
in01f80 g563131 ( .a(FE_OFN1198_n_13003), .o(n_6553) );
ao22s80 g563132 ( .a(n_5901), .b(n_5900), .c(n_5890), .d(x_in_21_5), .o(n_13003) );
in01f80 g563133 ( .a(n_6551), .o(n_6552) );
oa12f80 g563134 ( .a(n_4262), .b(n_5225), .c(n_5228), .o(n_6551) );
ao22s80 g563135 ( .a(n_12697), .b(n_2283), .c(n_10779), .d(n_2855), .o(n_8710) );
in01f80 g563136 ( .a(n_8066), .o(n_5899) );
oa12f80 g563137 ( .a(n_4005), .b(n_5701), .c(n_4004), .o(n_8066) );
in01f80 g563138 ( .a(n_8048), .o(n_5898) );
ao12f80 g563139 ( .a(n_3948), .b(n_3947), .c(n_3946), .o(n_8048) );
in01f80 g563140 ( .a(n_6989), .o(n_9307) );
oa22f80 g563141 ( .a(n_3217), .b(x_in_27_4), .c(n_3218), .d(n_5679), .o(n_6989) );
in01f80 g563142 ( .a(n_8879), .o(n_6550) );
ao22s80 g563143 ( .a(n_12697), .b(n_2734), .c(n_10779), .d(n_4801), .o(n_8879) );
in01f80 g563144 ( .a(n_8045), .o(n_5897) );
oa12f80 g563145 ( .a(n_3466), .b(n_3465), .c(n_3464), .o(n_8045) );
in01f80 g563146 ( .a(n_8043), .o(n_5896) );
ao12f80 g563147 ( .a(n_3945), .b(n_3944), .c(n_3943), .o(n_8043) );
in01f80 g563148 ( .a(n_8528), .o(n_8898) );
oa22f80 g563149 ( .a(n_6434), .b(n_2372), .c(n_6425), .d(n_2273), .o(n_8528) );
in01f80 g563150 ( .a(n_8035), .o(n_5895) );
oa12f80 g563151 ( .a(n_3565), .b(n_3564), .c(n_3563), .o(n_8035) );
in01f80 g563152 ( .a(n_8030), .o(n_5894) );
oa12f80 g563153 ( .a(n_3929), .b(n_3928), .c(n_3927), .o(n_8030) );
oa12f80 g563154 ( .a(n_3951), .b(n_3950), .c(n_3949), .o(n_8031) );
in01f80 g563155 ( .a(n_8811), .o(n_6549) );
oa22f80 g563156 ( .a(n_3677), .b(x_in_25_12), .c(n_3676), .d(n_5317), .o(n_8811) );
in01f80 g563157 ( .a(n_7045), .o(n_9332) );
oa22f80 g563158 ( .a(n_3213), .b(x_in_11_9), .c(n_3214), .d(n_5310), .o(n_7045) );
ao22s80 g563159 ( .a(n_5885), .b(n_5849), .c(n_5886), .d(x_in_37_12), .o(n_8855) );
in01f80 g563160 ( .a(n_7032), .o(n_9238) );
oa22f80 g563161 ( .a(n_2902), .b(x_in_11_7), .c(n_2903), .d(n_5089), .o(n_7032) );
in01f80 g563162 ( .a(n_11120), .o(n_12619) );
oa22f80 g563163 ( .a(n_5989), .b(x_in_21_2), .c(n_5915), .d(n_7434), .o(n_11120) );
in01f80 g563164 ( .a(n_7030), .o(n_9325) );
oa22f80 g563165 ( .a(n_2717), .b(x_in_11_6), .c(n_2718), .d(n_5309), .o(n_7030) );
oa12f80 g563166 ( .a(n_3539), .b(n_3538), .c(n_5308), .o(n_7094) );
in01f80 g563167 ( .a(FE_OFN1226_n_10183), .o(n_12157) );
oa22f80 g563168 ( .a(n_5750), .b(x_in_37_5), .c(n_5749), .d(n_5742), .o(n_10183) );
oa12f80 g563169 ( .a(n_5193), .b(n_5831), .c(n_5192), .o(n_8366) );
oa12f80 g563170 ( .a(n_3549), .b(n_3548), .c(n_4352), .o(n_7107) );
oa12f80 g563171 ( .a(n_3982), .b(n_3981), .c(n_4716), .o(n_7121) );
oa12f80 g563172 ( .a(n_3984), .b(n_3983), .c(n_4720), .o(n_7119) );
oa12f80 g563173 ( .a(n_3523), .b(n_3522), .c(n_4155), .o(n_7117) );
oa12f80 g563174 ( .a(n_3525), .b(n_3524), .c(n_4719), .o(n_7123) );
ao12f80 g563175 ( .a(n_3986), .b(n_3985), .c(n_4722), .o(n_7021) );
in01f80 g563176 ( .a(n_8455), .o(n_8881) );
oa12f80 g563177 ( .a(n_4708), .b(n_4760), .c(n_4707), .o(n_8455) );
in01f80 g563178 ( .a(n_7026), .o(n_9321) );
oa22f80 g563179 ( .a(n_2917), .b(x_in_11_4), .c(n_2918), .d(n_5387), .o(n_7026) );
ao12f80 g563180 ( .a(n_4133), .b(n_4132), .c(n_8191), .o(n_8588) );
in01f80 g563181 ( .a(n_7038), .o(n_9319) );
oa12f80 g563182 ( .a(n_3514), .b(n_3513), .c(x_in_11_3), .o(n_7038) );
in01f80 g563183 ( .a(n_7862), .o(n_9265) );
oa22f80 g563184 ( .a(n_4024), .b(x_in_19_3), .c(n_5893), .d(n_5252), .o(n_7862) );
oa22f80 g563185 ( .a(n_5307), .b(n_4668), .c(n_4669), .d(x_in_57_5), .o(n_7187) );
ao12f80 g563186 ( .a(n_3904), .b(n_5306), .c(x_in_57_6), .o(n_6939) );
ao12f80 g563187 ( .a(n_3905), .b(n_5305), .c(x_in_57_8), .o(n_6893) );
ao22s80 g563188 ( .a(n_2965), .b(x_in_57_10), .c(n_5304), .d(n_3409), .o(n_6815) );
ao22s80 g563189 ( .a(n_2954), .b(x_in_57_12), .c(n_5303), .d(n_5302), .o(n_6882) );
in01f80 g563190 ( .a(n_8448), .o(n_7819) );
oa22f80 g563191 ( .a(n_5026), .b(n_5025), .c(n_5024), .d(x_in_11_12), .o(n_8448) );
oa22f80 g563192 ( .a(n_9163), .b(FE_OFN292_n_3069), .c(n_761), .d(FE_OFN95_n_27449), .o(n_7387) );
in01f80 g563193 ( .a(n_8613), .o(n_6548) );
oa22f80 g563194 ( .a(n_5892), .b(n_3845), .c(n_5891), .d(n_5046), .o(n_8613) );
in01f80 g563195 ( .a(n_7060), .o(n_9235) );
oa12f80 g563196 ( .a(n_3935), .b(n_3934), .c(x_in_11_14), .o(n_7060) );
ao22s80 g563197 ( .a(n_4662), .b(x_in_25_3), .c(n_5704), .d(n_5703), .o(n_8106) );
oa22f80 g563198 ( .a(n_5890), .b(x_in_21_9), .c(n_5901), .d(n_3887), .o(n_7691) );
no02f80 g563199 ( .a(n_4357), .b(n_5054), .o(n_9403) );
ao22s80 g563200 ( .a(n_5024), .b(n_3389), .c(n_5026), .d(n_3806), .o(n_26273) );
in01f80 g563201 ( .a(n_7180), .o(n_9248) );
oa12f80 g563202 ( .a(n_3487), .b(n_3486), .c(x_in_51_14), .o(n_7180) );
oa22f80 g563203 ( .a(n_5298), .b(n_3245), .c(n_2964), .d(x_in_57_9), .o(n_6818) );
ao22s80 g563204 ( .a(FE_OFN726_n_5240), .b(n_4574), .c(n_5241), .d(n_2373), .o(n_6905) );
in01f80 g563205 ( .a(n_6546), .o(n_6547) );
oa12f80 g563206 ( .a(n_4690), .b(n_5227), .c(n_5224), .o(n_6546) );
oa12f80 g563207 ( .a(n_3356), .b(n_3355), .c(n_3354), .o(n_8055) );
in01f80 g563208 ( .a(n_8538), .o(n_6545) );
ao22s80 g563209 ( .a(n_5889), .b(n_5127), .c(n_5476), .d(n_2378), .o(n_8538) );
in01f80 g563210 ( .a(n_6987), .o(n_9240) );
oa22f80 g563211 ( .a(n_3029), .b(x_in_43_7), .c(n_3030), .d(n_5519), .o(n_6987) );
in01f80 g563212 ( .a(n_7746), .o(n_9251) );
oa22f80 g563213 ( .a(n_2849), .b(x_in_43_6), .c(n_2850), .d(n_5327), .o(n_7746) );
oa22f80 g563214 ( .a(n_5297), .b(n_5296), .c(n_5295), .d(x_in_5_5), .o(n_6809) );
ao22s80 g563215 ( .a(n_2988), .b(x_in_5_6), .c(n_5294), .d(n_3568), .o(n_6953) );
in01f80 g563216 ( .a(n_7011), .o(n_9312) );
oa22f80 g563217 ( .a(n_2726), .b(x_in_43_4), .c(n_2727), .d(n_5293), .o(n_7011) );
ao12f80 g563218 ( .a(n_3590), .b(n_5036), .c(x_in_5_7), .o(n_6927) );
oa22f80 g563219 ( .a(n_5292), .b(n_5291), .c(n_2966), .d(x_in_5_8), .o(n_6876) );
in01f80 g563220 ( .a(n_6997), .o(n_9303) );
oa12f80 g563221 ( .a(n_3921), .b(n_3920), .c(x_in_43_3), .o(n_6997) );
in01f80 g563222 ( .a(n_9591), .o(n_9001) );
oa12f80 g563223 ( .a(n_3503), .b(n_3502), .c(x_in_43_2), .o(n_9591) );
ao22s80 g563224 ( .a(n_2980), .b(x_in_5_11), .c(n_5290), .d(n_5754), .o(n_6806) );
oa22f80 g563225 ( .a(n_5811), .b(n_6458), .c(n_6457), .d(n_5810), .o(n_9352) );
ao22s80 g563226 ( .a(n_2955), .b(x_in_5_12), .c(n_5289), .d(n_5888), .o(n_6803) );
ao22s80 g563227 ( .a(n_2981), .b(x_in_5_13), .c(n_5288), .d(n_13241), .o(n_6924) );
ao22s80 g563228 ( .a(n_3396), .b(x_in_5_11), .c(n_5755), .d(n_5754), .o(n_7614) );
in01f80 g563229 ( .a(n_8531), .o(n_6544) );
ao22s80 g563230 ( .a(n_3765), .b(n_5888), .c(n_3766), .d(x_in_5_12), .o(n_8531) );
oa22f80 g563231 ( .a(n_4977), .b(n_5730), .c(n_8569), .d(n_4976), .o(n_7611) );
oa12f80 g563232 ( .a(n_5122), .b(n_5121), .c(n_5790), .o(n_8317) );
in01f80 g563233 ( .a(n_7024), .o(n_9229) );
oa22f80 g563234 ( .a(n_2970), .b(x_in_43_14), .c(n_2971), .d(n_7311), .o(n_7024) );
in01f80 g563235 ( .a(n_12160), .o(n_6543) );
ao12f80 g563236 ( .a(n_4368), .b(n_5409), .c(x_in_37_7), .o(n_12160) );
in01f80 g563237 ( .a(n_13001), .o(n_6542) );
oa22f80 g563238 ( .a(n_5887), .b(x_in_21_4), .c(n_5861), .d(n_8557), .o(n_13001) );
in01f80 g563239 ( .a(n_9227), .o(n_8442) );
ao12f80 g563240 ( .a(n_3623), .b(n_3622), .c(x_in_37_8), .o(n_9227) );
ao12f80 g563241 ( .a(n_5117), .b(n_5116), .c(n_5115), .o(n_8325) );
in01f80 g563242 ( .a(FE_OFN783_n_10771), .o(n_12602) );
oa22f80 g563243 ( .a(n_5886), .b(x_in_37_8), .c(n_5885), .d(n_5881), .o(n_10771) );
in01f80 g563244 ( .a(FE_OFN779_n_12158), .o(n_6541) );
oa22f80 g563245 ( .a(n_5883), .b(x_in_37_6), .c(n_5882), .d(n_5884), .o(n_12158) );
ao12f80 g563246 ( .a(n_4617), .b(n_5873), .c(n_4616), .o(n_7771) );
oa22f80 g563247 ( .a(n_5883), .b(x_in_37_10), .c(n_5882), .d(n_5745), .o(n_8858) );
in01f80 g563248 ( .a(n_8492), .o(n_5738) );
ao22s80 g563249 ( .a(n_5287), .b(n_2130), .c(n_5286), .d(n_2131), .o(n_8492) );
in01f80 g563250 ( .a(n_12154), .o(n_6540) );
oa12f80 g563251 ( .a(n_4676), .b(n_5880), .c(x_in_37_4), .o(n_12154) );
ao22s80 g563252 ( .a(n_4053), .b(n_5881), .c(n_5880), .d(x_in_37_8), .o(n_9053) );
in01f80 g563253 ( .a(n_12978), .o(n_6460) );
ao22s80 g563254 ( .a(n_5411), .b(n_4654), .c(n_5062), .d(x_in_37_3), .o(n_12978) );
in01f80 g563255 ( .a(n_13029), .o(n_12979) );
oa12f80 g563256 ( .a(n_4378), .b(n_5740), .c(x_in_37_2), .o(n_13029) );
oa12f80 g563257 ( .a(n_5878), .b(n_4862), .c(n_5871), .o(n_5879) );
ao22s80 g563258 ( .a(n_5877), .b(n_3780), .c(n_5876), .d(n_3729), .o(n_7827) );
in01f80 g563259 ( .a(n_9225), .o(n_5875) );
oa12f80 g563260 ( .a(n_3933), .b(n_3932), .c(x_in_37_15), .o(n_9225) );
oa22f80 g563261 ( .a(n_5874), .b(x_in_3_6), .c(n_3588), .d(n_5515), .o(n_7381) );
in01f80 g563262 ( .a(n_8533), .o(n_6539) );
oa22f80 g563263 ( .a(n_3678), .b(x_in_57_12), .c(n_3679), .d(n_5302), .o(n_8533) );
in01f80 g563264 ( .a(n_6974), .o(n_9222) );
oa22f80 g563265 ( .a(n_2787), .b(x_in_27_8), .c(n_2788), .d(n_7287), .o(n_6974) );
oa22f80 g563266 ( .a(n_5873), .b(x_in_21_11), .c(n_5087), .d(n_5872), .o(n_7684) );
in01f80 g563267 ( .a(n_7015), .o(n_9261) );
oa22f80 g563268 ( .a(n_2890), .b(x_in_27_9), .c(n_2891), .d(n_7289), .o(n_7015) );
oa12f80 g563269 ( .a(n_5147), .b(n_5146), .c(FE_OFN612_n_5698), .o(n_6538) );
in01f80 g563270 ( .a(n_6991), .o(n_9220) );
oa22f80 g563271 ( .a(n_3343), .b(x_in_27_6), .c(n_3344), .d(n_5677), .o(n_6991) );
oa12f80 g563272 ( .a(n_4229), .b(n_4706), .c(n_4228), .o(n_8954) );
in01f80 g563273 ( .a(n_9218), .o(n_8328) );
oa12f80 g563274 ( .a(n_3898), .b(n_3897), .c(x_in_27_5), .o(n_9218) );
oa22f80 g563275 ( .a(n_5751), .b(x_in_21_11), .c(n_3595), .d(n_5872), .o(n_8011) );
oa12f80 g563276 ( .a(n_5112), .b(n_5111), .c(n_5789), .o(n_8302) );
oa12f80 g563277 ( .a(n_3555), .b(n_3554), .c(x_in_11_1), .o(n_8639) );
in01f80 g563278 ( .a(n_6999), .o(n_8536) );
ao12f80 g563279 ( .a(n_3517), .b(n_4015), .c(n_3516), .o(n_6999) );
ao22s80 g563280 ( .a(n_3606), .b(x_in_37_2), .c(n_5871), .d(n_3011), .o(n_8570) );
ao22s80 g563281 ( .a(n_5870), .b(n_5869), .c(n_5903), .d(x_in_21_10), .o(n_7651) );
ao22s80 g563282 ( .a(n_5762), .b(n_5868), .c(n_5867), .d(n_5866), .o(n_7603) );
oa22f80 g563283 ( .a(n_2974), .b(x_in_25_10), .c(n_4909), .d(n_2743), .o(n_7068) );
oa22f80 g563284 ( .a(n_2915), .b(x_in_25_11), .c(n_5285), .d(n_3189), .o(n_7065) );
oa22f80 g563285 ( .a(n_5864), .b(n_5863), .c(n_5862), .d(n_3758), .o(n_7959) );
oa22f80 g563286 ( .a(n_5887), .b(x_in_21_8), .c(n_5861), .d(n_5860), .o(n_7688) );
ao22s80 g563287 ( .a(n_2937), .b(n_5293), .c(n_5284), .d(x_in_43_4), .o(n_7052) );
in01f80 g563288 ( .a(n_7036), .o(n_9224) );
oa22f80 g563289 ( .a(n_2968), .b(x_in_27_14), .c(n_2969), .d(n_14997), .o(n_7036) );
in01f80 g563290 ( .a(n_8444), .o(n_7786) );
oa22f80 g563291 ( .a(n_5273), .b(n_7263), .c(n_5274), .d(x_in_43_12), .o(n_8444) );
oa22f80 g563292 ( .a(n_4899), .b(n_5283), .c(FE_OFN931_n_4898), .d(x_in_51_10), .o(n_8470) );
in01f80 g563293 ( .a(n_12640), .o(n_9050) );
oa12f80 g563294 ( .a(n_3895), .b(n_3894), .c(x_in_61_9), .o(n_12640) );
oa22f80 g563295 ( .a(n_3993), .b(x_in_33_4), .c(n_5282), .d(n_5281), .o(n_10705) );
oa22f80 g563296 ( .a(n_2952), .b(n_6746), .c(n_5280), .d(x_in_3_13), .o(n_6798) );
oa12f80 g563297 ( .a(n_4227), .b(n_4236), .c(n_4226), .o(n_8943) );
ao12f80 g563298 ( .a(n_4150), .b(n_4149), .c(n_4148), .o(n_8558) );
ao22s80 g563299 ( .a(n_5279), .b(n_3500), .c(n_5278), .d(n_3788), .o(n_26266) );
ao22s80 g563300 ( .a(n_4230), .b(x_in_21_3), .c(n_4108), .d(n_6781), .o(n_7888) );
oa12f80 g563301 ( .a(n_3423), .b(n_5277), .c(x_in_25_4), .o(n_7142) );
ao22s80 g563302 ( .a(n_2957), .b(x_in_57_13), .c(n_5276), .d(n_3560), .o(n_6913) );
in01f80 g563303 ( .a(n_9676), .o(n_7660) );
oa12f80 g563304 ( .a(n_3815), .b(n_3814), .c(x_in_59_9), .o(n_9676) );
ao22s80 g563305 ( .a(n_5859), .b(n_3753), .c(n_5858), .d(n_3841), .o(n_7831) );
in01f80 g563306 ( .a(n_6536), .o(n_6537) );
oa12f80 g563307 ( .a(n_4691), .b(n_5229), .c(n_5231), .o(n_6536) );
ao22s80 g563308 ( .a(n_3165), .b(n_5275), .c(n_3164), .d(x_in_59_6), .o(n_9582) );
in01f80 g563309 ( .a(n_7127), .o(n_9214) );
oa22f80 g563310 ( .a(n_2907), .b(x_in_59_4), .c(n_2908), .d(n_5271), .o(n_7127) );
in01f80 g563311 ( .a(n_7000), .o(n_9282) );
oa12f80 g563312 ( .a(n_3419), .b(n_3418), .c(x_in_59_3), .o(n_7000) );
ao22s80 g563313 ( .a(n_5274), .b(n_3437), .c(n_5273), .d(n_3650), .o(n_26270) );
in01f80 g563314 ( .a(n_8521), .o(n_7779) );
oa22f80 g563315 ( .a(n_2802), .b(n_5272), .c(n_2803), .d(x_in_7_3), .o(n_8521) );
in01f80 g563316 ( .a(n_12586), .o(n_8980) );
oa12f80 g563317 ( .a(n_3627), .b(n_3626), .c(x_in_61_8), .o(n_12586) );
ao22s80 g563318 ( .a(n_2861), .b(n_5271), .c(n_5270), .d(x_in_59_4), .o(n_7077) );
ao12f80 g563319 ( .a(n_3883), .b(n_5269), .c(n_5268), .o(n_10083) );
in01f80 g563320 ( .a(n_5857), .o(n_7948) );
oa12f80 g563321 ( .a(n_3579), .b(n_3916), .c(n_5267), .o(n_5857) );
ao12f80 g563322 ( .a(n_4641), .b(n_4640), .c(n_4639), .o(n_8768) );
oa22f80 g563323 ( .a(n_5248), .b(FE_OFN256_n_4280), .c(n_1570), .d(FE_OFN1108_rst), .o(n_6535) );
oa22f80 g563324 ( .a(n_7385), .b(n_29046), .c(n_230), .d(FE_OFN1172_n_4860), .o(n_7386) );
in01f80 g563325 ( .a(n_8609), .o(n_6534) );
ao22s80 g563326 ( .a(n_3598), .b(n_5856), .c(n_5855), .d(n_5772), .o(n_8609) );
ao22s80 g563327 ( .a(n_6532), .b(n_4312), .c(x_out_57_21), .d(FE_OFN274_n_16893), .o(n_6533) );
ao22s80 g563328 ( .a(n_4921), .b(n_2800), .c(x_out_63_21), .d(FE_OFN271_n_16028), .o(n_4922) );
ao22s80 g563329 ( .a(n_6530), .b(n_4234), .c(x_out_58_21), .d(FE_OFN280_n_16656), .o(n_6531) );
ao22s80 g563330 ( .a(n_6528), .b(n_4222), .c(x_out_60_21), .d(FE_OFN271_n_16028), .o(n_6529) );
ao22s80 g563331 ( .a(n_6526), .b(n_4306), .c(x_out_61_21), .d(FE_OFN273_n_16893), .o(n_6527) );
ao22s80 g563332 ( .a(n_6524), .b(n_4294), .c(x_out_59_21), .d(n_16028), .o(n_6525) );
ao22s80 g563333 ( .a(n_6522), .b(n_4142), .c(x_out_62_21), .d(FE_OFN1162_n_5003), .o(n_6523) );
ao22s80 g563334 ( .a(n_10224), .b(n_4657), .c(n_10226), .d(n_6984), .o(n_9718) );
oa22f80 g563335 ( .a(n_5854), .b(n_5251), .c(n_5822), .d(n_5253), .o(n_7942) );
in01f80 g563336 ( .a(n_8118), .o(n_5266) );
oa22f80 g563337 ( .a(n_5329), .b(n_6350), .c(x_in_51_5), .d(x_in_51_3), .o(n_8118) );
ao22s80 g563338 ( .a(n_7211), .b(n_6478), .c(n_6477), .d(n_4970), .o(n_8337) );
ao22s80 g563339 ( .a(n_12366), .b(n_4929), .c(FE_OFN554_n_9468), .d(n_4928), .o(n_15651) );
ao22s80 g563340 ( .a(n_9034), .b(n_4476), .c(FE_OFN544_n_9030), .d(n_5265), .o(n_7114) );
oa22f80 g563341 ( .a(FE_OFN548_n_10452), .b(n_6372), .c(n_9638), .d(n_4481), .o(n_10325) );
ao22s80 g563342 ( .a(n_11700), .b(n_5264), .c(n_9480), .d(n_5263), .o(n_12860) );
ao22s80 g563343 ( .a(n_9042), .b(n_6032), .c(FE_OFN546_n_9036), .d(n_4170), .o(n_8807) );
oa22f80 g563344 ( .a(n_3529), .b(n_2645), .c(n_3113), .d(x_in_5_7), .o(n_7186) );
in01f80 g563345 ( .a(n_8345), .o(n_7384) );
oa22f80 g563346 ( .a(n_6521), .b(x_in_35_4), .c(n_4396), .d(n_5987), .o(n_8345) );
ao22s80 g563347 ( .a(n_3611), .b(x_in_17_4), .c(n_5853), .d(n_4021), .o(n_7729) );
oa22f80 g563348 ( .a(n_5852), .b(n_3024), .c(n_5851), .d(n_7653), .o(n_7794) );
ao22s80 g563349 ( .a(n_3612), .b(x_in_3_4), .c(n_5850), .d(n_5931), .o(n_7816) );
ao22s80 g563350 ( .a(n_3109), .b(x_in_43_7), .c(n_3404), .d(n_5519), .o(n_5262) );
oa22f80 g563351 ( .a(n_5261), .b(x_in_19_1), .c(n_5260), .d(n_3763), .o(n_8658) );
in01f80 g563352 ( .a(n_8084), .o(n_5259) );
oa22f80 g563353 ( .a(FE_OFN1246_n_4900), .b(n_6351), .c(x_in_51_7), .d(x_in_51_5), .o(n_8084) );
ao22s80 g563354 ( .a(n_3441), .b(x_in_59_3), .c(n_4288), .d(n_3260), .o(n_7920) );
ao22s80 g563355 ( .a(n_2885), .b(x_in_27_6), .c(n_3383), .d(n_5677), .o(n_5258) );
ao22s80 g563356 ( .a(n_3134), .b(x_in_7_5), .c(n_3996), .d(n_5256), .o(n_5257) );
ao22s80 g563357 ( .a(n_3439), .b(x_in_37_12), .c(n_3440), .d(n_5849), .o(n_7951) );
in01f80 g563358 ( .a(FE_OFN761_n_9661), .o(n_7752) );
oa22f80 g563359 ( .a(n_7086), .b(x_in_35_14), .c(n_3068), .d(n_2752), .o(n_9661) );
oa22f80 g563360 ( .a(n_5864), .b(n_5848), .c(n_5862), .d(x_in_9_1), .o(n_7965) );
in01f80 g563361 ( .a(n_8911), .o(n_6520) );
oa22f80 g563362 ( .a(n_6760), .b(n_10829), .c(n_7884), .d(x_in_41_12), .o(n_8911) );
in01f80 g563363 ( .a(n_9428), .o(n_7383) );
na02f80 g563364 ( .a(n_5168), .b(n_4342), .o(n_9428) );
in01f80 g563365 ( .a(n_6795), .o(n_9266) );
oa22f80 g563366 ( .a(n_5345), .b(x_in_19_2), .c(n_5347), .d(n_2440), .o(n_6795) );
ao22s80 g563367 ( .a(n_12197), .b(n_4042), .c(n_5558), .d(n_2672), .o(n_5255) );
ao22s80 g563368 ( .a(n_5253), .b(n_5252), .c(n_5251), .d(x_in_19_3), .o(n_7058) );
in01f80 g563369 ( .a(n_8906), .o(n_8904) );
oa22f80 g563370 ( .a(n_6285), .b(n_3077), .c(n_2843), .d(x_in_13_14), .o(n_8906) );
in01f80 g563371 ( .a(n_7457), .o(n_7619) );
ao22s80 g563372 ( .a(n_4892), .b(x_in_41_3), .c(n_5250), .d(n_2424), .o(n_7457) );
in01f80 g563373 ( .a(FE_OFN480_n_12184), .o(n_6519) );
ao22s80 g563374 ( .a(n_8092), .b(x_in_7_8), .c(n_5847), .d(n_7304), .o(n_12184) );
in01f80 g563375 ( .a(n_5845), .o(n_5846) );
oa22f80 g563376 ( .a(FE_OFN612_n_5698), .b(x_in_19_13), .c(n_5243), .d(n_5556), .o(n_5845) );
ao22s80 g563377 ( .a(n_4916), .b(x_in_49_5), .c(n_4562), .d(n_5095), .o(n_7022) );
ao22s80 g563378 ( .a(n_5844), .b(n_6750), .c(n_6751), .d(n_5443), .o(n_7962) );
in01f80 g563379 ( .a(FE_OFN1186_n_12201), .o(n_5843) );
oa22f80 g563380 ( .a(FE_OFN1188_n_5249), .b(n_5256), .c(n_5248), .d(x_in_7_5), .o(n_12201) );
in01f80 g563381 ( .a(FE_OFN456_n_8508), .o(n_5842) );
oa22f80 g563382 ( .a(FE_OFN458_n_5621), .b(n_5247), .c(n_4908), .d(x_in_3_12), .o(n_8508) );
in01f80 g563383 ( .a(FE_OFN963_n_9280), .o(n_5841) );
oa22f80 g563384 ( .a(n_5246), .b(n_2654), .c(n_6856), .d(x_in_53_8), .o(n_9280) );
in01f80 g563385 ( .a(FE_OFN1083_n_8877), .o(n_6518) );
ao22s80 g563386 ( .a(n_8089), .b(x_in_61_5), .c(n_5840), .d(n_5242), .o(n_8877) );
in01f80 g563387 ( .a(n_9270), .o(n_7875) );
oa22f80 g563388 ( .a(n_4915), .b(n_2655), .c(FE_OFN1091_n_8621), .d(x_in_61_15), .o(n_9270) );
ao22s80 g563389 ( .a(n_8971), .b(x_in_61_7), .c(n_4924), .d(n_5839), .o(n_8601) );
ao22s80 g563390 ( .a(n_4767), .b(n_5825), .c(n_3989), .d(x_in_3_3), .o(n_7133) );
in01f80 g563391 ( .a(n_8026), .o(n_8525) );
oa22f80 g563392 ( .a(FE_OFN765_n_5707), .b(n_5032), .c(n_5031), .d(x_in_35_12), .o(n_8026) );
oa22f80 g563393 ( .a(FE_OFN765_n_5707), .b(x_in_35_13), .c(n_5031), .d(n_5245), .o(n_8501) );
in01f80 g563394 ( .a(n_12684), .o(n_12690) );
oa22f80 g563395 ( .a(n_3392), .b(n_8165), .c(n_8157), .d(x_in_7_10), .o(n_12684) );
oa22f80 g563396 ( .a(n_6751), .b(n_5838), .c(n_5844), .d(n_8539), .o(n_7944) );
ao22s80 g563397 ( .a(n_4341), .b(n_5900), .c(n_5837), .d(x_in_21_5), .o(n_7673) );
in01f80 g563398 ( .a(n_8907), .o(n_8909) );
oa22f80 g563399 ( .a(FE_OFN612_n_5698), .b(n_5244), .c(n_5243), .d(x_in_19_12), .o(n_8907) );
in01f80 g563400 ( .a(FE_OFN967_n_9286), .o(n_5836) );
oa22f80 g563401 ( .a(n_4902), .b(n_2653), .c(FE_OFN973_n_6822), .d(x_in_53_10), .o(n_9286) );
in01f80 g563402 ( .a(n_8515), .o(n_7872) );
oa22f80 g563403 ( .a(n_4938), .b(n_4937), .c(FE_OFN1087_n_8974), .d(x_in_61_8), .o(n_8515) );
in01f80 g563404 ( .a(n_8468), .o(n_7867) );
oa22f80 g563405 ( .a(n_4652), .b(n_3833), .c(FE_OFN1274_n_8977), .d(x_in_61_10), .o(n_8468) );
in01f80 g563406 ( .a(n_11557), .o(n_6517) );
ao22s80 g563407 ( .a(n_5851), .b(x_in_9_2), .c(n_5852), .d(n_5216), .o(n_11557) );
ao22s80 g563408 ( .a(n_7581), .b(n_5723), .c(n_8477), .d(n_5835), .o(n_7974) );
in01f80 g563409 ( .a(n_6933), .o(n_5834) );
oa22f80 g563410 ( .a(FE_OFN458_n_5621), .b(x_in_3_13), .c(n_4908), .d(n_6746), .o(n_6933) );
in01f80 g563411 ( .a(n_12163), .o(n_5833) );
oa22f80 g563412 ( .a(n_6399), .b(n_5242), .c(FE_OFN1129_n_6399), .d(x_in_61_5), .o(n_12163) );
ao22s80 g563413 ( .a(n_3427), .b(x_in_35_4), .c(n_5832), .d(n_5987), .o(n_7856) );
oa22f80 g563414 ( .a(n_5241), .b(x_in_33_13), .c(FE_OFN726_n_5240), .d(n_2533), .o(n_7189) );
oa22f80 g563415 ( .a(n_5831), .b(x_in_57_11), .c(n_4739), .d(n_5313), .o(n_7703) );
oa22f80 g563416 ( .a(n_5239), .b(x_in_53_15), .c(FE_OFN971_n_6854), .d(n_3193), .o(n_8147) );
in01f80 g563417 ( .a(n_6515), .o(n_6516) );
ao22s80 g563418 ( .a(n_5826), .b(n_4419), .c(n_5830), .d(x_in_3_1), .o(n_6515) );
in01f80 g563419 ( .a(n_7740), .o(n_9285) );
oa22f80 g563420 ( .a(n_5828), .b(n_3608), .c(n_8142), .d(x_in_61_3), .o(n_7740) );
in01f80 g563421 ( .a(FE_OFN965_n_9283), .o(n_5829) );
oa22f80 g563422 ( .a(n_5239), .b(n_2550), .c(FE_OFN971_n_6854), .d(x_in_53_9), .o(n_9283) );
in01f80 g563423 ( .a(n_8565), .o(n_6514) );
oa22f80 g563424 ( .a(n_5743), .b(x_in_51_4), .c(n_5821), .d(n_5979), .o(n_8565) );
in01f80 g563425 ( .a(n_8111), .o(n_9242) );
oa22f80 g563426 ( .a(n_8295), .b(x_in_37_1), .c(n_8297), .d(n_4376), .o(n_8111) );
in01f80 g563427 ( .a(n_8074), .o(n_8523) );
oa22f80 g563428 ( .a(n_4915), .b(n_4914), .c(FE_OFN1091_n_8621), .d(x_in_61_9), .o(n_8074) );
in01f80 g563429 ( .a(n_12968), .o(n_6513) );
ao22s80 g563430 ( .a(n_8142), .b(x_in_61_8), .c(n_5828), .d(n_4937), .o(n_12968) );
in01f80 g563431 ( .a(n_12983), .o(n_12579) );
oa22f80 g563432 ( .a(n_8086), .b(n_4914), .c(n_5771), .d(x_in_61_9), .o(n_12983) );
ao22s80 g563433 ( .a(n_10216), .b(x_in_53_3), .c(n_10218), .d(n_5827), .o(n_8139) );
ao22s80 g563434 ( .a(n_5826), .b(n_5825), .c(n_5830), .d(x_in_3_3), .o(n_7663) );
in01f80 g563435 ( .a(n_8926), .o(n_8356) );
oa22f80 g563436 ( .a(n_8086), .b(n_8929), .c(n_5771), .d(x_in_61_4), .o(n_8926) );
oa22f80 g563437 ( .a(n_10222), .b(n_2525), .c(n_10220), .d(x_in_53_7), .o(n_8603) );
ao22s80 g563438 ( .a(n_11148), .b(x_in_53_4), .c(n_8503), .d(n_3038), .o(n_8599) );
ao22s80 g563439 ( .a(n_11168), .b(x_in_53_6), .c(n_8502), .d(n_2651), .o(n_8602) );
ao22s80 g563440 ( .a(n_8297), .b(n_5742), .c(n_8295), .d(x_in_37_5), .o(n_7606) );
ao22s80 g563441 ( .a(n_6760), .b(n_9608), .c(n_9604), .d(x_in_41_12), .o(n_7885) );
in01f80 g563442 ( .a(n_7091), .o(n_8878) );
oa22f80 g563443 ( .a(n_5241), .b(x_in_33_12), .c(FE_OFN726_n_5240), .d(n_12635), .o(n_7091) );
oa22f80 g563444 ( .a(n_8485), .b(n_2626), .c(n_11166), .d(x_in_53_5), .o(n_8605) );
oa22f80 g563445 ( .a(n_6751), .b(x_in_33_6), .c(n_5844), .d(n_12172), .o(n_8573) );
ao22s80 g563446 ( .a(n_10214), .b(x_in_53_3), .c(n_10212), .d(n_5827), .o(n_8594) );
ao22s80 g563447 ( .a(n_5824), .b(x_in_61_11), .c(n_9088), .d(n_4529), .o(n_8600) );
oa22f80 g563448 ( .a(n_5823), .b(x_in_9_12), .c(n_8704), .d(n_8957), .o(n_7735) );
oa22f80 g563449 ( .a(n_8477), .b(n_3186), .c(n_7581), .d(x_in_49_11), .o(n_7630) );
in01f80 g563450 ( .a(n_5235), .o(n_5236) );
oa22f80 g563451 ( .a(n_4793), .b(n_3173), .c(n_3370), .d(n_12178), .o(n_5235) );
ao22s80 g563452 ( .a(n_5854), .b(x_in_19_4), .c(n_5822), .d(n_5939), .o(n_7755) );
ao22s80 g563453 ( .a(n_5821), .b(x_in_51_3), .c(n_5743), .d(n_5180), .o(n_7908) );
ao22s80 g563454 ( .a(n_5980), .b(x_in_51_4), .c(n_10817), .d(n_5979), .o(n_7758) );
in01f80 g563455 ( .a(n_5233), .o(n_5234) );
oa22f80 g563456 ( .a(FE_OFN726_n_5240), .b(n_6904), .c(n_2538), .d(x_in_33_14), .o(n_5233) );
ao22s80 g563457 ( .a(n_4098), .b(x_in_33_6), .c(n_5230), .d(n_5820), .o(n_10773) );
oa22f80 g563458 ( .a(n_5232), .b(n_8885), .c(n_5231), .d(n_5230), .o(n_10798) );
in01f80 g563459 ( .a(n_5818), .o(n_5819) );
oa22f80 g563460 ( .a(n_5229), .b(n_12175), .c(n_5228), .d(n_3073), .o(n_5818) );
in01f80 g563461 ( .a(n_5816), .o(n_5817) );
oa22f80 g563462 ( .a(n_5227), .b(n_12634), .c(n_5226), .d(n_3311), .o(n_5816) );
oa22f80 g563463 ( .a(n_5225), .b(n_8884), .c(n_5224), .d(n_3106), .o(n_10785) );
oa22f80 g563464 ( .a(n_5223), .b(n_11297), .c(n_5820), .d(n_3015), .o(n_10775) );
no02f80 g563638 ( .a(n_4020), .b(n_7195), .o(n_7958) );
in01f80 g563639 ( .a(n_13251), .o(n_6660) );
na02f80 g563640 ( .a(n_8376), .b(x_in_38_0), .o(n_13251) );
na02f80 g563641 ( .a(n_3628), .b(n_1439), .o(n_5222) );
na02f80 g563642 ( .a(n_4790), .b(x_in_23_4), .o(n_10107) );
no02f80 g563643 ( .a(n_6577), .b(n_5221), .o(n_8406) );
na02f80 g563644 ( .a(n_4288), .b(x_in_59_3), .o(n_10091) );
na02f80 g563645 ( .a(n_4789), .b(x_in_47_4), .o(n_10101) );
na02f80 g563646 ( .a(n_4788), .b(x_in_55_4), .o(n_10103) );
na02f80 g563647 ( .a(n_4787), .b(x_in_31_4), .o(n_9385) );
na02f80 g563648 ( .a(n_4786), .b(x_in_63_4), .o(n_10097) );
na02f80 g563649 ( .a(n_2116), .b(n_2851), .o(n_7193) );
no02f80 g563650 ( .a(n_3646), .b(x_in_13_3), .o(n_4861) );
na02f80 g563651 ( .a(n_4016), .b(x_in_49_0), .o(n_4019) );
no02f80 g563652 ( .a(n_4018), .b(n_4017), .o(n_8397) );
no02f80 g563653 ( .a(n_4016), .b(x_in_49_0), .o(n_10983) );
na02f80 g563654 ( .a(n_3607), .b(x_in_28_0), .o(n_13246) );
na02f80 g563655 ( .a(n_7813), .b(n_1449), .o(n_5220) );
na02f80 g563656 ( .a(n_4785), .b(x_in_15_4), .o(n_10105) );
na02f80 g563657 ( .a(n_4783), .b(n_4782), .o(n_4784) );
na02f80 g563658 ( .a(n_4780), .b(n_4779), .o(n_4781) );
no02f80 g563659 ( .a(n_4828), .b(x_in_29_0), .o(n_11609) );
na03f80 g563660 ( .a(n_7099), .b(n_2185), .c(FE_OFN419_n_16909), .o(n_6070) );
na02f80 g563661 ( .a(n_4394), .b(n_4393), .o(n_4395) );
na02f80 g563662 ( .a(n_4777), .b(n_3162), .o(n_4778) );
na03f80 g563663 ( .a(n_7102), .b(n_2236), .c(FE_OFN384_n_16289), .o(n_7221) );
na02f80 g563664 ( .a(n_4775), .b(n_4774), .o(n_4776) );
no02f80 g563665 ( .a(n_4015), .b(n_6788), .o(n_12117) );
no02f80 g563666 ( .a(n_4916), .b(n_4013), .o(n_4014) );
no02f80 g563667 ( .a(n_6571), .b(n_5219), .o(n_8410) );
no02f80 g563668 ( .a(n_3253), .b(x_in_1_3), .o(n_5694) );
no02f80 g563669 ( .a(n_4772), .b(x_in_17_0), .o(n_4773) );
na02f80 g563670 ( .a(n_5215), .b(n_4011), .o(n_4012) );
no02f80 g563671 ( .a(n_5218), .b(n_5217), .o(n_8412) );
no02f80 g563672 ( .a(n_6563), .b(n_5023), .o(n_8416) );
no02f80 g563673 ( .a(n_5851), .b(n_5216), .o(n_8400) );
no02f80 g563674 ( .a(n_4771), .b(n_2331), .o(n_9191) );
no02f80 g563675 ( .a(n_4052), .b(n_5215), .o(n_10079) );
no02f80 g563676 ( .a(n_5891), .b(n_5213), .o(n_5214) );
na02f80 g563677 ( .a(n_2102), .b(n_7057), .o(n_7941) );
no02f80 g563678 ( .a(n_5197), .b(x_in_39_5), .o(n_6673) );
no02f80 g563679 ( .a(n_5212), .b(n_5211), .o(n_8408) );
in01f80 g563680 ( .a(n_6379), .o(n_4010) );
na02f80 g563681 ( .a(n_2081), .b(n_3530), .o(n_6379) );
in01f80 g563682 ( .a(n_6388), .o(n_4009) );
na02f80 g563683 ( .a(n_2294), .b(n_3399), .o(n_6388) );
in01f80 g563684 ( .a(n_4858), .o(n_6377) );
na02f80 g563685 ( .a(n_2137), .b(n_3535), .o(n_4858) );
no02f80 g563686 ( .a(n_5210), .b(n_5209), .o(n_8414) );
no02f80 g563687 ( .a(n_5814), .b(n_5813), .o(n_5815) );
in01f80 g563688 ( .a(n_4006), .o(n_8484) );
ao12f80 g563689 ( .a(n_4757), .b(n_1988), .c(x_in_19_14), .o(n_4006) );
in01f80 g563690 ( .a(n_4854), .o(n_6365) );
na02f80 g563691 ( .a(n_2292), .b(n_3968), .o(n_4854) );
na02f80 g563692 ( .a(n_6296), .b(x_in_13_3), .o(n_10073) );
in01f80 g563693 ( .a(n_6375), .o(n_3769) );
na02f80 g563694 ( .a(n_2203), .b(n_3545), .o(n_6375) );
na02f80 g563695 ( .a(n_5701), .b(n_4004), .o(n_4005) );
in01f80 g563696 ( .a(n_4769), .o(n_4770) );
no02f80 g563697 ( .a(n_4003), .b(n_2436), .o(n_4769) );
in01f80 g563698 ( .a(n_6368), .o(n_4002) );
na02f80 g563699 ( .a(n_2069), .b(n_3963), .o(n_6368) );
in01f80 g563700 ( .a(n_8459), .o(n_5208) );
no02f80 g563701 ( .a(n_2934), .b(n_4768), .o(n_8459) );
na02f80 g563702 ( .a(n_5322), .b(n_4768), .o(n_4137) );
no02f80 g563703 ( .a(n_7639), .b(n_4766), .o(n_10956) );
in01f80 g563704 ( .a(n_13282), .o(n_5006) );
no02f80 g563705 ( .a(n_4767), .b(n_4766), .o(n_13282) );
no02f80 g563706 ( .a(n_4251), .b(n_4250), .o(n_4252) );
in01f80 g563707 ( .a(n_6384), .o(n_4001) );
na02f80 g563708 ( .a(n_2079), .b(n_3954), .o(n_6384) );
no02f80 g563709 ( .a(n_4765), .b(n_4828), .o(n_14491) );
no02f80 g563710 ( .a(n_5701), .b(n_5700), .o(n_3478) );
no02f80 g563711 ( .a(n_7895), .b(x_in_13_12), .o(n_4764) );
na02f80 g563712 ( .a(n_7895), .b(x_in_13_12), .o(n_10948) );
no02f80 g563713 ( .a(n_6576), .b(n_5207), .o(n_7129) );
na02f80 g563714 ( .a(n_5205), .b(n_5204), .o(n_5206) );
no02f80 g563715 ( .a(n_6577), .b(n_5034), .o(n_5035) );
na02f80 g563716 ( .a(n_3355), .b(n_3354), .o(n_3356) );
no02f80 g563717 ( .a(n_7598), .b(n_4000), .o(n_8774) );
na02f80 g563718 ( .a(n_4891), .b(x_in_45_4), .o(n_10059) );
in01f80 g563719 ( .a(n_6082), .o(n_7218) );
no02f80 g563720 ( .a(n_4892), .b(n_4832), .o(n_6082) );
no02f80 g563721 ( .a(n_5811), .b(n_5810), .o(n_5812) );
no02f80 g563722 ( .a(n_5808), .b(n_5807), .o(n_5809) );
na02f80 g563723 ( .a(n_2790), .b(n_4763), .o(n_11615) );
no02f80 g563724 ( .a(n_9984), .b(n_7086), .o(n_4762) );
na02f80 g563725 ( .a(n_9984), .b(n_7086), .o(n_4761) );
na02f80 g563726 ( .a(n_4760), .b(n_4144), .o(n_6652) );
in01f80 g563727 ( .a(n_4989), .o(n_4990) );
no02f80 g563728 ( .a(n_4760), .b(n_4144), .o(n_4989) );
na02f80 g563729 ( .a(n_4895), .b(n_4894), .o(n_9422) );
na02f80 g563730 ( .a(n_5923), .b(x_in_53_12), .o(n_5203) );
na02f80 g563731 ( .a(n_3998), .b(n_4759), .o(n_3999) );
in01f80 g563732 ( .a(n_12091), .o(n_5202) );
no02f80 g563733 ( .a(n_3205), .b(n_4759), .o(n_12091) );
na02f80 g563734 ( .a(n_7847), .b(x_in_7_1), .o(n_4322) );
na02f80 g563735 ( .a(n_5928), .b(n_4757), .o(n_4758) );
in01f80 g563736 ( .a(n_6361), .o(n_3997) );
na02f80 g563737 ( .a(n_2202), .b(n_4138), .o(n_6361) );
no02f80 g563738 ( .a(n_3996), .b(x_in_7_5), .o(n_5702) );
na02f80 g563739 ( .a(n_3601), .b(n_5034), .o(n_7917) );
na02f80 g563740 ( .a(n_5200), .b(n_5199), .o(n_5201) );
na02f80 g563741 ( .a(n_5197), .b(n_4338), .o(n_5198) );
na02f80 g563742 ( .a(n_2754), .b(n_4755), .o(n_4756) );
no02f80 g563743 ( .a(n_5893), .b(n_4325), .o(n_4326) );
na02f80 g563744 ( .a(n_3382), .b(n_5195), .o(n_5196) );
no02f80 g563745 ( .a(n_6477), .b(n_5805), .o(n_5806) );
in01f80 g563746 ( .a(n_3995), .o(n_5692) );
oa12f80 g563747 ( .a(n_2878), .b(n_2016), .c(x_in_59_3), .o(n_3995) );
na02f80 g563748 ( .a(n_5824), .b(n_5929), .o(n_4754) );
na02f80 g563749 ( .a(n_6296), .b(FE_OFN27_n_13676), .o(n_7225) );
no02f80 g563750 ( .a(n_3993), .b(n_5281), .o(n_3994) );
no02f80 g563751 ( .a(n_5039), .b(n_2392), .o(n_3992) );
no02f80 g563752 ( .a(n_3018), .b(n_3292), .o(n_4753) );
na02f80 g563753 ( .a(n_3510), .b(x_in_49_0), .o(n_10920) );
na02f80 g563754 ( .a(n_4751), .b(x_in_1_3), .o(n_4752) );
na02f80 g563755 ( .a(n_4748), .b(n_5961), .o(n_4749) );
no02f80 g563756 ( .a(n_10553), .b(n_5961), .o(n_5194) );
no02f80 g563757 ( .a(n_5824), .b(n_2141), .o(n_4747) );
na02f80 g563758 ( .a(n_6528), .b(n_4746), .o(n_6293) );
na02f80 g563759 ( .a(n_4921), .b(n_4745), .o(n_6294) );
na02f80 g563760 ( .a(n_6524), .b(n_4329), .o(n_5711) );
na02f80 g563761 ( .a(n_6530), .b(n_4744), .o(n_6295) );
na02f80 g563762 ( .a(n_4772), .b(n_3363), .o(n_12281) );
no02f80 g563763 ( .a(n_5918), .b(n_4742), .o(n_4743) );
na02f80 g563764 ( .a(n_8157), .b(n_4740), .o(n_4331) );
no02f80 g563765 ( .a(n_8157), .b(n_4740), .o(n_4741) );
no02f80 g563766 ( .a(n_4739), .b(n_5192), .o(n_8195) );
na02f80 g563767 ( .a(n_6522), .b(n_4738), .o(n_6291) );
na02f80 g563768 ( .a(n_6526), .b(n_4737), .o(n_5712) );
in01f80 g563769 ( .a(n_6719), .o(n_4736) );
na02f80 g563770 ( .a(FE_OFN676_n_6824), .b(n_3364), .o(n_6719) );
na02f80 g563771 ( .a(n_5831), .b(n_5192), .o(n_5193) );
no02f80 g563772 ( .a(n_2993), .b(n_4734), .o(n_4735) );
no02f80 g563773 ( .a(n_8618), .b(n_4732), .o(n_4733) );
na02f80 g563774 ( .a(n_10048), .b(n_4057), .o(n_4731) );
in01f80 g563775 ( .a(n_6512), .o(n_10849) );
na02f80 g563776 ( .a(n_6521), .b(x_in_35_3), .o(n_6512) );
na02f80 g563777 ( .a(n_2895), .b(n_11148), .o(n_4730) );
in01f80 g563778 ( .a(n_4729), .o(n_6680) );
no02f80 g563779 ( .a(n_3370), .b(n_2078), .o(n_4729) );
no02f80 g563780 ( .a(n_4808), .b(x_in_0_1), .o(n_3991) );
no02f80 g563781 ( .a(n_3989), .b(x_in_3_0), .o(n_3990) );
na02f80 g563782 ( .a(n_4727), .b(x_in_45_15), .o(n_4728) );
no02f80 g563783 ( .a(n_4872), .b(x_in_4_1), .o(n_3520) );
in01f80 g563784 ( .a(n_5803), .o(n_5804) );
na02f80 g563785 ( .a(n_5191), .b(x_in_41_1), .o(n_5803) );
no02f80 g563786 ( .a(n_5850), .b(n_4725), .o(n_4726) );
no02f80 g563787 ( .a(n_2812), .b(n_2287), .o(n_4724) );
no02f80 g563788 ( .a(n_3602), .b(n_2288), .o(n_3521) );
na02f80 g563789 ( .a(n_4956), .b(n_3987), .o(n_3988) );
na02f80 g563790 ( .a(n_3488), .b(n_5161), .o(n_7170) );
no02f80 g563791 ( .a(n_9010), .b(n_7481), .o(n_4723) );
no02f80 g563792 ( .a(n_3985), .b(n_4722), .o(n_3986) );
na02f80 g563793 ( .a(n_3522), .b(n_4155), .o(n_3523) );
no02f80 g563794 ( .a(n_2897), .b(n_4155), .o(n_7118) );
no02f80 g563795 ( .a(n_2872), .b(n_4722), .o(n_7122) );
na02f80 g563796 ( .a(n_3524), .b(n_4719), .o(n_3525) );
no02f80 g563797 ( .a(n_3216), .b(n_4720), .o(n_7120) );
no02f80 g563798 ( .a(n_2896), .b(n_4719), .o(n_7116) );
na02f80 g563799 ( .a(n_3983), .b(n_4720), .o(n_3984) );
na02f80 g563800 ( .a(n_9146), .b(n_4717), .o(n_4718) );
no02f80 g563801 ( .a(n_3383), .b(x_in_27_6), .o(n_4974) );
na02f80 g563802 ( .a(n_5980), .b(n_4163), .o(n_4164) );
na02f80 g563803 ( .a(n_3981), .b(n_4716), .o(n_3982) );
no02f80 g563804 ( .a(n_2782), .b(n_4716), .o(n_7106) );
no02f80 g563805 ( .a(n_3529), .b(x_in_5_7), .o(n_5619) );
no02f80 g563806 ( .a(n_4714), .b(x_in_17_15), .o(n_4715) );
na02f80 g563807 ( .a(n_5099), .b(n_3978), .o(n_3979) );
na02f80 g563808 ( .a(n_2853), .b(n_6856), .o(n_4174) );
no02f80 g563809 ( .a(n_5076), .b(n_3558), .o(n_3559) );
no02f80 g563810 ( .a(n_3400), .b(n_3399), .o(n_3401) );
na02f80 g563811 ( .a(n_3536), .b(n_3535), .o(n_3537) );
na02f80 g563812 ( .a(n_2779), .b(n_11168), .o(n_4713) );
na02f80 g563813 ( .a(n_3531), .b(n_3530), .o(n_3532) );
no02f80 g563814 ( .a(n_3975), .b(n_7099), .o(n_3976) );
na02f80 g563815 ( .a(FE_OFN933_n_4950), .b(x_in_51_15), .o(n_3974) );
no02f80 g563816 ( .a(n_3533), .b(n_7102), .o(n_3534) );
no02f80 g563817 ( .a(n_5189), .b(n_6641), .o(n_5190) );
no02f80 g563818 ( .a(n_4182), .b(x_in_25_1), .o(n_4712) );
in01f80 g563819 ( .a(n_5187), .o(n_5188) );
na02f80 g563820 ( .a(n_4182), .b(x_in_25_1), .o(n_5187) );
no02f80 g563821 ( .a(n_2731), .b(n_5308), .o(n_8365) );
na02f80 g563822 ( .a(n_3538), .b(n_5308), .o(n_3539) );
no02f80 g563823 ( .a(n_4710), .b(n_5902), .o(n_4711) );
na02f80 g563824 ( .a(n_5367), .b(n_3971), .o(n_3972) );
na02f80 g563825 ( .a(n_2836), .b(FE_OFN973_n_6822), .o(n_4709) );
no02f80 g563826 ( .a(n_9082), .b(n_7551), .o(n_3540) );
na02f80 g563827 ( .a(n_4760), .b(n_4707), .o(n_4708) );
no02f80 g563828 ( .a(n_4706), .b(n_4027), .o(n_7096) );
no02f80 g563829 ( .a(n_3404), .b(x_in_43_7), .o(n_5608) );
na02f80 g563830 ( .a(n_3969), .b(n_3968), .o(n_3970) );
na02f80 g563831 ( .a(n_3062), .b(n_10220), .o(n_4705) );
no02f80 g563832 ( .a(n_3476), .b(n_4967), .o(n_4968) );
no02f80 g563833 ( .a(n_4123), .b(n_5185), .o(n_5186) );
no02f80 g563834 ( .a(n_3337), .b(n_4352), .o(n_7093) );
na02f80 g563835 ( .a(n_3548), .b(n_4352), .o(n_3549) );
na02f80 g563836 ( .a(n_5223), .b(n_4203), .o(n_4204) );
na02f80 g563837 ( .a(n_3546), .b(n_3545), .o(n_3547) );
na02f80 g563838 ( .a(n_3059), .b(FE_OFN971_n_6854), .o(n_4704) );
no02f80 g563839 ( .a(n_3320), .b(n_4355), .o(n_4356) );
no02f80 g563840 ( .a(n_4702), .b(n_6653), .o(n_4703) );
no02f80 g563841 ( .a(n_3966), .b(n_4903), .o(n_3967) );
no02f80 g563842 ( .a(n_10020), .b(n_3551), .o(n_3552) );
no02f80 g563843 ( .a(n_4977), .b(n_4976), .o(n_4978) );
na02f80 g563844 ( .a(n_3964), .b(n_3963), .o(n_3965) );
no02f80 g563845 ( .a(n_3961), .b(x_in_35_15), .o(n_3962) );
na02f80 g563846 ( .a(n_3554), .b(x_in_11_1), .o(n_3555) );
no02f80 g563847 ( .a(n_3959), .b(x_in_43_1), .o(n_3960) );
in01f80 g563848 ( .a(n_9543), .o(n_5183) );
no02f80 g563849 ( .a(n_5852), .b(n_7653), .o(n_9543) );
na02f80 g563850 ( .a(n_4700), .b(n_5938), .o(n_4701) );
no02f80 g563851 ( .a(n_5928), .b(n_4698), .o(n_4699) );
no02f80 g563852 ( .a(n_10013), .b(n_8485), .o(n_5182) );
na02f80 g563853 ( .a(n_2847), .b(n_4358), .o(n_4359) );
na02f80 g563854 ( .a(n_4706), .b(n_4228), .o(n_4229) );
na02f80 g563855 ( .a(n_4696), .b(n_5820), .o(n_4697) );
no02f80 g563856 ( .a(n_10007), .b(n_3957), .o(n_3958) );
no02f80 g563857 ( .a(n_3658), .b(n_4694), .o(n_4695) );
na02f80 g563858 ( .a(n_4230), .b(n_6781), .o(n_10847) );
na02f80 g563859 ( .a(n_10820), .b(n_6359), .o(n_5181) );
no02f80 g563860 ( .a(n_5821), .b(n_5180), .o(n_10887) );
no02f80 g563861 ( .a(n_4655), .b(x_in_37_3), .o(n_4362) );
na02f80 g563862 ( .a(n_3955), .b(n_3954), .o(n_3956) );
na02f80 g563863 ( .a(FE_OFN1188_n_5249), .b(x_in_7_1), .o(n_10885) );
no02f80 g563864 ( .a(FE_OFN1188_n_5249), .b(x_in_7_1), .o(n_3557) );
na02f80 g563865 ( .a(n_3952), .b(x_in_7_1), .o(n_3953) );
na02f80 g563866 ( .a(n_5425), .b(x_in_21_15), .o(n_5426) );
na02f80 g563867 ( .a(n_3457), .b(x_in_59_1), .o(n_3458) );
na02f80 g563868 ( .a(n_5232), .b(n_4692), .o(n_4693) );
na02f80 g563869 ( .a(n_5229), .b(n_5231), .o(n_4691) );
na02f80 g563870 ( .a(n_3950), .b(n_3949), .o(n_3951) );
no02f80 g563871 ( .a(n_3947), .b(n_3946), .o(n_3948) );
na02f80 g563872 ( .a(n_3057), .b(n_4289), .o(n_4290) );
na02f80 g563873 ( .a(n_5225), .b(n_5228), .o(n_4262) );
na02f80 g563874 ( .a(n_5227), .b(n_5224), .o(n_4690) );
no02f80 g563875 ( .a(n_3944), .b(n_3943), .o(n_3945) );
na02f80 g563876 ( .a(n_2899), .b(n_4688), .o(n_4689) );
na02f80 g563877 ( .a(n_3465), .b(n_3464), .o(n_3466) );
na02f80 g563878 ( .a(n_3473), .b(n_3472), .o(n_3474) );
no02f80 g563879 ( .a(n_3657), .b(x_in_29_10), .o(n_4263) );
in01f80 g563880 ( .a(n_5178), .o(n_5179) );
no02f80 g563881 ( .a(n_5853), .b(n_4687), .o(n_5178) );
na02f80 g563882 ( .a(n_2926), .b(FE_OFN676_n_6824), .o(n_4686) );
na02f80 g563883 ( .a(n_3564), .b(n_3563), .o(n_3565) );
na02f80 g563884 ( .a(n_2916), .b(n_4264), .o(n_4265) );
na02f80 g563885 ( .a(n_3940), .b(x_in_27_2), .o(n_3941) );
na02f80 g563886 ( .a(FE_OFN1073_n_6399), .b(x_in_61_0), .o(n_9987) );
na02f80 g563887 ( .a(n_11201), .b(x_in_53_0), .o(n_8562) );
in01f80 g563888 ( .a(n_4685), .o(n_10872) );
na02f80 g563889 ( .a(n_3566), .b(n_5848), .o(n_4685) );
na02f80 g563890 ( .a(n_3938), .b(x_in_9_15), .o(n_3939) );
na02f80 g563891 ( .a(n_3486), .b(x_in_51_14), .o(n_3487) );
na02f80 g563892 ( .a(n_3936), .b(x_in_11_2), .o(n_3937) );
na02f80 g563893 ( .a(n_3934), .b(x_in_11_14), .o(n_3935) );
na02f80 g563894 ( .a(n_3932), .b(x_in_37_15), .o(n_3933) );
na02f80 g563895 ( .a(n_3502), .b(x_in_43_2), .o(n_3503) );
na02f80 g563896 ( .a(n_3930), .b(x_in_27_1), .o(n_3931) );
na02f80 g563897 ( .a(n_3928), .b(n_3927), .o(n_3929) );
na02f80 g563898 ( .a(n_5443), .b(n_4317), .o(n_4318) );
no02f80 g563899 ( .a(n_3925), .b(x_in_49_4), .o(n_3926) );
na02f80 g563900 ( .a(n_4683), .b(n_5319), .o(n_4684) );
no02f80 g563901 ( .a(n_3365), .b(n_5176), .o(n_5177) );
na02f80 g563902 ( .a(n_3394), .b(n_4737), .o(n_5175) );
na02f80 g563903 ( .a(n_3682), .b(n_4329), .o(n_5174) );
na02f80 g563904 ( .a(n_3684), .b(n_4746), .o(n_5055) );
na02f80 g563905 ( .a(n_3683), .b(n_4745), .o(n_5038) );
na02f80 g563906 ( .a(n_3685), .b(n_4744), .o(n_5173) );
na02f80 g563907 ( .a(n_4120), .b(n_4738), .o(n_5172) );
no02f80 g563908 ( .a(n_5261), .b(n_3146), .o(n_3506) );
no02f80 g563909 ( .a(n_5261), .b(n_5342), .o(n_3924) );
na02f80 g563910 ( .a(n_8734), .b(n_6709), .o(n_4682) );
na02f80 g563911 ( .a(n_3922), .b(x_in_3_14), .o(n_3923) );
na02f80 g563912 ( .a(n_3513), .b(x_in_11_3), .o(n_3514) );
no02f80 g563913 ( .a(n_3493), .b(n_5170), .o(n_5171) );
na02f80 g563914 ( .a(n_8731), .b(n_6715), .o(n_5169) );
na02f80 g563915 ( .a(n_3571), .b(x_in_59_14), .o(n_3572) );
in01f80 g563916 ( .a(n_6725), .o(n_4681) );
no02f80 g563917 ( .a(n_3518), .b(n_4948), .o(n_6725) );
na02f80 g563918 ( .a(n_3920), .b(x_in_43_3), .o(n_3921) );
na02f80 g563920 ( .a(n_3916), .b(n_2277), .o(n_7043) );
na02f80 g563921 ( .a(n_3916), .b(n_5267), .o(n_3579) );
na02f80 g563923 ( .a(n_2328), .b(n_3424), .o(n_4332) );
no02f80 g563924 ( .a(n_5826), .b(x_in_3_3), .o(n_4334) );
na02f80 g563925 ( .a(n_5837), .b(x_in_21_1), .o(n_5168) );
na02f80 g563926 ( .a(n_4341), .b(n_3746), .o(n_4342) );
no02f80 g563927 ( .a(n_5943), .b(x_in_21_13), .o(n_4335) );
na02f80 g563928 ( .a(n_8728), .b(FE_OFN692_n_6708), .o(n_5043) );
na02f80 g563929 ( .a(n_2972), .b(n_4343), .o(n_4344) );
no02f80 g563930 ( .a(n_3494), .b(n_5166), .o(n_5167) );
no02f80 g563931 ( .a(n_4956), .b(x_in_35_2), .o(n_3544) );
na02f80 g563932 ( .a(n_5269), .b(x_in_59_2), .o(n_3574) );
no02f80 g563933 ( .a(n_3414), .b(x_in_39_10), .o(n_5045) );
in01f80 g563934 ( .a(n_5164), .o(n_5165) );
na02f80 g563935 ( .a(n_4347), .b(x_in_37_13), .o(n_5164) );
na02f80 g563936 ( .a(n_5163), .b(n_4343), .o(n_7204) );
na02f80 g563937 ( .a(n_3866), .b(x_in_37_13), .o(n_3541) );
na02f80 g563938 ( .a(n_3577), .b(x_in_37_14), .o(n_3578) );
no02f80 g563939 ( .a(n_3542), .b(x_in_5_3), .o(n_9982) );
in01f80 g563940 ( .a(n_4680), .o(n_10864) );
na02f80 g563941 ( .a(n_3989), .b(n_4419), .o(n_4680) );
na02f80 g563942 ( .a(n_5930), .b(x_in_3_2), .o(n_6030) );
no02f80 g563943 ( .a(n_5478), .b(x_in_17_5), .o(n_4360) );
no02f80 g563944 ( .a(n_5049), .b(n_5048), .o(n_5050) );
no02f80 g563945 ( .a(n_6576), .b(n_5161), .o(n_5162) );
no02f80 g563946 ( .a(n_4998), .b(x_in_17_10), .o(n_4679) );
no02f80 g563947 ( .a(n_5740), .b(x_in_37_6), .o(n_4357) );
no02f80 g563948 ( .a(n_3596), .b(n_5884), .o(n_5054) );
no02f80 g563949 ( .a(n_3008), .b(x_in_21_12), .o(n_6763) );
no02f80 g563950 ( .a(n_3436), .b(n_4677), .o(n_4678) );
na02f80 g563951 ( .a(n_5253), .b(x_in_19_3), .o(n_10856) );
na02f80 g563952 ( .a(n_3620), .b(x_in_19_14), .o(n_3621) );
no02f80 g563953 ( .a(n_5669), .b(x_in_17_3), .o(n_3915) );
na02f80 g563954 ( .a(n_3613), .b(x_in_49_3), .o(n_3614) );
no02f80 g563955 ( .a(n_4655), .b(n_4376), .o(n_4377) );
no02f80 g563956 ( .a(n_3009), .b(n_5977), .o(n_6764) );
no02f80 g563957 ( .a(n_3649), .b(n_5159), .o(n_5160) );
na02f80 g563958 ( .a(n_5880), .b(x_in_37_4), .o(n_4676) );
no02f80 g563959 ( .a(n_5780), .b(n_4037), .o(n_5781) );
na02f80 g563960 ( .a(n_5740), .b(x_in_37_2), .o(n_4378) );
na02f80 g563961 ( .a(n_11201), .b(x_in_53_1), .o(n_12820) );
na02f80 g563962 ( .a(n_7602), .b(x_in_61_1), .o(n_4382) );
no02f80 g563963 ( .a(n_3912), .b(x_in_49_10), .o(n_3913) );
na02f80 g563964 ( .a(n_3653), .b(x_in_49_8), .o(n_3654) );
na02f80 g563965 ( .a(n_3911), .b(x_in_57_4), .o(n_7020) );
no02f80 g563966 ( .a(n_3909), .b(x_in_57_3), .o(n_3910) );
no02f80 g563967 ( .a(n_3726), .b(x_in_49_6), .o(n_3727) );
no02f80 g563968 ( .a(n_2730), .b(x_in_57_3), .o(n_9967) );
na02f80 g563969 ( .a(n_4084), .b(x_in_11_5), .o(n_4085) );
na02f80 g563970 ( .a(n_3907), .b(x_in_61_1), .o(n_3908) );
na02f80 g563971 ( .a(n_3584), .b(x_in_49_7), .o(n_3585) );
na02f80 g563972 ( .a(n_9120), .b(n_4674), .o(n_4675) );
no02f80 g563973 ( .a(n_4128), .b(n_5068), .o(n_5069) );
no02f80 g563974 ( .a(n_5036), .b(x_in_5_7), .o(n_3590) );
na02f80 g563975 ( .a(n_3778), .b(x_in_27_3), .o(n_3779) );
no02f80 g563976 ( .a(FE_OFN1073_n_6399), .b(x_in_61_1), .o(n_3768) );
na02f80 g563977 ( .a(FE_OFN1073_n_6399), .b(x_in_61_1), .o(n_10851) );
na02f80 g563978 ( .a(n_7419), .b(n_4672), .o(n_4673) );
na02f80 g563979 ( .a(n_5751), .b(x_in_21_7), .o(n_4517) );
in01f80 g563980 ( .a(n_4510), .o(n_6271) );
no02f80 g563981 ( .a(n_2441), .b(n_9207), .o(n_4510) );
na02f80 g563982 ( .a(n_5922), .b(x_in_21_7), .o(n_4671) );
na02f80 g563983 ( .a(n_4669), .b(n_4668), .o(n_4670) );
na02f80 g563984 ( .a(n_5411), .b(n_3318), .o(n_4528) );
no02f80 g563985 ( .a(n_5305), .b(x_in_57_8), .o(n_3905) );
na02f80 g563986 ( .a(n_5391), .b(x_in_61_12), .o(n_3790) );
no02f80 g563987 ( .a(n_3602), .b(x_in_35_1), .o(n_3603) );
na02f80 g563988 ( .a(n_5157), .b(n_5156), .o(n_5158) );
no02f80 g563989 ( .a(n_5918), .b(x_in_51_2), .o(n_4169) );
na02f80 g563990 ( .a(n_3604), .b(x_in_33_5), .o(n_5432) );
no02f80 g563991 ( .a(n_5306), .b(x_in_57_6), .o(n_3904) );
na02f80 g563992 ( .a(n_4025), .b(x_in_43_5), .o(n_4026) );
no02f80 g563993 ( .a(n_5409), .b(x_in_37_7), .o(n_4368) );
na02f80 g563994 ( .a(n_5062), .b(x_in_37_7), .o(n_5063) );
na02f80 g563995 ( .a(n_3814), .b(x_in_59_9), .o(n_3815) );
na02f80 g563996 ( .a(n_5943), .b(x_in_21_9), .o(n_4666) );
na02f80 g563997 ( .a(n_5801), .b(n_9961), .o(n_5802) );
no02f80 g563998 ( .a(n_5934), .b(n_4664), .o(n_4665) );
no02f80 g563999 ( .a(n_3016), .b(n_4579), .o(n_4580) );
no02f80 g564000 ( .a(n_6573), .b(n_5153), .o(n_5154) );
na02f80 g564001 ( .a(n_3824), .b(x_in_59_5), .o(n_3825) );
na02f80 g564002 ( .a(n_2923), .b(n_3608), .o(n_3609) );
na02f80 g564003 ( .a(n_4101), .b(x_in_37_5), .o(n_5151) );
na02f80 g564004 ( .a(n_5732), .b(x_in_3_6), .o(n_6014) );
na02f80 g564005 ( .a(n_5149), .b(n_9958), .o(n_5150) );
na02f80 g564006 ( .a(n_5934), .b(x_in_19_5), .o(n_4886) );
na02f80 g564007 ( .a(n_4662), .b(n_5703), .o(n_4663) );
na02f80 g564008 ( .a(n_4936), .b(x_in_51_3), .o(n_4114) );
na02f80 g564009 ( .a(n_2924), .b(x_in_61_3), .o(n_4896) );
na02f80 g564010 ( .a(n_5956), .b(x_in_3_8), .o(n_6001) );
na02f80 g564011 ( .a(n_3918), .b(x_in_53_4), .o(n_3901) );
na02f80 g564012 ( .a(n_5277), .b(x_in_25_4), .o(n_3423) );
na02f80 g564013 ( .a(n_4640), .b(n_5742), .o(n_4371) );
no02f80 g564014 ( .a(n_4132), .b(n_8191), .o(n_4133) );
na02f80 g564015 ( .a(n_3276), .b(n_4660), .o(n_4661) );
no02f80 g564016 ( .a(n_5854), .b(n_5074), .o(n_5075) );
no02f80 g564017 ( .a(n_6216), .b(n_4659), .o(n_8358) );
no02f80 g564018 ( .a(n_3618), .b(n_3617), .o(n_3619) );
no02f80 g564019 ( .a(n_4015), .b(n_3516), .o(n_3517) );
na02f80 g564020 ( .a(n_3455), .b(x_in_61_7), .o(n_3456) );
no02f80 g564021 ( .a(n_5799), .b(n_3361), .o(n_5800) );
na02f80 g564022 ( .a(n_5076), .b(x_in_35_5), .o(n_3471) );
na02f80 g564023 ( .a(n_3624), .b(x_in_53_14), .o(n_3625) );
no02f80 g564024 ( .a(n_3989), .b(n_5825), .o(n_10839) );
na02f80 g564025 ( .a(n_3418), .b(x_in_59_3), .o(n_3419) );
no02f80 g564026 ( .a(n_3622), .b(x_in_37_8), .o(n_3623) );
no02f80 g564027 ( .a(n_8561), .b(n_4657), .o(n_4658) );
no02f80 g564028 ( .a(n_5797), .b(n_4070), .o(n_5798) );
na02f80 g564029 ( .a(n_4139), .b(n_4138), .o(n_4140) );
na02f80 g564030 ( .a(n_5874), .b(x_in_3_4), .o(n_6010) );
no02f80 g564031 ( .a(n_4206), .b(n_4205), .o(n_4207) );
na02f80 g564032 ( .a(n_5771), .b(n_5431), .o(n_5148) );
no02f80 g564033 ( .a(n_4341), .b(x_in_21_5), .o(n_4147) );
na02f80 g564034 ( .a(n_3897), .b(x_in_27_5), .o(n_3898) );
na02f80 g564035 ( .a(n_3680), .b(n_4180), .o(n_4181) );
na02f80 g564036 ( .a(n_5146), .b(FE_OFN612_n_5698), .o(n_5147) );
in01f80 g564037 ( .a(n_9932), .o(n_4656) );
na02f80 g564038 ( .a(n_5322), .b(n_3387), .o(n_9932) );
na02f80 g564039 ( .a(n_3896), .b(x_in_33_4), .o(n_5427) );
na02f80 g564040 ( .a(n_3626), .b(x_in_61_8), .o(n_3627) );
na02f80 g564041 ( .a(n_3894), .b(x_in_61_9), .o(n_3895) );
no02f80 g564042 ( .a(n_4149), .b(n_4148), .o(n_4150) );
na02f80 g564043 ( .a(n_4655), .b(n_4654), .o(n_10777) );
na02f80 g564044 ( .a(n_4700), .b(n_7765), .o(n_4219) );
no02f80 g564045 ( .a(n_4652), .b(n_4651), .o(n_4653) );
no02f80 g564046 ( .a(n_5616), .b(x_in_17_7), .o(n_4208) );
na02f80 g564047 ( .a(n_4927), .b(x_in_51_5), .o(n_3893) );
na02f80 g564048 ( .a(n_3636), .b(x_in_33_10), .o(n_5423) );
na02f80 g564049 ( .a(n_4969), .b(x_in_33_9), .o(n_6636) );
na02f80 g564050 ( .a(n_3891), .b(x_in_33_8), .o(n_5064) );
na02f80 g564051 ( .a(n_3403), .b(x_in_33_7), .o(n_5422) );
na02f80 g564052 ( .a(n_3359), .b(x_in_33_6), .o(n_5424) );
na02f80 g564053 ( .a(FE_OFN933_n_4950), .b(x_in_51_9), .o(n_5421) );
na02f80 g564054 ( .a(n_5144), .b(n_7434), .o(n_5145) );
na02f80 g564055 ( .a(n_4821), .b(x_in_25_9), .o(n_3371) );
no02f80 g564056 ( .a(n_5611), .b(x_in_17_9), .o(n_4154) );
na02f80 g564057 ( .a(n_10216), .b(n_5827), .o(n_5143) );
na02f80 g564058 ( .a(n_5299), .b(x_in_21_2), .o(n_4152) );
na02f80 g564059 ( .a(n_3435), .b(n_7434), .o(n_4918) );
no02f80 g564060 ( .a(n_7648), .b(x_in_33_12), .o(n_4153) );
na02f80 g564061 ( .a(n_12697), .b(x_in_33_11), .o(n_5759) );
in01f80 g564062 ( .a(n_11346), .o(n_5142) );
na02f80 g564063 ( .a(n_2766), .b(n_4386), .o(n_11346) );
no02f80 g564064 ( .a(n_4924), .b(n_4923), .o(n_4925) );
na02f80 g564065 ( .a(n_8287), .b(x_in_17_4), .o(n_3690) );
no02f80 g564066 ( .a(n_3593), .b(x_in_17_4), .o(n_4650) );
no02f80 g564067 ( .a(n_8287), .b(n_4021), .o(n_7838) );
no02f80 g564068 ( .a(n_5140), .b(x_in_3_13), .o(n_5141) );
na02f80 g564069 ( .a(n_3637), .b(n_5866), .o(n_5139) );
no02f80 g564070 ( .a(n_3376), .b(n_5868), .o(n_3377) );
na02f80 g564071 ( .a(n_4953), .b(n_9896), .o(n_4954) );
no02f80 g564072 ( .a(n_3586), .b(x_in_17_8), .o(n_4649) );
no02f80 g564073 ( .a(n_3589), .b(x_in_17_6), .o(n_4648) );
no02f80 g564074 ( .a(n_4915), .b(n_4397), .o(n_4398) );
na02f80 g564075 ( .a(n_4793), .b(n_5226), .o(n_3515) );
na02f80 g564076 ( .a(n_3889), .b(n_8336), .o(n_3890) );
no02f80 g564077 ( .a(n_4041), .b(x_in_21_3), .o(n_4931) );
no02f80 g564078 ( .a(n_4040), .b(n_6781), .o(n_4647) );
in01f80 g564079 ( .a(n_4933), .o(n_4934) );
na02f80 g564080 ( .a(n_4160), .b(n_2476), .o(n_4933) );
na02f80 g564081 ( .a(n_6573), .b(n_5137), .o(n_5138) );
no02f80 g564082 ( .a(n_5795), .b(x_in_17_13), .o(n_5796) );
na02f80 g564083 ( .a(n_6958), .b(x_in_51_11), .o(n_6628) );
no02f80 g564084 ( .a(n_4160), .b(n_4159), .o(n_4161) );
na02f80 g564085 ( .a(n_5135), .b(n_3277), .o(n_5136) );
na02f80 g564086 ( .a(n_4714), .b(n_4176), .o(n_4177) );
in01f80 g564087 ( .a(n_6775), .o(n_5134) );
no02f80 g564088 ( .a(n_6219), .b(n_4146), .o(n_6775) );
na02f80 g564089 ( .a(n_6219), .b(n_4146), .o(n_6777) );
na02f80 g564090 ( .a(n_5132), .b(n_6425), .o(n_5133) );
na02f80 g564091 ( .a(n_4183), .b(n_4172), .o(n_4173) );
na02f80 g564092 ( .a(n_4646), .b(n_4645), .o(n_9426) );
na02f80 g564093 ( .a(n_3553), .b(n_5130), .o(n_7865) );
no02f80 g564094 ( .a(n_6563), .b(n_5130), .o(n_5131) );
in01f80 g564095 ( .a(n_5128), .o(n_5129) );
no02f80 g564096 ( .a(n_7499), .b(n_2808), .o(n_5128) );
no02f80 g564097 ( .a(n_7498), .b(n_2411), .o(n_6648) );
na02f80 g564098 ( .a(n_6707), .b(n_8701), .o(n_3884) );
in01f80 g564099 ( .a(n_5793), .o(n_5794) );
na02f80 g564100 ( .a(n_3581), .b(n_4957), .o(n_5793) );
na02f80 g564101 ( .a(n_3580), .b(n_4232), .o(n_6646) );
na02f80 g564102 ( .a(n_5482), .b(n_2437), .o(n_6443) );
no02f80 g564103 ( .a(n_4183), .b(n_2443), .o(n_7751) );
na02f80 g564104 ( .a(n_5822), .b(n_5251), .o(n_11524) );
in01f80 g564105 ( .a(n_8896), .o(n_5792) );
no02f80 g564106 ( .a(n_4959), .b(n_4958), .o(n_8896) );
na02f80 g564107 ( .a(n_4867), .b(n_2390), .o(n_5791) );
in01f80 g564108 ( .a(n_4962), .o(n_4963) );
na02f80 g564109 ( .a(n_5436), .b(n_2857), .o(n_4962) );
na02f80 g564110 ( .a(n_4960), .b(n_2662), .o(n_6647) );
na02f80 g564111 ( .a(n_3774), .b(n_3773), .o(n_3775) );
no02f80 g564112 ( .a(n_5269), .b(n_5268), .o(n_3883) );
na02f80 g564113 ( .a(n_4643), .b(n_4642), .o(n_4644) );
in01f80 g564114 ( .a(n_7599), .o(n_5760) );
no02f80 g564115 ( .a(n_5476), .b(n_5127), .o(n_7599) );
no02f80 g564116 ( .a(n_4640), .b(n_4639), .o(n_4641) );
na02f80 g564117 ( .a(n_3828), .b(n_3827), .o(n_3829) );
na02f80 g564118 ( .a(n_4367), .b(n_5790), .o(n_8324) );
na02f80 g564119 ( .a(n_3475), .b(n_5126), .o(n_7744) );
na02f80 g564120 ( .a(n_6437), .b(n_4213), .o(n_4214) );
no02f80 g564121 ( .a(n_3425), .b(n_2374), .o(n_3426) );
no02f80 g564122 ( .a(n_4638), .b(n_2508), .o(n_7743) );
na02f80 g564123 ( .a(n_4638), .b(n_4636), .o(n_4637) );
na02f80 g564124 ( .a(n_4634), .b(n_5125), .o(n_4635) );
no02f80 g564125 ( .a(n_3597), .b(n_5125), .o(n_7742) );
in01f80 g564126 ( .a(n_8892), .o(n_5124) );
no02f80 g564127 ( .a(n_6209), .b(n_4220), .o(n_8892) );
no02f80 g564128 ( .a(FE_OFN1234_n_4979), .b(n_3796), .o(n_3797) );
in01f80 g564129 ( .a(n_4632), .o(n_4633) );
na02f80 g564130 ( .a(FE_OFN1234_n_4979), .b(n_5401), .o(n_4632) );
na02f80 g564131 ( .a(n_3582), .b(n_4980), .o(n_7738) );
no02f80 g564132 ( .a(n_4643), .b(n_2447), .o(n_6910) );
no02f80 g564133 ( .a(n_6571), .b(n_4980), .o(n_4981) );
na02f80 g564134 ( .a(n_4630), .b(n_8693), .o(n_4631) );
no02f80 g564135 ( .a(n_5123), .b(n_3477), .o(n_10810) );
na02f80 g564136 ( .a(n_5121), .b(n_5790), .o(n_5122) );
na02f80 g564137 ( .a(n_4236), .b(n_4226), .o(n_4227) );
no02f80 g564138 ( .a(n_4109), .b(n_2564), .o(n_6461) );
no02f80 g564139 ( .a(n_6204), .b(n_3045), .o(n_6776) );
na02f80 g564140 ( .a(n_4554), .b(n_5126), .o(n_4555) );
in01f80 g564141 ( .a(n_7489), .o(n_5120) );
no02f80 g564142 ( .a(n_4629), .b(n_2472), .o(n_7489) );
no02f80 g564143 ( .a(n_4629), .b(n_5904), .o(n_4235) );
in01f80 g564144 ( .a(n_5118), .o(n_5119) );
na02f80 g564145 ( .a(n_4236), .b(n_2316), .o(n_5118) );
no02f80 g564146 ( .a(n_6437), .b(n_2498), .o(n_7763) );
no02f80 g564147 ( .a(n_5384), .b(n_5383), .o(n_3882) );
na02f80 g564148 ( .a(FE_OFN1184_n_6701), .b(n_8690), .o(n_3835) );
no02f80 g564149 ( .a(n_7474), .b(n_3643), .o(n_6651) );
na02f80 g564150 ( .a(n_4627), .b(n_4626), .o(n_4628) );
na02f80 g564151 ( .a(n_4624), .b(n_4623), .o(n_4625) );
na02f80 g564152 ( .a(n_4248), .b(n_4247), .o(n_4249) );
na02f80 g564153 ( .a(n_5855), .b(n_4253), .o(n_4254) );
na02f80 g564154 ( .a(n_5928), .b(n_4621), .o(n_4622) );
no02f80 g564155 ( .a(n_5913), .b(n_4997), .o(n_4620) );
na02f80 g564156 ( .a(n_3357), .b(n_4997), .o(n_8013) );
na02f80 g564157 ( .a(n_3462), .b(n_4903), .o(n_26869) );
no02f80 g564158 ( .a(n_6204), .b(n_4618), .o(n_4619) );
no02f80 g564159 ( .a(n_5116), .b(n_5115), .o(n_5117) );
na02f80 g564160 ( .a(n_4876), .b(n_5772), .o(n_5773) );
na02f80 g564161 ( .a(n_5645), .b(n_3326), .o(n_19015) );
in01f80 g564162 ( .a(n_5113), .o(n_5114) );
na02f80 g564163 ( .a(n_5685), .b(n_3019), .o(n_5113) );
na02f80 g564164 ( .a(n_3880), .b(n_3879), .o(n_3881) );
no02f80 g564165 ( .a(n_5873), .b(n_4616), .o(n_4617) );
in01f80 g564166 ( .a(n_4266), .o(n_4267) );
na02f80 g564167 ( .a(n_3880), .b(n_2609), .o(n_4266) );
no02f80 g564168 ( .a(n_4615), .b(n_4089), .o(n_7720) );
na02f80 g564169 ( .a(n_4615), .b(n_4291), .o(n_4292) );
no02f80 g564170 ( .a(n_5116), .b(n_3592), .o(n_8301) );
na02f80 g564171 ( .a(n_5391), .b(n_3885), .o(n_3886) );
na02f80 g564172 ( .a(n_4613), .b(n_2398), .o(n_4614) );
no02f80 g564173 ( .a(n_4991), .b(n_4121), .o(n_3489) );
na02f80 g564174 ( .a(n_9032), .b(n_3878), .o(n_6203) );
in01f80 g564175 ( .a(n_4611), .o(n_4612) );
no02f80 g564176 ( .a(n_9032), .b(n_3878), .o(n_4611) );
na02f80 g564177 ( .a(n_5916), .b(n_3039), .o(n_4610) );
no02f80 g564178 ( .a(n_5916), .b(n_4323), .o(n_4324) );
no02f80 g564179 ( .a(n_3899), .b(n_2361), .o(n_3900) );
no02f80 g564180 ( .a(n_4852), .b(n_5789), .o(n_7686) );
na02f80 g564181 ( .a(n_5111), .b(n_5789), .o(n_5112) );
na02f80 g564182 ( .a(n_6081), .b(n_13676), .o(n_7409) );
na02f80 g564184 ( .a(n_4609), .b(n_4608), .o(n_9424) );
in01f80 g564185 ( .a(n_6338), .o(n_3906) );
oa12f80 g564186 ( .a(n_2714), .b(n_2713), .c(x_in_37_5), .o(n_6338) );
in01f80 g564187 ( .a(n_6334), .o(n_3877) );
oa12f80 g564188 ( .a(n_2733), .b(n_2732), .c(x_in_37_9), .o(n_6334) );
in01f80 g564189 ( .a(n_5788), .o(n_11860) );
na02f80 g564190 ( .a(n_6580), .b(n_5039), .o(n_5788) );
na02f80 g564191 ( .a(n_4820), .b(n_3527), .o(n_3528) );
na02f80 g564192 ( .a(n_4606), .b(n_4605), .o(n_4607) );
ao12f80 g564193 ( .a(n_3876), .b(n_2610), .c(x_in_41_6), .o(n_5643) );
oa12f80 g564194 ( .a(n_2057), .b(n_3207), .c(x_in_61_2), .o(n_6047) );
na02f80 g564195 ( .a(n_4598), .b(n_4336), .o(n_4337) );
in01f80 g564196 ( .a(n_5662), .o(n_3874) );
oa12f80 g564197 ( .a(n_2939), .b(n_2938), .c(x_in_51_0), .o(n_5662) );
oa12f80 g564198 ( .a(n_4097), .b(n_2625), .c(x_in_39_15), .o(n_8787) );
no02f80 g564199 ( .a(n_3181), .b(n_4604), .o(n_12342) );
no02f80 g564202 ( .a(n_3573), .b(n_5108), .o(n_7626) );
na03f80 g564203 ( .a(x_in_35_0), .b(n_5832), .c(x_in_35_2), .o(n_14103) );
na03f80 g564204 ( .a(x_in_17_0), .b(n_4772), .c(x_in_17_1), .o(n_14115) );
ao12f80 g564206 ( .a(n_3869), .b(n_3868), .c(x_in_41_4), .o(n_5640) );
ao12f80 g564207 ( .a(n_7215), .b(n_2617), .c(x_in_41_8), .o(n_5646) );
na02f80 g564208 ( .a(n_3866), .b(n_8441), .o(n_3867) );
na02f80 g564209 ( .a(n_4606), .b(n_2883), .o(n_8280) );
in01f80 g564210 ( .a(n_4353), .o(n_4354) );
na02f80 g564211 ( .a(FE_OFN552_n_9482), .b(n_4455), .o(n_4353) );
na02f80 g564212 ( .a(n_4603), .b(n_4454), .o(n_5729) );
in01f80 g564213 ( .a(n_3865), .o(n_5652) );
oa12f80 g564214 ( .a(n_2939), .b(n_2938), .c(x_in_51_1), .o(n_3865) );
in01f80 g564215 ( .a(n_6297), .o(n_6451) );
na03f80 g564216 ( .a(n_7987), .b(n_2299), .c(n_2320), .o(n_6297) );
ao12f80 g564217 ( .a(n_3864), .b(n_7855), .c(x_in_35_4), .o(n_6371) );
no02f80 g564219 ( .a(n_5109), .b(n_5108), .o(n_5110) );
oa12f80 g564220 ( .a(n_3170), .b(n_4602), .c(n_4601), .o(n_7973) );
ao12f80 g564221 ( .a(n_2740), .b(n_2362), .c(x_in_45_1), .o(n_7191) );
na02f80 g564222 ( .a(n_4599), .b(n_5107), .o(n_4600) );
no02f80 g564223 ( .a(n_3495), .b(n_5107), .o(n_7624) );
oa12f80 g564224 ( .a(n_3993), .b(n_2851), .c(n_2573), .o(n_7961) );
oa12f80 g564225 ( .a(n_2724), .b(n_2723), .c(x_in_7_2), .o(n_6389) );
no02f80 g564226 ( .a(FE_OFN845_n_7616), .b(n_4604), .o(n_3862) );
no02f80 g564227 ( .a(n_4598), .b(n_3725), .o(n_7390) );
no02f80 g564228 ( .a(n_3860), .b(n_3859), .o(n_3861) );
ao12f80 g564229 ( .a(n_2042), .b(n_3143), .c(x_in_33_14), .o(n_8453) );
in01f80 g564230 ( .a(n_4830), .o(n_3858) );
oa12f80 g564231 ( .a(n_5700), .b(n_2144), .c(x_in_25_0), .o(n_4830) );
na02f80 g564232 ( .a(n_4862), .b(n_5871), .o(n_5878) );
na03f80 g564233 ( .a(n_5105), .b(n_5743), .c(x_in_51_1), .o(n_5106) );
in01f80 g564234 ( .a(n_6344), .o(n_5653) );
oa12f80 g564235 ( .a(n_3204), .b(n_3203), .c(x_in_37_6), .o(n_6344) );
in01f80 g564236 ( .a(n_6450), .o(n_3857) );
oa12f80 g564237 ( .a(n_3202), .b(n_3201), .c(x_in_37_3), .o(n_6450) );
in01f80 g564238 ( .a(n_4088), .o(n_5717) );
na03f80 g564239 ( .a(n_4863), .b(n_7893), .c(n_3151), .o(n_4088) );
ao12f80 g564240 ( .a(n_2486), .b(n_2143), .c(n_5745), .o(n_10666) );
oa12f80 g564241 ( .a(n_2772), .b(n_2771), .c(x_in_37_15), .o(n_7950) );
in01f80 g564242 ( .a(n_6342), .o(n_3856) );
oa12f80 g564243 ( .a(n_3197), .b(n_3196), .c(x_in_37_4), .o(n_6342) );
in01f80 g564244 ( .a(n_16637), .o(n_5104) );
na02f80 g564245 ( .a(n_5642), .b(n_3252), .o(n_16637) );
ao12f80 g564246 ( .a(n_2557), .b(n_7172), .c(n_2382), .o(n_7947) );
no02f80 g564248 ( .a(n_4016), .b(n_2030), .o(n_13232) );
oa12f80 g564249 ( .a(n_3124), .b(n_3755), .c(x_in_53_0), .o(n_4826) );
in01f80 g564250 ( .a(n_6339), .o(n_5656) );
oa12f80 g564251 ( .a(n_2720), .b(n_2719), .c(x_in_37_7), .o(n_6339) );
no03m80 g564252 ( .a(n_4391), .b(n_4392), .c(x_in_11_3), .o(n_7595) );
no03m80 g564253 ( .a(n_4534), .b(n_4533), .c(x_in_43_3), .o(n_7592) );
in01f80 g564254 ( .a(n_5102), .o(n_5103) );
oa12f80 g564255 ( .a(n_4585), .b(n_5407), .c(n_9329), .o(n_5102) );
ao12f80 g564256 ( .a(n_2738), .b(n_2641), .c(x_in_41_7), .o(n_5686) );
in01f80 g564257 ( .a(n_7429), .o(n_7209) );
oa12f80 g564258 ( .a(n_4573), .b(n_2547), .c(x_in_37_2), .o(n_7429) );
oa12f80 g564259 ( .a(n_3210), .b(n_3209), .c(x_in_61_1), .o(n_6366) );
ao12f80 g564260 ( .a(n_6285), .b(n_4929), .c(n_3853), .o(n_3854) );
no03m80 g564261 ( .a(n_4595), .b(n_4804), .c(x_in_27_3), .o(n_7589) );
ao12f80 g564262 ( .a(n_4029), .b(n_2584), .c(x_in_41_5), .o(n_5635) );
oa12f80 g564263 ( .a(n_3048), .b(n_3818), .c(x_in_47_2), .o(n_5778) );
oa12f80 g564264 ( .a(n_3049), .b(n_3491), .c(x_in_31_2), .o(n_6318) );
in01f80 g564265 ( .a(n_3852), .o(n_5693) );
oa12f80 g564266 ( .a(n_3170), .b(n_4601), .c(n_3186), .o(n_3852) );
oa12f80 g564267 ( .a(n_3185), .b(n_4801), .c(n_4800), .o(n_10085) );
in01f80 g564268 ( .a(n_3851), .o(n_4995) );
oa12f80 g564269 ( .a(n_2669), .b(n_2695), .c(x_in_51_5), .o(n_3851) );
in01f80 g564270 ( .a(n_3850), .o(n_5638) );
oa12f80 g564271 ( .a(n_2647), .b(n_3212), .c(x_in_51_3), .o(n_3850) );
in01f80 g564272 ( .a(n_3484), .o(n_5067) );
oa12f80 g564273 ( .a(n_2682), .b(n_3199), .c(x_in_51_7), .o(n_3484) );
in01f80 g564274 ( .a(n_6335), .o(n_6333) );
oa12f80 g564275 ( .a(n_3342), .b(n_3242), .c(n_4180), .o(n_6335) );
in01f80 g564276 ( .a(n_4039), .o(n_5668) );
oa12f80 g564277 ( .a(n_3315), .b(n_3314), .c(x_in_51_6), .o(n_4039) );
in01f80 g564278 ( .a(n_5101), .o(n_13687) );
no03m80 g564279 ( .a(n_4592), .b(n_4828), .c(n_491), .o(n_5101) );
ao12f80 g564280 ( .a(n_4030), .b(n_2594), .c(x_in_11_14), .o(n_5650) );
ao12f80 g564281 ( .a(x_in_41_15), .b(n_3485), .c(n_9608), .o(n_3071) );
in01f80 g564282 ( .a(n_5626), .o(n_4591) );
ao12f80 g564283 ( .a(n_3848), .b(n_2649), .c(x_in_3_14), .o(n_5626) );
in01f80 g564284 ( .a(n_3892), .o(n_5690) );
oa12f80 g564285 ( .a(n_2357), .b(n_3198), .c(x_in_51_8), .o(n_3892) );
ao12f80 g564286 ( .a(n_3847), .b(n_3811), .c(x_in_51_14), .o(n_6311) );
in01f80 g564287 ( .a(n_5440), .o(n_3846) );
oa12f80 g564288 ( .a(n_3185), .b(n_4800), .c(n_12178), .o(n_5440) );
in01f80 g564289 ( .a(n_10069), .o(n_7593) );
oa12f80 g564290 ( .a(x_in_43_3), .b(n_4533), .c(n_4534), .o(n_10069) );
in01f80 g564291 ( .a(n_10071), .o(n_7596) );
oa12f80 g564292 ( .a(x_in_11_3), .b(n_4392), .c(n_4391), .o(n_10071) );
oa22f80 g564293 ( .a(n_3845), .b(n_2002), .c(n_3736), .d(n_1250), .o(n_8266) );
ao12f80 g564294 ( .a(n_5786), .b(n_2614), .c(x_in_41_10), .o(n_7420) );
in01f80 g564295 ( .a(n_9783), .o(n_10558) );
oa12f80 g564296 ( .a(n_3052), .b(n_5153), .c(x_in_53_11), .o(n_9783) );
oa12f80 g564297 ( .a(n_3384), .b(n_4034), .c(x_in_3_15), .o(n_5622) );
in01f80 g564298 ( .a(n_3842), .o(n_3843) );
oa12f80 g564299 ( .a(n_2696), .b(n_2220), .c(n_5689), .o(n_3842) );
in01f80 g564300 ( .a(n_7430), .o(n_7208) );
oa12f80 g564301 ( .a(n_3202), .b(n_3201), .c(n_3318), .o(n_7430) );
in01f80 g564302 ( .a(n_4588), .o(n_4589) );
ao12f80 g564303 ( .a(n_3642), .b(n_2570), .c(n_3641), .o(n_4588) );
ao12f80 g564304 ( .a(n_6219), .b(n_4448), .c(n_4445), .o(n_4810) );
na03f80 g564305 ( .a(x_in_17_0), .b(n_3689), .c(x_in_17_2), .o(n_10944) );
in01f80 g564306 ( .a(n_10063), .o(n_7590) );
oa12f80 g564307 ( .a(x_in_27_3), .b(n_4804), .c(n_4595), .o(n_10063) );
in01f80 g564308 ( .a(n_6336), .o(n_6337) );
oa12f80 g564309 ( .a(n_3204), .b(n_3203), .c(n_5745), .o(n_6336) );
in01f80 g564310 ( .a(n_6449), .o(n_3840) );
oa12f80 g564311 ( .a(n_3197), .b(n_3196), .c(n_5881), .o(n_6449) );
in01f80 g564312 ( .a(n_5614), .o(n_4587) );
ao12f80 g564313 ( .a(n_4080), .b(n_2324), .c(x_in_27_14), .o(n_5614) );
in01f80 g564314 ( .a(n_5340), .o(n_4586) );
ao12f80 g564315 ( .a(n_3839), .b(n_2338), .c(x_in_43_14), .o(n_5340) );
ao12f80 g564316 ( .a(n_3903), .b(n_3902), .c(x_in_35_14), .o(n_6447) );
in01f80 g564317 ( .a(n_6340), .o(n_5657) );
oa12f80 g564318 ( .a(n_2772), .b(n_2771), .c(n_5962), .o(n_6340) );
ao12f80 g564319 ( .a(n_6209), .b(n_4438), .c(n_4435), .o(n_4584) );
in01f80 g564320 ( .a(n_7435), .o(n_5097) );
na02f80 g564321 ( .a(n_2889), .b(n_2099), .o(n_7435) );
ao12f80 g564322 ( .a(n_6437), .b(n_4434), .c(n_4431), .o(n_4581) );
in01f80 g564323 ( .a(n_6341), .o(n_3369) );
oa12f80 g564324 ( .a(n_2714), .b(n_2713), .c(n_5962), .o(n_6341) );
in01f80 g564325 ( .a(n_6044), .o(n_3375) );
oa12f80 g564326 ( .a(n_2724), .b(n_2723), .c(n_2408), .o(n_6044) );
oa12f80 g564327 ( .a(n_2746), .b(n_2044), .c(n_1), .o(n_6509) );
in01f80 g564328 ( .a(n_6345), .o(n_5654) );
oa12f80 g564329 ( .a(n_2720), .b(n_2719), .c(n_4180), .o(n_6345) );
in01f80 g564330 ( .a(n_6042), .o(n_3836) );
oa22f80 g564331 ( .a(n_3207), .b(n_3237), .c(n_3608), .d(n_5242), .o(n_6042) );
in01f80 g564332 ( .a(n_6357), .o(n_3380) );
oa12f80 g564333 ( .a(n_2733), .b(n_2732), .c(n_4343), .o(n_6357) );
ao12f80 g564334 ( .a(n_2817), .b(n_3242), .c(n_3241), .o(n_3243) );
oa12f80 g564335 ( .a(n_2237), .b(n_2737), .c(n_2691), .o(n_7629) );
in01f80 g564336 ( .a(n_4577), .o(n_4578) );
ao12f80 g564337 ( .a(n_3777), .b(n_2795), .c(x_in_35_0), .o(n_4577) );
no02f80 g564338 ( .a(n_3279), .b(x_in_29_14), .o(n_4167) );
ao12f80 g564339 ( .a(n_5913), .b(n_4423), .c(n_4420), .o(n_4576) );
na03f80 g564340 ( .a(n_6904), .b(n_4574), .c(x_in_33_14), .o(n_4575) );
oa12f80 g564341 ( .a(n_6125), .b(n_4170), .c(n_4165), .o(n_4171) );
in01f80 g564342 ( .a(n_6304), .o(n_7456) );
na02f80 g564343 ( .a(n_2811), .b(n_4573), .o(n_6304) );
ao12f80 g564344 ( .a(n_5713), .b(n_4571), .c(n_4570), .o(n_4572) );
oa12f80 g564345 ( .a(n_2415), .b(n_3498), .c(x_in_35_15), .o(n_5708) );
oa12f80 g564346 ( .a(n_3210), .b(n_3209), .c(n_5242), .o(n_4850) );
oa12f80 g564347 ( .a(n_6769), .b(n_3195), .c(n_4529), .o(n_4848) );
in01f80 g564348 ( .a(n_7453), .o(n_6668) );
na02f80 g564349 ( .a(n_2742), .b(n_4573), .o(n_7453) );
ao12f80 g564350 ( .a(n_2763), .b(n_5153), .c(n_3193), .o(n_3194) );
oa12f80 g564351 ( .a(n_2715), .b(n_2716), .c(x_in_57_13), .o(n_3395) );
ao12f80 g564352 ( .a(n_3834), .b(n_2368), .c(x_in_59_14), .o(n_5624) );
in01f80 g564353 ( .a(n_6288), .o(n_4569) );
ao12f80 g564354 ( .a(n_3398), .b(n_3397), .c(x_in_7_14), .o(n_6288) );
oa22f80 g564355 ( .a(n_2010), .b(n_3833), .c(n_3832), .d(x_in_61_10), .o(n_7891) );
ao12f80 g564356 ( .a(n_2769), .b(n_2768), .c(n_5311), .o(n_2770) );
ao12f80 g564357 ( .a(n_2579), .b(n_3322), .c(x_in_7_6), .o(n_5593) );
ao12f80 g564358 ( .a(n_6172), .b(n_4567), .c(n_4566), .o(n_4568) );
ao12f80 g564359 ( .a(n_6193), .b(n_4260), .c(n_4257), .o(n_4565) );
oa12f80 g564360 ( .a(n_2284), .b(n_3188), .c(n_3191), .o(n_6833) );
ao22s80 g564361 ( .a(n_2225), .b(x_in_49_4), .c(x_in_49_7), .d(x_in_49_6), .o(n_6792) );
oa12f80 g564362 ( .a(n_2204), .b(n_3191), .c(n_3187), .o(n_6867) );
ao22s80 g564363 ( .a(n_2218), .b(x_in_49_5), .c(x_in_49_8), .d(x_in_49_7), .o(n_6860) );
ao12f80 g564364 ( .a(n_5763), .b(n_4428), .c(n_4426), .o(n_4564) );
ao22s80 g564365 ( .a(n_2216), .b(x_in_49_3), .c(x_in_49_6), .d(x_in_49_5), .o(n_6831) );
ao12f80 g564366 ( .a(FE_OFN991_n_5720), .b(n_4513), .c(n_4511), .o(n_4563) );
oa12f80 g564367 ( .a(n_4562), .b(n_3238), .c(x_in_49_1), .o(n_7877) );
ao12f80 g564368 ( .a(n_5850), .b(n_2393), .c(x_in_3_4), .o(n_4561) );
ao22s80 g564369 ( .a(n_2249), .b(x_in_49_9), .c(x_in_49_12), .d(x_in_49_11), .o(n_6835) );
ao12f80 g564370 ( .a(n_6098), .b(n_4463), .c(n_4460), .o(n_4560) );
ao12f80 g564371 ( .a(n_6175), .b(n_4452), .c(n_4449), .o(n_4559) );
ao12f80 g564372 ( .a(n_2211), .b(n_2768), .c(n_3189), .o(n_3190) );
no02f80 g564373 ( .a(n_3269), .b(n_6049), .o(n_4558) );
no02f80 g564374 ( .a(n_2792), .b(n_6184), .o(n_4557) );
ao12f80 g564375 ( .a(n_6055), .b(n_4494), .c(n_4491), .o(n_4556) );
oa22f80 g564376 ( .a(n_2011), .b(n_5761), .c(n_4923), .d(x_in_61_6), .o(n_7889) );
in01f80 g564377 ( .a(n_8596), .o(n_6441) );
oa22f80 g564378 ( .a(n_2012), .b(n_5242), .c(n_6731), .d(x_in_61_5), .o(n_8596) );
oa22f80 g564379 ( .a(n_2021), .b(n_3188), .c(n_3187), .d(n_3186), .o(n_7632) );
ao12f80 g564380 ( .a(n_2820), .b(n_2493), .c(x_in_25_12), .o(n_6414) );
oa12f80 g564381 ( .a(x_in_57_4), .b(n_2219), .c(n_4668), .o(n_10095) );
in01f80 g564382 ( .a(n_4553), .o(n_8876) );
oa22f80 g564383 ( .a(n_1985), .b(n_8929), .c(n_3447), .d(x_in_61_4), .o(n_4553) );
ao12f80 g564384 ( .a(n_6164), .b(n_4240), .c(n_4239), .o(n_4241) );
ao12f80 g564385 ( .a(n_4710), .b(n_3809), .c(n_5281), .o(n_4552) );
in01f80 g564386 ( .a(n_8469), .o(n_4551) );
oa22f80 g564387 ( .a(n_2027), .b(n_4914), .c(n_4651), .d(x_in_61_9), .o(n_8469) );
in01f80 g564388 ( .a(n_8516), .o(n_4256) );
oa22f80 g564389 ( .a(n_2020), .b(n_5839), .c(n_7445), .d(x_in_61_7), .o(n_8516) );
ao12f80 g564390 ( .a(n_2832), .b(n_2113), .c(n_23944), .o(n_2833) );
in01f80 g564391 ( .a(n_6352), .o(n_3826) );
oa12f80 g564392 ( .a(n_2798), .b(n_5820), .c(n_12175), .o(n_6352) );
in01f80 g564393 ( .a(n_8075), .o(n_4550) );
oa22f80 g564394 ( .a(n_2005), .b(n_4937), .c(n_4397), .d(x_in_61_8), .o(n_8075) );
oa12f80 g564395 ( .a(n_5450), .b(n_3762), .c(x_in_23_2), .o(n_3823) );
ao12f80 g564396 ( .a(n_3822), .b(n_3716), .c(x_in_61_14), .o(n_5769) );
oa12f80 g564397 ( .a(n_3821), .b(n_3820), .c(x_in_57_12), .o(n_5428) );
ao12f80 g564398 ( .a(n_3526), .b(n_3233), .c(x_in_35_3), .o(n_5606) );
oa12f80 g564399 ( .a(n_11226), .b(n_2676), .c(n_5245), .o(n_8499) );
ao12f80 g564400 ( .a(n_5777), .b(n_3818), .c(n_5365), .o(n_3819) );
ao12f80 g564401 ( .a(n_6317), .b(n_3491), .c(n_5373), .o(n_3492) );
ao12f80 g564402 ( .a(n_3055), .b(n_3634), .c(x_in_27_1), .o(n_6299) );
in01f80 g564403 ( .a(n_6381), .o(n_3817) );
oa12f80 g564404 ( .a(n_3052), .b(n_5153), .c(n_2870), .o(n_6381) );
in01f80 g564405 ( .a(n_6343), .o(n_3816) );
oa12f80 g564406 ( .a(n_2877), .b(n_4203), .c(n_8885), .o(n_6343) );
in01f80 g564407 ( .a(n_6348), .o(n_4054) );
oa12f80 g564408 ( .a(n_2879), .b(n_5228), .c(n_12178), .o(n_6348) );
in01f80 g564409 ( .a(n_6346), .o(n_3813) );
oa12f80 g564410 ( .a(n_3072), .b(n_4692), .c(n_8884), .o(n_6346) );
in01f80 g564411 ( .a(n_6347), .o(n_3519) );
oa12f80 g564412 ( .a(n_3070), .b(n_5231), .c(n_12634), .o(n_6347) );
in01f80 g564413 ( .a(n_5094), .o(n_7217) );
oa12f80 g564414 ( .a(n_3324), .b(n_2659), .c(x_in_45_15), .o(n_5094) );
in01f80 g564415 ( .a(n_5597), .o(n_6730) );
ao12f80 g564416 ( .a(n_2384), .b(n_2906), .c(x_in_61_6), .o(n_5597) );
in01f80 g564417 ( .a(n_6349), .o(n_3812) );
oa12f80 g564418 ( .a(n_2805), .b(n_5224), .c(n_12635), .o(n_6349) );
in01f80 g564419 ( .a(n_5093), .o(n_7478) );
oa12f80 g564420 ( .a(n_3980), .b(n_21777), .c(x_in_25_12), .o(n_5093) );
ao12f80 g564421 ( .a(n_4970), .b(n_4410), .c(x_in_59_15), .o(n_6278) );
ao12f80 g564422 ( .a(n_3847), .b(n_3811), .c(n_8420), .o(n_5601) );
in01f80 g564423 ( .a(n_4546), .o(n_6272) );
oa12f80 g564424 ( .a(n_3054), .b(n_3634), .c(n_5677), .o(n_4546) );
in01f80 g564425 ( .a(n_4544), .o(n_4545) );
ao12f80 g564426 ( .a(n_3239), .b(n_3838), .c(n_4325), .o(n_4544) );
oa12f80 g564427 ( .a(n_6475), .b(n_5046), .c(x_in_29_10), .o(n_9540) );
ao12f80 g564428 ( .a(n_3543), .b(n_2827), .c(x_in_35_9), .o(n_5437) );
ao22s80 g564429 ( .a(n_2244), .b(n_5387), .c(x_in_11_7), .d(x_in_11_5), .o(n_5660) );
in01f80 g564430 ( .a(n_4844), .o(n_6354) );
oa22f80 g564431 ( .a(n_2032), .b(x_in_7_4), .c(n_5256), .d(n_6494), .o(n_4844) );
in01f80 g564432 ( .a(n_4543), .o(n_7201) );
ao12f80 g564433 ( .a(n_4401), .b(n_3809), .c(x_in_33_6), .o(n_4543) );
in01f80 g564434 ( .a(n_3808), .o(n_5514) );
oa22f80 g564435 ( .a(n_1978), .b(x_in_11_9), .c(n_3229), .d(n_5025), .o(n_3808) );
ao12f80 g564436 ( .a(n_5943), .b(n_2464), .c(n_2310), .o(n_4542) );
oa12f80 g564437 ( .a(n_5639), .b(n_2280), .c(x_in_41_4), .o(n_4366) );
ao12f80 g564438 ( .a(n_5832), .b(n_4035), .c(x_in_35_4), .o(n_4541) );
ao12f80 g564439 ( .a(n_2551), .b(x_in_11_8), .c(x_in_11_6), .o(n_5661) );
ao12f80 g564440 ( .a(n_3051), .b(n_4540), .c(x_in_17_14), .o(n_6231) );
oa12f80 g564441 ( .a(n_5752), .b(n_2473), .c(x_in_21_12), .o(n_4539) );
ao12f80 g564442 ( .a(n_2405), .b(n_3330), .c(x_in_21_9), .o(n_6011) );
no03m80 g564443 ( .a(n_3803), .b(n_5772), .c(x_in_45_1), .o(n_3807) );
oa12f80 g564444 ( .a(n_5855), .b(n_2107), .c(x_in_45_2), .o(n_4538) );
oa12f80 g564445 ( .a(n_3806), .b(n_3388), .c(x_in_11_10), .o(n_9977) );
in01f80 g564446 ( .a(n_3805), .o(n_5301) );
oa22f80 g564447 ( .a(n_2008), .b(x_in_11_6), .c(n_5089), .d(n_5310), .o(n_3805) );
ao22s80 g564448 ( .a(n_2274), .b(n_5089), .c(x_in_11_10), .d(x_in_11_8), .o(n_5561) );
oa12f80 g564449 ( .a(x_in_45_1), .b(n_5772), .c(n_3803), .o(n_3804) );
in01f80 g564450 ( .a(n_4387), .o(n_5741) );
ao12f80 g564451 ( .a(n_3386), .b(n_3090), .c(x_in_35_10), .o(n_4387) );
in01f80 g564452 ( .a(n_6747), .o(n_4537) );
ao12f80 g564453 ( .a(n_2485), .b(n_3333), .c(x_in_7_9), .o(n_6747) );
in01f80 g564454 ( .a(n_6308), .o(n_7559) );
ao12f80 g564455 ( .a(n_2844), .b(n_2307), .c(x_in_7_11), .o(n_6308) );
oa12f80 g564456 ( .a(n_3655), .b(n_3298), .c(x_in_61_10), .o(n_9972) );
in01f80 g564457 ( .a(n_6770), .o(n_5092) );
ao12f80 g564458 ( .a(n_3081), .b(n_2622), .c(x_in_61_12), .o(n_6770) );
in01f80 g564459 ( .a(n_3750), .o(n_5525) );
oa22f80 g564460 ( .a(n_1999), .b(x_in_3_4), .c(n_5963), .d(n_5757), .o(n_3750) );
oa12f80 g564461 ( .a(n_6230), .b(n_2087), .c(x_in_17_12), .o(n_3754) );
in01f80 g564462 ( .a(n_4536), .o(n_5746) );
ao12f80 g564463 ( .a(n_2347), .b(n_3875), .c(x_in_59_12), .o(n_4536) );
ao12f80 g564464 ( .a(n_3782), .b(n_3222), .c(x_in_35_4), .o(n_5587) );
in01f80 g564465 ( .a(n_5091), .o(n_6654) );
ao12f80 g564466 ( .a(n_2848), .b(n_2482), .c(x_in_7_10), .o(n_5091) );
in01f80 g564467 ( .a(n_6722), .o(n_4535) );
ao12f80 g564468 ( .a(n_2675), .b(n_3083), .c(x_in_61_9), .o(n_6722) );
ao12f80 g564469 ( .a(n_2396), .b(n_3691), .c(x_in_59_8), .o(n_5585) );
in01f80 g564470 ( .a(n_3802), .o(n_5492) );
oa22f80 g564471 ( .a(n_1998), .b(x_in_43_9), .c(n_6496), .d(n_7263), .o(n_3802) );
in01f80 g564472 ( .a(n_3837), .o(n_5683) );
oa22f80 g564473 ( .a(n_1986), .b(x_in_27_9), .c(n_7417), .d(n_7402), .o(n_3837) );
oa12f80 g564474 ( .a(n_5749), .b(n_2689), .c(x_in_37_9), .o(n_4590) );
ao22s80 g564475 ( .a(n_2048), .b(n_5963), .c(x_in_3_8), .d(x_in_3_6), .o(n_5667) );
in01f80 g564476 ( .a(n_6785), .o(n_5090) );
ao12f80 g564477 ( .a(n_2728), .b(n_2381), .c(x_in_7_12), .o(n_6785) );
in01f80 g564478 ( .a(n_3801), .o(n_5065) );
oa22f80 g564479 ( .a(n_1976), .b(x_in_27_5), .c(n_5677), .d(n_7287), .o(n_3801) );
oa12f80 g564480 ( .a(n_5882), .b(n_3040), .c(x_in_37_10), .o(n_4750) );
oa12f80 g564481 ( .a(n_5087), .b(n_2477), .c(x_in_21_11), .o(n_5088) );
in01f80 g564482 ( .a(n_4879), .o(n_3800) );
oa22f80 g564483 ( .a(n_1982), .b(x_in_3_6), .c(n_5757), .d(n_5905), .o(n_4879) );
ao22s80 g564484 ( .a(n_2047), .b(n_5757), .c(x_in_3_10), .d(x_in_3_8), .o(n_5675) );
in01f80 g564485 ( .a(n_7540), .o(n_5085) );
ao12f80 g564486 ( .a(n_3334), .b(n_2371), .c(x_in_21_7), .o(n_7540) );
ao12f80 g564487 ( .a(n_2665), .b(n_3368), .c(x_in_59_10), .o(n_5581) );
in01f80 g564488 ( .a(n_4158), .o(n_6402) );
oa12f80 g564489 ( .a(n_2340), .b(n_3366), .c(n_4942), .o(n_4158) );
ao22s80 g564490 ( .a(n_2208), .b(n_5352), .c(x_in_11_11), .d(x_in_11_9), .o(n_5569) );
in01f80 g564491 ( .a(n_3799), .o(n_5041) );
oa22f80 g564492 ( .a(n_1991), .b(x_in_3_9), .c(n_5666), .d(n_5247), .o(n_3799) );
in01f80 g564493 ( .a(n_3798), .o(n_5494) );
oa22f80 g564494 ( .a(n_2019), .b(x_in_43_6), .c(n_5519), .d(n_7268), .o(n_3798) );
in01f80 g564495 ( .a(n_5496), .o(n_4796) );
ao12f80 g564496 ( .a(n_3632), .b(n_2466), .c(x_in_59_9), .o(n_5496) );
in01f80 g564497 ( .a(n_6768), .o(n_5084) );
ao12f80 g564498 ( .a(n_3332), .b(n_2458), .c(x_in_61_10), .o(n_6768) );
in01f80 g564499 ( .a(n_3795), .o(n_5152) );
oa22f80 g564500 ( .a(n_1996), .b(x_in_27_4), .c(n_3747), .d(n_5680), .o(n_3795) );
oa12f80 g564501 ( .a(n_2475), .b(n_3082), .c(x_in_19_10), .o(n_9937) );
ao12f80 g564502 ( .a(n_5880), .b(n_2303), .c(n_5881), .o(n_4799) );
oa12f80 g564503 ( .a(n_4739), .b(n_2465), .c(x_in_57_11), .o(n_4175) );
oa12f80 g564505 ( .a(n_2613), .b(n_4122), .c(x_in_59_10), .o(n_9929) );
in01f80 g564506 ( .a(n_6358), .o(n_6356) );
oa22f80 g564507 ( .a(n_2031), .b(x_in_37_8), .c(n_4180), .d(n_5962), .o(n_6358) );
oa12f80 g564508 ( .a(n_3650), .b(n_3438), .c(x_in_43_10), .o(n_9943) );
in01f80 g564509 ( .a(n_3791), .o(n_5100) );
oa22f80 g564510 ( .a(n_2018), .b(x_in_27_7), .c(n_7287), .d(n_7417), .o(n_3791) );
ao12f80 g564511 ( .a(n_3353), .b(n_3257), .c(x_in_35_6), .o(n_5663) );
ao12f80 g564512 ( .a(n_3449), .b(n_3255), .c(x_in_35_8), .o(n_5576) );
ao12f80 g564513 ( .a(n_3453), .b(n_2468), .c(x_in_51_5), .o(n_5574) );
in01f80 g564514 ( .a(n_4156), .o(n_6733) );
ao12f80 g564515 ( .a(n_4063), .b(n_4062), .c(n_5977), .o(n_4156) );
ao22s80 g564516 ( .a(n_2062), .b(n_5156), .c(x_in_35_4), .d(x_in_35_2), .o(n_5659) );
in01f80 g564517 ( .a(n_4530), .o(n_6474) );
oa12f80 g564518 ( .a(n_2407), .b(n_3313), .c(n_5869), .o(n_4530) );
in01f80 g564519 ( .a(n_5579), .o(n_4215) );
ao12f80 g564520 ( .a(n_3903), .b(n_3902), .c(n_8524), .o(n_5579) );
ao12f80 g564521 ( .a(n_3248), .b(n_2298), .c(x_in_21_6), .o(n_6282) );
ao12f80 g564522 ( .a(n_5751), .b(n_8010), .c(n_5872), .o(n_4597) );
ao12f80 g564523 ( .a(n_2432), .b(x_in_11_5), .c(x_in_11_3), .o(n_5549) );
in01f80 g564524 ( .a(n_4072), .o(n_5445) );
oa22f80 g564525 ( .a(n_1990), .b(x_in_43_7), .c(n_5501), .d(n_6496), .o(n_4072) );
in01f80 g564526 ( .a(n_4083), .o(n_5493) );
oa22f80 g564527 ( .a(n_2024), .b(x_in_27_6), .c(n_5680), .d(n_7289), .o(n_4083) );
ao12f80 g564528 ( .a(n_5922), .b(n_7715), .c(n_3036), .o(n_4791) );
ao12f80 g564529 ( .a(n_2577), .b(n_3084), .c(x_in_21_8), .o(n_5589) );
oa12f80 g564530 ( .a(n_3789), .b(n_2868), .c(x_in_7_10), .o(n_9910) );
ao22s80 g564531 ( .a(n_2094), .b(n_5825), .c(x_in_3_6), .d(x_in_3_4), .o(n_5528) );
oa12f80 g564532 ( .a(n_3788), .b(n_3501), .c(x_in_27_10), .o(n_9907) );
ao12f80 g564533 ( .a(n_2553), .b(x_in_27_4), .c(x_in_27_2), .o(n_5678) );
ao12f80 g564534 ( .a(n_3220), .b(n_2337), .c(x_in_7_8), .o(n_6276) );
in01f80 g564535 ( .a(n_3787), .o(n_5509) );
oa22f80 g564536 ( .a(n_1989), .b(x_in_43_5), .c(n_5327), .d(n_5501), .o(n_3787) );
ao12f80 g564537 ( .a(n_2412), .b(x_in_43_5), .c(x_in_43_3), .o(n_5520) );
ao12f80 g564538 ( .a(n_5822), .b(n_3104), .c(x_in_19_4), .o(n_4806) );
ao12f80 g564539 ( .a(n_3629), .b(n_2559), .c(x_in_3_4), .o(n_5516) );
in01f80 g564540 ( .a(n_4058), .o(n_5548) );
oa22f80 g564541 ( .a(n_1993), .b(x_in_43_8), .c(n_7268), .d(n_8443), .o(n_4058) );
in01f80 g564542 ( .a(n_3583), .o(n_5502) );
oa22f80 g564543 ( .a(n_2006), .b(x_in_27_8), .c(n_7289), .d(n_8513), .o(n_3583) );
in01f80 g564544 ( .a(n_5081), .o(n_7555) );
oa12f80 g564545 ( .a(n_3078), .b(n_2450), .c(n_4529), .o(n_5081) );
in01f80 g564546 ( .a(n_6364), .o(n_3786) );
na02f80 g564547 ( .a(n_2199), .b(n_2001), .o(n_6364) );
in01f80 g564548 ( .a(n_5734), .o(n_4973) );
oa12f80 g564549 ( .a(n_3223), .b(n_2313), .c(n_5900), .o(n_5734) );
ao12f80 g564550 ( .a(n_2804), .b(n_2639), .c(x_in_61_8), .o(n_6223) );
ao12f80 g564551 ( .a(n_3358), .b(n_2591), .c(x_in_59_11), .o(n_5583) );
in01f80 g564552 ( .a(n_5500), .o(n_4893) );
oa12f80 g564553 ( .a(n_2345), .b(n_3448), .c(n_5519), .o(n_5500) );
na03f80 g564554 ( .a(n_2529), .b(n_4403), .c(n_4138), .o(n_5433) );
in01f80 g564555 ( .a(n_3785), .o(n_5096) );
oa22f80 g564556 ( .a(n_2015), .b(x_in_3_8), .c(n_5905), .d(n_6380), .o(n_3785) );
ao12f80 g564558 ( .a(n_2435), .b(x_in_11_6), .c(x_in_11_4), .o(n_5546) );
in01f80 g564559 ( .a(n_4527), .o(n_6739) );
oa12f80 g564560 ( .a(n_3235), .b(n_3362), .c(x_in_53_12), .o(n_4527) );
ao12f80 g564561 ( .a(n_3331), .b(n_2456), .c(x_in_51_7), .o(n_6429) );
ao12f80 g564562 ( .a(n_2359), .b(n_3784), .c(x_in_35_5), .o(n_5565) );
oa12f80 g564563 ( .a(n_2661), .b(n_3379), .c(x_in_35_10), .o(n_9883) );
in01f80 g564564 ( .a(n_4935), .o(n_7442) );
oa12f80 g564565 ( .a(n_2901), .b(n_2356), .c(n_5839), .o(n_4935) );
in01f80 g564566 ( .a(n_3783), .o(n_5530) );
oa22f80 g564567 ( .a(n_1987), .b(x_in_3_2), .c(n_5825), .d(n_5963), .o(n_3783) );
ao12f80 g564568 ( .a(n_2333), .b(x_in_11_4), .c(x_in_11_2), .o(n_5551) );
in01f80 g564569 ( .a(n_5080), .o(n_7479) );
oa12f80 g564570 ( .a(n_2888), .b(n_2461), .c(n_8557), .o(n_5080) );
oa12f80 g564571 ( .a(n_2873), .b(n_2377), .c(n_5987), .o(n_11157) );
ao12f80 g564572 ( .a(n_4034), .b(n_3384), .c(n_5666), .o(n_9875) );
ao12f80 g564573 ( .a(n_2552), .b(x_in_43_4), .c(x_in_43_2), .o(n_5498) );
oa12f80 g564574 ( .a(n_3599), .b(n_3591), .c(x_in_29_1), .o(n_8316) );
ao12f80 g564575 ( .a(n_3385), .b(n_2496), .c(n_5283), .o(n_9878) );
ao12f80 g564576 ( .a(n_2402), .b(x_in_27_5), .c(x_in_27_3), .o(n_5681) );
in01f80 g564577 ( .a(n_5572), .o(n_6717) );
no02f80 g564578 ( .a(n_2502), .b(n_2206), .o(n_5572) );
ao12f80 g564579 ( .a(n_3822), .b(n_3716), .c(n_4529), .o(n_5784) );
ao12f80 g564580 ( .a(n_2489), .b(x_in_43_6), .c(x_in_43_4), .o(n_5505) );
in01f80 g564581 ( .a(n_6385), .o(n_4912) );
oa22f80 g564582 ( .a(n_2000), .b(x_in_7_1), .c(n_8522), .d(n_2699), .o(n_6385) );
ao12f80 g564583 ( .a(n_3108), .b(n_3781), .c(n_3753), .o(n_10804) );
ao12f80 g564584 ( .a(n_2446), .b(x_in_59_4), .c(x_in_59_2), .o(n_5532) );
in01f80 g564585 ( .a(n_6391), .o(n_4190) );
ao22s80 g564586 ( .a(n_2056), .b(n_5849), .c(n_3241), .d(x_in_37_14), .o(n_6391) );
oa12f80 g564587 ( .a(n_3047), .b(n_3781), .c(n_5938), .o(n_10812) );
ao12f80 g564588 ( .a(n_7211), .b(n_4970), .c(n_8336), .o(n_4971) );
in01f80 g564589 ( .a(n_8925), .o(n_5079) );
oa12f80 g564590 ( .a(n_4197), .b(n_4196), .c(x_in_61_3), .o(n_8925) );
in01f80 g564591 ( .a(n_9091), .o(n_5783) );
ao12f80 g564592 ( .a(n_6884), .b(n_4972), .c(n_8851), .o(n_9091) );
in01f80 g564593 ( .a(n_4525), .o(n_4526) );
ao12f80 g564594 ( .a(n_3034), .b(n_4664), .c(n_3415), .o(n_4525) );
oa12f80 g564595 ( .a(n_3026), .b(n_4664), .c(n_3780), .o(n_10781) );
in01f80 g564596 ( .a(n_7557), .o(n_5078) );
ao22s80 g564597 ( .a(n_2690), .b(x_in_3_13), .c(n_3321), .d(n_6746), .o(n_7557) );
oa22f80 g564598 ( .a(n_4524), .b(n_3122), .c(n_4523), .d(n_4522), .o(n_6120) );
ao22s80 g564599 ( .a(n_2259), .b(n_5293), .c(n_3178), .d(x_in_43_4), .o(n_5670) );
ao22s80 g564600 ( .a(n_2765), .b(n_5271), .c(n_2051), .d(x_in_59_4), .o(n_5672) );
ao22s80 g564601 ( .a(n_4218), .b(n_3431), .c(n_3432), .d(n_4217), .o(n_6108) );
ao22s80 g564602 ( .a(n_4521), .b(n_4093), .c(n_4094), .d(n_4520), .o(n_6191) );
in01f80 g564603 ( .a(n_6395), .o(n_4519) );
ao22s80 g564604 ( .a(n_2281), .b(x_in_55_11), .c(n_5376), .d(x_in_55_12), .o(n_6395) );
ao22s80 g564605 ( .a(n_8058), .b(n_3694), .c(n_3695), .d(n_4518), .o(n_6864) );
oa22f80 g564606 ( .a(n_3178), .b(n_3177), .c(n_5293), .d(n_3176), .o(n_11683) );
in01f80 g564607 ( .a(n_6393), .o(n_4874) );
ao22s80 g564608 ( .a(n_2212), .b(x_in_63_11), .c(n_5042), .d(x_in_63_12), .o(n_6393) );
ao12f80 g564609 ( .a(n_2351), .b(x_in_11_5), .c(x_in_11_4), .o(n_11115) );
oa22f80 g564610 ( .a(n_3485), .b(x_in_41_12), .c(n_2151), .d(n_9608), .o(n_5563) );
oa22f80 g564611 ( .a(n_2679), .b(n_4516), .c(n_4515), .d(n_2245), .o(n_6185) );
in01f80 g564612 ( .a(n_6772), .o(n_4988) );
oa22f80 g564613 ( .a(n_2685), .b(x_in_39_11), .c(n_2809), .d(n_7317), .o(n_6772) );
in01f80 g564614 ( .a(n_7467), .o(n_4994) );
ao22s80 g564615 ( .a(n_2767), .b(n_4514), .c(n_2582), .d(x_in_39_9), .o(n_7467) );
oa22f80 g564616 ( .a(n_4260), .b(n_4259), .c(n_4258), .d(n_4257), .o(n_6194) );
ao22s80 g564617 ( .a(n_2239), .b(n_5387), .c(n_2350), .d(x_in_11_4), .o(n_5542) );
ao22s80 g564618 ( .a(n_3777), .b(n_5987), .c(n_2794), .d(x_in_35_4), .o(n_5507) );
oa22f80 g564619 ( .a(n_3776), .b(x_in_17_8), .c(n_2084), .d(n_5360), .o(n_5461) );
in01f80 g564620 ( .a(n_7448), .o(n_5001) );
ao22s80 g564621 ( .a(n_2750), .b(n_8851), .c(n_2677), .d(x_in_39_10), .o(n_7448) );
oa22f80 g564622 ( .a(n_4346), .b(n_3273), .c(n_3274), .d(n_4345), .o(n_6217) );
ao12f80 g564623 ( .a(n_4077), .b(n_4076), .c(x_in_39_4), .o(n_5022) );
ao22s80 g564624 ( .a(n_4065), .b(n_5336), .c(n_2565), .d(x_in_55_2), .o(n_4906) );
oa22f80 g564625 ( .a(n_4310), .b(n_3300), .c(n_3301), .d(n_4309), .o(n_6170) );
ao22s80 g564626 ( .a(n_4068), .b(n_4687), .c(n_2837), .d(x_in_17_2), .o(n_5454) );
in01f80 g564627 ( .a(n_6780), .o(n_5665) );
ao22s80 g564628 ( .a(n_3346), .b(n_4338), .c(n_2344), .d(x_in_39_5), .o(n_6780) );
ao22s80 g564629 ( .a(n_2315), .b(x_in_61_1), .c(n_2998), .d(n_3237), .o(n_10765) );
ao12f80 g564630 ( .a(n_3033), .b(n_3849), .c(n_3780), .o(n_10737) );
ao22s80 g564631 ( .a(n_3177), .b(x_in_43_6), .c(n_2092), .d(n_5327), .o(n_3772) );
oa22f80 g564632 ( .a(n_4513), .b(n_4512), .c(n_6022), .d(n_4511), .o(n_5721) );
oa22f80 g564633 ( .a(n_4509), .b(n_3306), .c(n_3307), .d(n_4508), .o(n_6182) );
oa22f80 g564634 ( .a(n_4507), .b(n_2838), .c(n_2839), .d(n_4506), .o(n_6143) );
na03f80 g564635 ( .a(n_4763), .b(n_2586), .c(n_4870), .o(n_11449) );
in01f80 g564636 ( .a(n_6397), .o(n_4505) );
ao22s80 g564637 ( .a(n_2100), .b(x_in_15_11), .c(n_5368), .d(x_in_15_12), .o(n_6397) );
in01f80 g564638 ( .a(n_5517), .o(n_4873) );
oa22f80 g564639 ( .a(n_2556), .b(x_in_25_6), .c(n_2080), .d(n_3771), .o(n_5517) );
oa22f80 g564640 ( .a(n_4504), .b(n_3140), .c(n_3141), .d(n_4503), .o(n_6062) );
oa22f80 g564641 ( .a(n_4370), .b(n_4129), .c(n_4130), .d(n_4369), .o(n_6167) );
oa22f80 g564642 ( .a(n_2302), .b(n_4374), .c(n_4373), .d(n_2275), .o(n_6050) );
oa22f80 g564643 ( .a(n_4240), .b(n_4502), .c(n_6013), .d(n_4239), .o(n_6165) );
oa22f80 g564644 ( .a(n_4390), .b(n_3110), .c(n_4389), .d(n_4388), .o(n_6162) );
oa22f80 g564645 ( .a(n_4501), .b(n_3327), .c(n_3328), .d(n_4500), .o(n_6179) );
ao22s80 g564646 ( .a(n_8071), .b(n_4102), .c(n_4103), .d(n_4405), .o(n_6858) );
oa22f80 g564647 ( .a(n_4499), .b(n_2693), .c(n_4498), .d(n_4497), .o(n_6096) );
oa22f80 g564648 ( .a(n_4532), .b(n_3294), .c(n_3295), .d(n_4531), .o(n_6158) );
oa22f80 g564649 ( .a(n_4496), .b(n_4134), .c(n_4135), .d(n_4495), .o(n_6155) );
oa22f80 g564650 ( .a(n_4494), .b(n_4493), .c(n_4492), .d(n_4491), .o(n_6056) );
oa22f80 g564651 ( .a(n_4549), .b(n_2866), .c(n_4548), .d(n_4547), .o(n_6152) );
ao22s80 g564652 ( .a(n_4490), .b(n_3459), .c(n_3460), .d(n_4489), .o(n_6149) );
oa22f80 g564653 ( .a(n_4567), .b(n_4583), .c(n_4582), .d(n_4566), .o(n_6173) );
oa22f80 g564654 ( .a(n_4488), .b(n_3281), .c(n_3282), .d(n_4487), .o(n_6146) );
ao22s80 g564655 ( .a(n_8069), .b(n_4115), .c(n_4116), .d(n_4596), .o(n_6852) );
ao22s80 g564656 ( .a(n_3417), .b(n_5931), .c(n_3234), .d(x_in_3_4), .o(n_5510) );
in01f80 g564657 ( .a(n_6396), .o(n_4667) );
ao22s80 g564658 ( .a(n_2133), .b(x_in_47_11), .c(n_5363), .d(x_in_47_12), .o(n_6396) );
oa22f80 g564659 ( .a(n_3770), .b(x_in_17_11), .c(n_2091), .d(n_5418), .o(n_5490) );
oa22f80 g564660 ( .a(n_4022), .b(x_in_17_4), .c(n_2064), .d(n_4021), .o(n_5469) );
in01f80 g564661 ( .a(n_9855), .o(n_5238) );
ao22s80 g564662 ( .a(n_2620), .b(x_in_17_14), .c(n_2751), .d(n_4794), .o(n_9855) );
in01f80 g564663 ( .a(n_6789), .o(n_5073) );
oa12f80 g564664 ( .a(n_3097), .b(n_3096), .c(x_in_29_4), .o(n_6789) );
ao22s80 g564665 ( .a(n_5048), .b(n_2121), .c(n_3363), .d(x_in_17_3), .o(n_6849) );
oa22f80 g564666 ( .a(n_4571), .b(n_4798), .c(n_4797), .d(n_4570), .o(n_5714) );
oa12f80 g564667 ( .a(n_3125), .b(n_3481), .c(n_4486), .o(n_6027) );
in01f80 g564668 ( .a(n_7518), .o(n_5072) );
ao22s80 g564669 ( .a(n_4540), .b(x_in_17_13), .c(n_3638), .d(n_10477), .o(n_7518) );
oa22f80 g564670 ( .a(n_4929), .b(n_4890), .c(n_4928), .d(n_3853), .o(n_6286) );
oa22f80 g564671 ( .a(n_4885), .b(n_2815), .c(n_4884), .d(n_4883), .o(n_6134) );
oa22f80 g564672 ( .a(n_4485), .b(n_3114), .c(n_3115), .d(n_4484), .o(n_6090) );
ao22s80 g564673 ( .a(n_4483), .b(n_4059), .c(n_4060), .d(n_4482), .o(n_6214) );
ao22s80 g564674 ( .a(n_6372), .b(n_3692), .c(n_4481), .d(n_4480), .o(n_6131) );
in01f80 g564675 ( .a(n_3767), .o(n_11150) );
oa22f80 g564676 ( .a(n_3175), .b(n_2009), .c(n_3174), .d(n_5939), .o(n_3767) );
ao22s80 g564677 ( .a(n_2068), .b(n_5939), .c(n_3175), .d(x_in_19_4), .o(n_5521) );
oa12f80 g564678 ( .a(n_3145), .b(n_3144), .c(n_4479), .o(n_6073) );
in01f80 g564679 ( .a(n_6394), .o(n_4478) );
ao22s80 g564680 ( .a(n_2063), .b(x_in_31_11), .c(n_5355), .d(x_in_31_12), .o(n_6394) );
in01f80 g564681 ( .a(n_6398), .o(n_4477) );
ao22s80 g564682 ( .a(n_2059), .b(x_in_23_11), .c(n_5371), .d(x_in_23_12), .o(n_6398) );
ao22s80 g564683 ( .a(n_5265), .b(n_3511), .c(n_4476), .d(n_4475), .o(n_6059) );
oa22f80 g564684 ( .a(n_4474), .b(n_3686), .c(n_3687), .d(n_4473), .o(n_6123) );
oa22f80 g564685 ( .a(n_4472), .b(n_2759), .c(n_2760), .d(n_4471), .o(n_6117) );
oa22f80 g564686 ( .a(n_4470), .b(n_2881), .c(n_4469), .d(n_4468), .o(n_6114) );
oa22f80 g564687 ( .a(n_4467), .b(n_3338), .c(n_3339), .d(n_4466), .o(n_6111) );
oa22f80 g564688 ( .a(n_4465), .b(n_3284), .c(n_3285), .d(n_4464), .o(n_6102) );
oa22f80 g564689 ( .a(n_4463), .b(n_4462), .c(n_4461), .d(n_4460), .o(n_6099) );
ao22s80 g564690 ( .a(n_3764), .b(n_5351), .c(n_2571), .d(x_in_63_2), .o(n_5448) );
oa22f80 g564691 ( .a(n_4459), .b(n_3467), .c(n_3468), .d(n_4458), .o(n_6445) );
oa12f80 g564692 ( .a(n_3147), .b(n_3287), .c(n_4457), .o(n_6439) );
ao22s80 g564693 ( .a(n_5074), .b(n_2123), .c(n_3763), .d(x_in_19_3), .o(n_6837) );
ao22s80 g564694 ( .a(n_3762), .b(n_5430), .c(n_3761), .d(x_in_23_2), .o(n_5451) );
ao22s80 g564695 ( .a(n_2038), .b(n_9646), .c(n_3760), .d(x_in_17_5), .o(n_5479) );
oa12f80 g564696 ( .a(n_3064), .b(n_5979), .c(n_3792), .o(n_10194) );
oa12f80 g564697 ( .a(n_2531), .b(n_2628), .c(x_in_1_2), .o(n_4949) );
ao22s80 g564698 ( .a(n_2364), .b(x_in_7_4), .c(n_2260), .d(n_8522), .o(n_3759) );
ao22s80 g564699 ( .a(n_5263), .b(n_2705), .c(n_5264), .d(n_4456), .o(n_6137) );
ao22s80 g564700 ( .a(n_4455), .b(n_2845), .c(n_4454), .d(n_4453), .o(n_6140) );
oa22f80 g564701 ( .a(n_4452), .b(n_4451), .c(n_4450), .d(n_4449), .o(n_6176) );
oa22f80 g564702 ( .a(n_4448), .b(n_4447), .c(n_4446), .d(n_4445), .o(n_6220) );
oa22f80 g564703 ( .a(n_4444), .b(n_3372), .c(n_3373), .d(n_4443), .o(n_6079) );
oa22f80 g564704 ( .a(n_2318), .b(x_in_9_1), .c(n_3758), .d(x_in_9_0), .o(n_7964) );
oa22f80 g564705 ( .a(n_4442), .b(n_3135), .c(n_3136), .d(n_4441), .o(n_6129) );
oa22f80 g564706 ( .a(n_4440), .b(n_3420), .c(n_3421), .d(n_4439), .o(n_5725) );
oa22f80 g564707 ( .a(n_4438), .b(n_4437), .c(n_4436), .d(n_4435), .o(n_6210) );
oa22f80 g564708 ( .a(n_4434), .b(n_4433), .c(n_4432), .d(n_4431), .o(n_6207) );
oa22f80 g564709 ( .a(n_4430), .b(n_3665), .c(n_3666), .d(n_4429), .o(n_6198) );
ao22s80 g564710 ( .a(n_3757), .b(n_5381), .c(n_2633), .d(x_in_41_4), .o(n_5483) );
oa12f80 g564711 ( .a(n_3102), .b(n_3101), .c(n_3100), .o(n_6087) );
oa22f80 g564712 ( .a(n_4428), .b(n_4427), .c(n_6023), .d(n_4426), .o(n_5764) );
ao22s80 g564713 ( .a(n_6015), .b(n_4110), .c(n_4111), .d(n_4425), .o(n_6076) );
ao22s80 g564714 ( .a(n_8061), .b(n_3697), .c(n_3698), .d(n_4424), .o(n_6790) );
in01f80 g564715 ( .a(n_6783), .o(n_5071) );
oa22f80 g564716 ( .a(n_2515), .b(x_in_39_7), .c(n_3098), .d(n_7325), .o(n_6783) );
oa22f80 g564717 ( .a(n_4423), .b(n_4422), .c(n_4421), .d(n_4420), .o(n_5718) );
oa12f80 g564718 ( .a(n_3352), .b(n_3351), .c(x_in_7_0), .o(n_6313) );
ao12f80 g564719 ( .a(n_2999), .b(n_4419), .c(x_in_3_3), .o(n_7662) );
oa22f80 g564720 ( .a(n_3156), .b(n_3756), .c(n_3157), .d(n_3755), .o(n_7404) );
oa12f80 g564721 ( .a(n_3021), .b(n_3849), .c(n_3753), .o(n_10739) );
in01f80 g564722 ( .a(n_4417), .o(n_4418) );
oa22f80 g564723 ( .a(n_3752), .b(x_in_41_11), .c(n_3751), .d(n_11409), .o(n_4417) );
ao22s80 g564724 ( .a(n_8063), .b(n_3507), .c(n_3508), .d(n_4416), .o(n_6862) );
in01f80 g564725 ( .a(n_7502), .o(n_4947) );
ao22s80 g564726 ( .a(n_4168), .b(n_8133), .c(n_2491), .d(x_in_39_8), .o(n_7502) );
ao22s80 g564727 ( .a(n_4170), .b(n_4166), .c(n_6032), .d(n_4165), .o(n_6126) );
ao22s80 g564728 ( .a(n_3749), .b(n_4946), .c(n_2686), .d(x_in_15_2), .o(n_5457) );
ao22s80 g564729 ( .a(n_2562), .b(x_in_27_5), .c(n_2050), .d(n_3747), .o(n_3748) );
ao22s80 g564730 ( .a(n_8067), .b(n_4105), .c(n_4106), .d(n_4415), .o(n_6841) );
oa22f80 g564731 ( .a(n_4414), .b(n_3119), .c(n_3120), .d(n_4413), .o(n_6188) );
oa22f80 g564732 ( .a(n_3393), .b(x_in_17_6), .c(n_2035), .d(n_5362), .o(n_5465) );
oa22f80 g564733 ( .a(n_4186), .b(n_4090), .c(n_4091), .d(n_4185), .o(n_6205) );
ao22s80 g564734 ( .a(n_4639), .b(n_2278), .c(n_4376), .d(x_in_37_3), .o(n_7605) );
oa22f80 g564735 ( .a(n_4199), .b(n_3450), .c(n_3451), .d(n_4198), .o(n_6105) );
oa22f80 g564736 ( .a(n_2017), .b(n_2004), .c(n_5679), .d(n_3747), .o(n_11679) );
ao22s80 g564737 ( .a(n_4210), .b(n_3662), .c(n_3663), .d(n_4209), .o(n_6092) );
ao22s80 g564738 ( .a(n_2149), .b(n_4148), .c(n_3746), .d(x_in_21_3), .o(n_7672) );
ao22s80 g564739 ( .a(n_3417), .b(n_2233), .c(x_in_3_5), .d(x_in_3_4), .o(n_11163) );
ao12f80 g564740 ( .a(n_3099), .b(n_3291), .c(x_in_39_4), .o(n_7019) );
ao22s80 g564741 ( .a(n_6021), .b(n_3669), .c(n_3670), .d(n_4145), .o(n_6065) );
oa22f80 g564742 ( .a(n_4412), .b(n_3672), .c(n_3673), .d(n_4411), .o(n_6053) );
oa22f80 g564743 ( .a(n_4410), .b(n_4409), .c(n_4122), .d(x_in_59_15), .o(n_6234) );
oa12f80 g564744 ( .a(n_3350), .b(n_3741), .c(n_4408), .o(n_6068) );
oa22f80 g564745 ( .a(n_4225), .b(n_2886), .c(n_4224), .d(n_4223), .o(n_6084) );
oa12f80 g564746 ( .a(n_2729), .b(n_2540), .c(x_in_5_1), .o(n_6808) );
in01f80 g564747 ( .a(n_4985), .o(n_4986) );
oa22f80 g564748 ( .a(n_4232), .b(n_4231), .c(n_4957), .d(n_4099), .o(n_4985) );
in01f80 g564749 ( .a(n_7552), .o(n_4987) );
ao22s80 g564750 ( .a(n_2708), .b(n_6500), .c(n_2322), .d(x_in_39_6), .o(n_7552) );
ao22s80 g564751 ( .a(n_3076), .b(n_3744), .c(n_4492), .d(n_5430), .o(n_3745) );
ao22s80 g564752 ( .a(n_2781), .b(n_3482), .c(n_3481), .d(n_4946), .o(n_3483) );
ao22s80 g564753 ( .a(n_2753), .b(n_3445), .c(n_4490), .d(n_5365), .o(n_3446) );
ao22s80 g564754 ( .a(n_3131), .b(n_3742), .c(n_3741), .d(n_5336), .o(n_3743) );
ao22s80 g564755 ( .a(n_3293), .b(n_3739), .c(n_4210), .d(n_5373), .o(n_3740) );
ao22s80 g564756 ( .a(n_3289), .b(n_3737), .c(n_4218), .d(n_5351), .o(n_3738) );
oa22f80 g564757 ( .a(n_2835), .b(x_in_13_11), .c(n_3077), .d(n_2834), .o(n_4836) );
in01f80 g564758 ( .a(n_4406), .o(n_4407) );
oa22f80 g564759 ( .a(n_5716), .b(n_3126), .c(n_3127), .d(x_in_37_0), .o(n_4406) );
oa22f80 g564760 ( .a(n_2453), .b(x_in_5_6), .c(n_6875), .d(x_in_5_5), .o(n_5649) );
oa22f80 g564761 ( .a(n_2330), .b(n_5271), .c(n_2226), .d(x_in_59_4), .o(n_5503) );
in01f80 g564762 ( .a(n_8952), .o(n_6225) );
oa22f80 g564763 ( .a(n_2033), .b(x_in_53_14), .c(n_2656), .d(n_2762), .o(n_8952) );
in01f80 g564764 ( .a(n_4303), .o(n_4304) );
ao22s80 g564765 ( .a(n_3025), .b(n_2834), .c(n_4231), .d(n_5926), .o(n_4303) );
oa22f80 g564766 ( .a(n_3170), .b(n_3186), .c(x_in_49_14), .d(x_in_49_11), .o(n_3171) );
ao22s80 g564767 ( .a(n_2267), .b(n_3043), .c(n_2268), .d(x_in_21_14), .o(n_8627) );
oa22f80 g564768 ( .a(n_2599), .b(n_3736), .c(n_2247), .d(x_in_29_14), .o(n_6476) );
oa22f80 g564769 ( .a(n_2198), .b(n_4042), .c(n_2949), .d(x_in_53_0), .o(n_5559) );
oa22f80 g564770 ( .a(n_2122), .b(n_2605), .c(n_3309), .d(x_in_61_0), .o(n_5603) );
in01f80 g564771 ( .a(n_3735), .o(n_4961) );
oa22f80 g564772 ( .a(n_4325), .b(x_in_19_2), .c(n_3174), .d(n_5252), .o(n_3735) );
in01f80 g564773 ( .a(n_9840), .o(n_4404) );
ao22s80 g564774 ( .a(n_5723), .b(x_in_49_14), .c(n_5835), .d(n_9118), .o(n_9840) );
ao22s80 g564775 ( .a(n_6843), .b(x_in_17_9), .c(n_3734), .d(x_in_17_10), .o(n_4999) );
in01f80 g564776 ( .a(n_3733), .o(n_5591) );
oa22f80 g564777 ( .a(n_3261), .b(x_in_59_2), .c(n_3260), .d(n_3259), .o(n_3733) );
ao22s80 g564778 ( .a(n_6878), .b(x_in_17_6), .c(n_3732), .d(x_in_17_7), .o(n_5617) );
oa22f80 g564779 ( .a(n_4403), .b(x_in_53_13), .c(n_4402), .d(n_5988), .o(n_6201) );
ao22s80 g564780 ( .a(n_6872), .b(x_in_17_8), .c(n_3731), .d(x_in_17_9), .o(n_5612) );
ao22s80 g564781 ( .a(n_4401), .b(n_5838), .c(n_8539), .d(n_3659), .o(n_7622) );
ao22s80 g564782 ( .a(n_5344), .b(n_3763), .c(x_in_19_4), .d(x_in_19_2), .o(n_5535) );
in01f80 g564783 ( .a(n_3730), .o(n_5684) );
oa22f80 g564784 ( .a(n_3262), .b(x_in_51_9), .c(n_5283), .d(n_6420), .o(n_3730) );
in01f80 g564785 ( .a(n_7455), .o(n_6303) );
no02f80 g564786 ( .a(n_2619), .b(n_2241), .o(n_7455) );
ao22s80 g564787 ( .a(n_3838), .b(n_5252), .c(x_in_19_6), .d(x_in_19_4), .o(n_5555) );
ao22s80 g564788 ( .a(n_3841), .b(n_5940), .c(x_in_19_10), .d(x_in_19_8), .o(n_5682) );
in01f80 g564789 ( .a(n_5487), .o(n_4400) );
ao22s80 g564790 ( .a(n_3849), .b(n_5326), .c(x_in_19_9), .d(x_in_19_7), .o(n_5487) );
ao22s80 g564791 ( .a(n_3729), .b(n_3174), .c(x_in_19_8), .d(x_in_19_6), .o(n_5664) );
ao22s80 g564792 ( .a(n_4664), .b(n_5939), .c(x_in_19_7), .d(x_in_19_5), .o(n_5538) );
in01f80 g564793 ( .a(n_3728), .o(n_5488) );
oa22f80 g564794 ( .a(n_5938), .b(x_in_19_9), .c(n_3020), .d(n_5244), .o(n_3728) );
ao22s80 g564795 ( .a(n_3781), .b(n_5554), .c(x_in_19_11), .d(x_in_19_9), .o(n_5557) );
in01f80 g564796 ( .a(n_6728), .o(n_4399) );
ao22s80 g564797 ( .a(n_4027), .b(n_2864), .c(n_3056), .d(x_in_29_11), .o(n_6728) );
oa22f80 g564798 ( .a(n_5115), .b(x_in_29_2), .c(n_3172), .d(n_3470), .o(n_6626) );
oa22f80 g564799 ( .a(n_15752), .b(x_in_5_12), .c(n_3169), .d(x_in_5_15), .o(n_5540) );
ao22s80 g564800 ( .a(n_4226), .b(n_3390), .c(n_2543), .d(x_in_29_9), .o(n_6007) );
ao22s80 g564801 ( .a(n_3725), .b(n_3724), .c(n_2876), .d(x_in_29_7), .o(n_5471) );
oa22f80 g564802 ( .a(n_4172), .b(x_in_29_7), .c(n_3225), .d(n_8537), .o(n_6629) );
oa22f80 g564803 ( .a(n_2644), .b(x_in_29_3), .c(n_3206), .d(n_3390), .o(n_6005) );
oa22f80 g564804 ( .a(n_9336), .b(n_4021), .c(n_3723), .d(x_in_17_4), .o(n_8662) );
in01f80 g564805 ( .a(n_6743), .o(n_4802) );
ao22s80 g564806 ( .a(n_4089), .b(n_3470), .c(n_2865), .d(x_in_29_8), .o(n_6743) );
in01f80 g564807 ( .a(n_4805), .o(n_5736) );
oa22f80 g564808 ( .a(n_3477), .b(n_5699), .c(n_3259), .d(x_in_59_4), .o(n_4805) );
no02f80 g564809 ( .a(n_4076), .b(x_in_39_4), .o(n_4077) );
na02f80 g564810 ( .a(n_4521), .b(x_in_23_0), .o(n_3219) );
na02f80 g564811 ( .a(n_3872), .b(x_in_15_15), .o(n_3873) );
na02f80 g564812 ( .a(n_4582), .b(x_in_47_0), .o(n_3168) );
na02f80 g564813 ( .a(n_3870), .b(x_in_47_15), .o(n_3871) );
na02f80 g564814 ( .a(n_2628), .b(x_in_1_2), .o(n_2531) );
na02f80 g564815 ( .a(n_4450), .b(x_in_55_0), .o(n_3167) );
na02f80 g564816 ( .a(n_4258), .b(x_in_31_0), .o(n_3166) );
na02f80 g564817 ( .a(n_3504), .b(x_in_63_15), .o(n_3505) );
no02f80 g564818 ( .a(n_2382), .b(x_in_57_2), .o(n_10986) );
na02f80 g564819 ( .a(n_4461), .b(x_in_63_0), .o(n_3163) );
in01f80 g564820 ( .a(n_3993), .o(n_5282) );
na02f80 g564821 ( .a(n_2851), .b(n_2573), .o(n_3993) );
na02f80 g564822 ( .a(n_2625), .b(x_in_39_15), .o(n_4097) );
in01f80 g564823 ( .a(n_10970), .o(n_3162) );
no02f80 g564824 ( .a(n_2599), .b(x_in_29_14), .o(n_10970) );
na02f80 g564825 ( .a(n_3287), .b(x_in_15_0), .o(n_3161) );
in01f80 g564826 ( .a(n_4043), .o(n_4044) );
na02f80 g564827 ( .a(n_2161), .b(n_3224), .o(n_4043) );
in01f80 g564828 ( .a(n_3721), .o(n_3722) );
na02f80 g564829 ( .a(n_2157), .b(n_3160), .o(n_3721) );
in01f80 g564830 ( .a(n_3719), .o(n_3720) );
na02f80 g564831 ( .a(n_2170), .b(n_2810), .o(n_3719) );
in01f80 g564832 ( .a(n_3717), .o(n_3718) );
na02f80 g564833 ( .a(n_2187), .b(n_2755), .o(n_3717) );
in01f80 g564834 ( .a(n_4046), .o(n_4047) );
na02f80 g564835 ( .a(n_2193), .b(n_3065), .o(n_4046) );
no02f80 g564836 ( .a(n_2172), .b(n_2813), .o(n_6403) );
in01f80 g564837 ( .a(n_3714), .o(n_3715) );
na02f80 g564838 ( .a(n_2176), .b(n_2703), .o(n_3714) );
in01f80 g564839 ( .a(n_3712), .o(n_3713) );
na02f80 g564840 ( .a(n_2153), .b(n_2709), .o(n_3712) );
in01f80 g564841 ( .a(n_3710), .o(n_3711) );
na02f80 g564842 ( .a(n_2228), .b(n_3341), .o(n_3710) );
in01f80 g564843 ( .a(n_3830), .o(n_3831) );
na02f80 g564844 ( .a(n_2163), .b(n_2748), .o(n_3830) );
no02f80 g564845 ( .a(n_2159), .b(n_3267), .o(n_28024) );
in01f80 g564846 ( .a(n_3708), .o(n_3709) );
na02f80 g564847 ( .a(n_2180), .b(n_3230), .o(n_3708) );
in01f80 g564848 ( .a(n_4118), .o(n_4119) );
na02f80 g564849 ( .a(n_2262), .b(n_3249), .o(n_4118) );
in01f80 g564850 ( .a(n_4007), .o(n_4008) );
na02f80 g564851 ( .a(n_2167), .b(n_3155), .o(n_4007) );
in01f80 g564852 ( .a(n_3406), .o(n_3407) );
na02f80 g564853 ( .a(n_2195), .b(n_2874), .o(n_3406) );
in01f80 g564854 ( .a(n_4050), .o(n_4051) );
na02f80 g564855 ( .a(n_2197), .b(n_3247), .o(n_4050) );
in01f80 g564856 ( .a(n_4048), .o(n_4049) );
na02f80 g564857 ( .a(n_2178), .b(n_3268), .o(n_4048) );
in01f80 g564858 ( .a(n_3706), .o(n_3707) );
na02f80 g564859 ( .a(n_2165), .b(n_3060), .o(n_3706) );
in01f80 g564860 ( .a(n_3615), .o(n_3616) );
na02f80 g564861 ( .a(n_2155), .b(n_3154), .o(n_3615) );
in01f80 g564862 ( .a(n_4066), .o(n_4067) );
na02f80 g564863 ( .a(n_2189), .b(n_2704), .o(n_4066) );
in01f80 g564864 ( .a(n_4074), .o(n_4075) );
na02f80 g564865 ( .a(n_2174), .b(n_3153), .o(n_4074) );
in01f80 g564866 ( .a(n_4126), .o(n_4127) );
na02f80 g564867 ( .a(n_2258), .b(n_3254), .o(n_4126) );
in01f80 g564868 ( .a(n_3704), .o(n_3705) );
na02f80 g564869 ( .a(n_2191), .b(n_3272), .o(n_3704) );
in01f80 g564870 ( .a(n_3702), .o(n_3703) );
na02f80 g564871 ( .a(n_2182), .b(n_3271), .o(n_3702) );
in01f80 g564872 ( .a(n_4086), .o(n_4087) );
na02f80 g564873 ( .a(n_2251), .b(n_3152), .o(n_4086) );
no02f80 g564874 ( .a(n_2266), .b(n_3256), .o(n_6412) );
in01f80 g564875 ( .a(n_3700), .o(n_3701) );
na02f80 g564876 ( .a(n_2184), .b(n_3258), .o(n_3700) );
na02f80 g564877 ( .a(n_2532), .b(x_in_55_15), .o(n_3855) );
na02f80 g564878 ( .a(n_2401), .b(x_in_23_15), .o(n_3863) );
na02f80 g564879 ( .a(n_2596), .b(x_in_31_15), .o(n_3973) );
in01f80 g564880 ( .a(n_5250), .o(n_4892) );
na02f80 g564881 ( .a(n_2590), .b(n_5435), .o(n_5250) );
in01f80 g564882 ( .a(n_3253), .o(n_4751) );
na02f80 g564883 ( .a(n_2628), .b(n_1036), .o(n_3253) );
in01f80 g564884 ( .a(n_4832), .o(n_3150) );
no02f80 g564885 ( .a(n_2590), .b(n_5435), .o(n_4832) );
no02f80 g564886 ( .a(n_5105), .b(x_in_51_2), .o(n_11603) );
in01f80 g564887 ( .a(n_7385), .o(n_6580) );
na02f80 g564888 ( .a(n_3215), .b(n_9187), .o(n_7385) );
in01f80 g564889 ( .a(n_6532), .o(n_5197) );
no02f80 g564890 ( .a(n_3215), .b(x_in_39_4), .o(n_6532) );
in01f80 g564891 ( .a(n_4396), .o(n_6521) );
no02f80 g564892 ( .a(n_4035), .b(n_3864), .o(n_4396) );
in01f80 g564893 ( .a(n_9429), .o(n_3221) );
no02f80 g564894 ( .a(n_7887), .b(x_in_21_0), .o(n_9429) );
no02f80 g564895 ( .a(n_4763), .b(x_in_21_2), .o(n_11597) );
na02f80 g564896 ( .a(n_3101), .b(n_3100), .o(n_3102) );
no02f80 g564897 ( .a(n_4863), .b(x_in_37_2), .o(n_11594) );
no02f80 g564898 ( .a(n_2617), .b(x_in_41_8), .o(n_7215) );
no02f80 g564899 ( .a(n_2610), .b(x_in_41_6), .o(n_3876) );
no02f80 g564900 ( .a(n_4822), .b(x_in_41_5), .o(n_4003) );
in01f80 g564901 ( .a(n_3869), .o(n_3148) );
no02f80 g564902 ( .a(n_3868), .b(x_in_41_4), .o(n_3869) );
no02f80 g564903 ( .a(n_3274), .b(n_3273), .o(n_3275) );
na02f80 g564904 ( .a(n_4060), .b(n_4059), .o(n_4061) );
no02f80 g564905 ( .a(n_3157), .b(n_3156), .o(n_3158) );
na02f80 g564906 ( .a(n_2656), .b(x_in_53_14), .o(n_8769) );
na02f80 g564907 ( .a(n_2686), .b(n_4946), .o(n_2687) );
na02f80 g564908 ( .a(n_2565), .b(n_5336), .o(n_2566) );
na02f80 g564909 ( .a(n_2571), .b(n_5351), .o(n_2572) );
na02f80 g564910 ( .a(n_3287), .b(n_4457), .o(n_3147) );
na02f80 g564911 ( .a(n_4103), .b(n_4102), .o(n_4104) );
na02f80 g564912 ( .a(n_4116), .b(n_4115), .o(n_4117) );
na02f80 g564913 ( .a(n_4106), .b(n_4105), .o(n_4107) );
in01f80 g564914 ( .a(n_10121), .o(n_2884) );
no02f80 g564915 ( .a(n_2851), .b(n_2636), .o(n_10121) );
na02f80 g564916 ( .a(n_2630), .b(n_448), .o(n_2631) );
na02f80 g564917 ( .a(n_23345), .b(n_2096), .o(n_23072) );
na02f80 g564918 ( .a(n_4476), .b(n_3511), .o(n_3512) );
na02f80 g564919 ( .a(n_4454), .b(n_2845), .o(n_2846) );
no02f80 g564920 ( .a(n_3144), .b(n_2040), .o(n_3080) );
na02f80 g564921 ( .a(n_3698), .b(n_3697), .o(n_3699) );
na02f80 g564922 ( .a(n_3695), .b(n_3694), .o(n_3696) );
na02f80 g564923 ( .a(n_3508), .b(n_3507), .o(n_3509) );
in01f80 g564924 ( .a(n_5822), .o(n_5854) );
na02f80 g564925 ( .a(n_3146), .b(n_3175), .o(n_5822) );
na02f80 g564926 ( .a(n_3773), .b(x_in_29_15), .o(n_3279) );
no02f80 g564927 ( .a(n_2570), .b(n_3641), .o(n_3642) );
na02f80 g564928 ( .a(n_2145), .b(n_5700), .o(n_4760) );
na02f80 g564929 ( .a(n_4481), .b(n_3692), .o(n_3693) );
na02f80 g564930 ( .a(n_3144), .b(n_4479), .o(n_3145) );
no02f80 g564931 ( .a(n_2132), .b(n_3771), .o(n_2862) );
na02f80 g564932 ( .a(n_2043), .b(n_3143), .o(n_8114) );
no02f80 g564933 ( .a(n_3141), .b(n_3140), .o(n_3142) );
no02f80 g564934 ( .a(n_2839), .b(n_2838), .o(n_2840) );
in01f80 g564935 ( .a(n_3689), .o(n_5049) );
na02f80 g564936 ( .a(n_2045), .b(n_2746), .o(n_3689) );
no02f80 g564937 ( .a(n_3285), .b(n_3284), .o(n_3286) );
no02f80 g564938 ( .a(n_3282), .b(n_3281), .o(n_3283) );
na02f80 g564939 ( .a(n_2276), .b(n_3138), .o(n_3139) );
no02f80 g564940 ( .a(n_3136), .b(n_3135), .o(n_3137) );
in01f80 g564941 ( .a(n_3996), .o(n_3134) );
na02f80 g564942 ( .a(n_2364), .b(n_8522), .o(n_3996) );
no02f80 g564943 ( .a(n_3687), .b(n_3686), .o(n_3688) );
no02f80 g564944 ( .a(n_2054), .b(n_3132), .o(n_3133) );
in01f80 g564945 ( .a(n_6530), .o(n_3685) );
no02f80 g564946 ( .a(n_3076), .b(x_in_23_4), .o(n_6530) );
in01f80 g564947 ( .a(n_6528), .o(n_3684) );
no02f80 g564948 ( .a(n_2781), .b(x_in_15_4), .o(n_6528) );
no02f80 g564949 ( .a(n_3287), .b(n_2207), .o(n_3288) );
in01f80 g564950 ( .a(n_4921), .o(n_3683) );
no02f80 g564951 ( .a(n_3289), .b(x_in_63_4), .o(n_4921) );
in01f80 g564952 ( .a(n_6526), .o(n_3394) );
no02f80 g564953 ( .a(n_2753), .b(x_in_47_4), .o(n_6526) );
in01f80 g564954 ( .a(n_6524), .o(n_3682) );
no02f80 g564955 ( .a(n_3131), .b(x_in_55_4), .o(n_6524) );
in01f80 g564956 ( .a(n_6522), .o(n_4120) );
no02f80 g564957 ( .a(n_3293), .b(x_in_31_4), .o(n_6522) );
na02f80 g564958 ( .a(n_4094), .b(n_4093), .o(n_4095) );
na02f80 g564959 ( .a(n_5264), .b(n_2705), .o(n_2706) );
no02f80 g564960 ( .a(n_4091), .b(n_4090), .o(n_4092) );
na02f80 g564961 ( .a(n_3292), .b(n_3291), .o(n_8367) );
na02f80 g564962 ( .a(n_3351), .b(x_in_7_0), .o(n_3352) );
in01f80 g564963 ( .a(n_3680), .o(n_3681) );
no02f80 g564964 ( .a(n_2142), .b(n_3242), .o(n_3680) );
in01f80 g564965 ( .a(n_3678), .o(n_3679) );
na02f80 g564966 ( .a(n_2716), .b(n_2715), .o(n_3678) );
no02f80 g564967 ( .a(n_2129), .b(n_5317), .o(n_2722) );
no02f80 g564968 ( .a(n_2074), .b(n_3129), .o(n_3130) );
in01f80 g564969 ( .a(n_3676), .o(n_3677) );
no02f80 g564970 ( .a(n_2103), .b(n_2768), .o(n_3676) );
in01f80 g564971 ( .a(n_5980), .o(n_10817) );
no02f80 g564972 ( .a(n_4742), .b(n_7840), .o(n_5980) );
na02f80 g564973 ( .a(n_2633), .b(n_5381), .o(n_2634) );
na02f80 g564974 ( .a(n_2617), .b(n_9612), .o(n_2569) );
no02f80 g564975 ( .a(n_3127), .b(n_3126), .o(n_3128) );
na02f80 g564976 ( .a(n_7070), .b(x_in_25_9), .o(n_2568) );
no02f80 g564977 ( .a(n_7070), .b(x_in_25_9), .o(n_2295) );
in01f80 g564978 ( .a(n_4585), .o(n_3675) );
na02f80 g564979 ( .a(n_5407), .b(n_9329), .o(n_4585) );
na02f80 g564980 ( .a(n_2610), .b(n_9610), .o(n_2314) );
in01f80 g564981 ( .a(n_2738), .o(n_2739) );
no02f80 g564982 ( .a(n_2641), .b(x_in_41_7), .o(n_2738) );
na02f80 g564983 ( .a(n_3481), .b(n_4486), .o(n_3125) );
na02f80 g564984 ( .a(n_3741), .b(n_4408), .o(n_3350) );
no02f80 g564985 ( .a(n_2126), .b(n_2743), .o(n_2744) );
in01f80 g564986 ( .a(n_6434), .o(n_6425) );
na02f80 g564987 ( .a(n_3156), .b(n_3124), .o(n_6434) );
no02f80 g564988 ( .a(n_4130), .b(n_4129), .o(n_4131) );
no02f80 g564989 ( .a(n_3295), .b(n_3294), .o(n_3296) );
no02f80 g564990 ( .a(n_2760), .b(n_2759), .o(n_2761) );
in01f80 g564991 ( .a(n_5755), .o(n_3396) );
na02f80 g564992 ( .a(n_2114), .b(n_4151), .o(n_5755) );
no02f80 g564993 ( .a(n_2127), .b(n_3189), .o(n_2778) );
no02f80 g564994 ( .a(n_9975), .b(x_in_49_5), .o(n_2637) );
no02f80 g564995 ( .a(n_6667), .b(x_in_37_1), .o(n_2619) );
in01f80 g564996 ( .a(n_5832), .o(n_3427) );
na02f80 g564997 ( .a(n_2795), .b(n_2794), .o(n_5832) );
no02f80 g564998 ( .a(n_3481), .b(n_2217), .o(n_3297) );
no02f80 g564999 ( .a(n_7099), .b(n_2567), .o(n_4814) );
no02f80 g565000 ( .a(n_4523), .b(n_3122), .o(n_3123) );
no02f80 g565001 ( .a(n_3120), .b(n_3119), .o(n_3121) );
no02f80 g565002 ( .a(n_4515), .b(n_4516), .o(n_2792) );
na02f80 g565003 ( .a(n_7099), .b(n_2567), .o(n_4813) );
no02f80 g565004 ( .a(n_3673), .b(n_3672), .o(n_3674) );
no02f80 g565005 ( .a(n_3421), .b(n_3420), .o(n_3422) );
no02f80 g565006 ( .a(n_4498), .b(n_2693), .o(n_2694) );
na02f80 g565007 ( .a(n_3670), .b(n_3669), .o(n_3671) );
no02f80 g565008 ( .a(n_3328), .b(n_3327), .o(n_3329) );
no02f80 g565009 ( .a(n_3339), .b(n_3338), .o(n_3340) );
na02f80 g565010 ( .a(n_3432), .b(n_3431), .o(n_3433) );
na02f80 g565011 ( .a(n_2146), .b(x_in_19_0), .o(n_9205) );
na02f80 g565012 ( .a(n_7102), .b(n_2434), .o(n_4807) );
no02f80 g565013 ( .a(n_7102), .b(n_2434), .o(n_4809) );
na02f80 g565014 ( .a(n_2389), .b(x_in_45_15), .o(n_3668) );
no02f80 g565015 ( .a(n_4884), .b(n_2815), .o(n_2816) );
no02f80 g565016 ( .a(n_3741), .b(n_2055), .o(n_3118) );
in01f80 g565017 ( .a(n_4029), .o(n_3117) );
no02f80 g565018 ( .a(n_2584), .b(x_in_41_5), .o(n_4029) );
na02f80 g565019 ( .a(n_3025), .b(x_in_13_13), .o(n_7895) );
in01f80 g565020 ( .a(n_8519), .o(n_7723) );
na02f80 g565021 ( .a(n_2221), .b(n_2696), .o(n_8519) );
na02f80 g565022 ( .a(n_7124), .b(n_5311), .o(n_2640) );
no02f80 g565023 ( .a(n_3373), .b(n_3372), .o(n_3374) );
no02f80 g565024 ( .a(n_3451), .b(n_3450), .o(n_3452) );
no02f80 g565025 ( .a(n_3666), .b(n_3665), .o(n_3667) );
no02f80 g565026 ( .a(n_4135), .b(n_4134), .o(n_4136) );
na02f80 g565027 ( .a(n_3460), .b(n_3459), .o(n_3461) );
no02f80 g565028 ( .a(n_3468), .b(n_3467), .o(n_3469) );
na02f80 g565029 ( .a(n_3663), .b(n_3662), .o(n_3664) );
no02f80 g565030 ( .a(n_4373), .b(n_4374), .o(n_3269) );
in01f80 g565031 ( .a(n_7807), .o(n_8451) );
na02f80 g565032 ( .a(n_2700), .b(n_3351), .o(n_7807) );
in01f80 g565033 ( .a(n_11226), .o(n_3277) );
na02f80 g565034 ( .a(n_2676), .b(n_5245), .o(n_11226) );
na02f80 g565035 ( .a(n_2614), .b(n_7915), .o(n_2615) );
no02f80 g565036 ( .a(n_3115), .b(n_3114), .o(n_3116) );
no02f80 g565037 ( .a(n_3301), .b(n_3300), .o(n_3302) );
no02f80 g565038 ( .a(n_3307), .b(n_3306), .o(n_3308) );
in01f80 g565039 ( .a(n_3529), .o(n_3113) );
na02f80 g565040 ( .a(n_2453), .b(n_3568), .o(n_3529) );
in01f80 g565041 ( .a(n_3661), .o(n_10897) );
no02f80 g565042 ( .a(n_2856), .b(n_2855), .o(n_3661) );
in01f80 g565043 ( .a(n_9146), .o(n_3490) );
na02f80 g565044 ( .a(n_2708), .b(x_in_39_6), .o(n_9146) );
no02f80 g565045 ( .a(n_3617), .b(x_in_57_3), .o(n_3112) );
na02f80 g565046 ( .a(n_7887), .b(n_2066), .o(n_2586) );
na02f80 g565047 ( .a(n_2880), .b(x_in_41_13), .o(n_7884) );
na02f80 g565048 ( .a(n_4111), .b(n_4110), .o(n_4112) );
no02f80 g565049 ( .a(n_4548), .b(n_2866), .o(n_2867) );
na02f80 g565050 ( .a(n_4903), .b(x_in_49_15), .o(n_2871) );
no02f80 g565051 ( .a(n_4224), .b(n_2886), .o(n_2887) );
no02f80 g565052 ( .a(n_4469), .b(n_2881), .o(n_2882) );
no02f80 g565053 ( .a(n_4389), .b(n_3110), .o(n_3111) );
in01f80 g565054 ( .a(n_3383), .o(n_2885) );
na02f80 g565055 ( .a(n_2562), .b(n_3747), .o(n_3383) );
na02f80 g565056 ( .a(n_2255), .b(x_in_21_5), .o(n_2889) );
no02f80 g565057 ( .a(n_2789), .b(n_2254), .o(n_4149) );
no02f80 g565058 ( .a(n_7776), .b(n_3261), .o(n_7932) );
in01f80 g565059 ( .a(n_3404), .o(n_3109) );
na02f80 g565060 ( .a(n_3177), .b(n_5327), .o(n_3404) );
na02f80 g565061 ( .a(n_2135), .b(n_2798), .o(n_5223) );
na02f80 g565062 ( .a(n_2587), .b(n_3568), .o(n_3569) );
na02f80 g565063 ( .a(n_3659), .b(n_5838), .o(n_3660) );
in01f80 g565064 ( .a(n_10299), .o(n_2900) );
no02f80 g565065 ( .a(n_7554), .b(x_in_61_10), .o(n_10299) );
na02f80 g565066 ( .a(n_2741), .b(x_in_37_6), .o(n_2811) );
na02f80 g565067 ( .a(n_2741), .b(x_in_37_1), .o(n_2742) );
in01f80 g565068 ( .a(n_10017), .o(n_2922) );
no02f80 g565069 ( .a(n_7443), .b(x_in_61_6), .o(n_10017) );
no02f80 g565070 ( .a(n_7054), .b(n_2365), .o(n_11568) );
no02f80 g565071 ( .a(n_7051), .b(n_2664), .o(n_11565) );
no02f80 g565072 ( .a(n_5596), .b(x_in_61_5), .o(n_10894) );
in01f80 g565073 ( .a(n_4783), .o(n_5908) );
na02f80 g565074 ( .a(n_2950), .b(n_2949), .o(n_4783) );
no02f80 g565075 ( .a(n_4004), .b(n_5703), .o(n_6966) );
in01f80 g565076 ( .a(n_3658), .o(n_9139) );
no02f80 g565077 ( .a(n_3291), .b(n_3107), .o(n_3658) );
in01f80 g565078 ( .a(n_7844), .o(n_8509) );
na02f80 g565079 ( .a(n_3310), .b(n_3309), .o(n_7844) );
in01f80 g565080 ( .a(n_10004), .o(n_4385) );
no02f80 g565081 ( .a(n_3576), .b(x_in_61_7), .o(n_10004) );
no02f80 g565082 ( .a(n_6767), .b(x_in_61_9), .o(n_10889) );
na02f80 g565083 ( .a(n_3015), .b(n_2877), .o(n_4710) );
na02f80 g565084 ( .a(n_2471), .b(x_in_59_4), .o(n_3594) );
in01f80 g565085 ( .a(n_3657), .o(n_10879) );
no02f80 g565086 ( .a(n_3056), .b(n_2875), .o(n_3657) );
no02f80 g565087 ( .a(n_4011), .b(x_in_33_3), .o(n_3066) );
no02f80 g565088 ( .a(n_7076), .b(n_2509), .o(n_10622) );
in01f80 g565089 ( .a(n_4696), .o(n_4098) );
na02f80 g565090 ( .a(n_5230), .b(n_3072), .o(n_4696) );
na02f80 g565092 ( .a(n_3073), .b(n_3070), .o(n_5232) );
na02f80 g565094 ( .a(n_3106), .b(n_2879), .o(n_5229) );
no02f80 g565095 ( .a(n_3723), .b(n_4021), .o(n_3094) );
na02f80 g565096 ( .a(n_3173), .b(n_2077), .o(n_5227) );
no02f80 g565097 ( .a(n_2243), .b(x_in_45_12), .o(n_3105) );
in01f80 g565098 ( .a(n_9998), .o(n_3312) );
no02f80 g565099 ( .a(n_6723), .b(x_in_61_8), .o(n_9998) );
in01f80 g565100 ( .a(n_10882), .o(n_3149) );
no02f80 g565101 ( .a(n_6387), .b(x_in_61_4), .o(n_10882) );
na02f80 g565102 ( .a(n_3311), .b(n_2805), .o(n_5225) );
na02f80 g565104 ( .a(n_3104), .b(x_in_19_1), .o(n_9964) );
no02f80 g565105 ( .a(n_2319), .b(x_in_9_1), .o(n_7793) );
no02f80 g565106 ( .a(n_7048), .b(n_2420), .o(n_11548) );
na02f80 g565107 ( .a(n_3655), .b(x_in_61_15), .o(n_3656) );
no02f80 g565108 ( .a(n_7855), .b(n_5156), .o(n_12862) );
no02f80 g565109 ( .a(n_6938), .b(x_in_57_6), .o(n_2854) );
na02f80 g565110 ( .a(n_6938), .b(x_in_57_6), .o(n_3244) );
na02f80 g565112 ( .a(n_4232), .b(n_4099), .o(n_4100) );
in01f80 g565113 ( .a(n_9135), .o(n_3365) );
na02f80 g565114 ( .a(n_2767), .b(x_in_39_9), .o(n_9135) );
in01f80 g565115 ( .a(n_8737), .o(n_3570) );
na02f80 g565116 ( .a(n_3206), .b(x_in_29_6), .o(n_8737) );
na02f80 g565117 ( .a(n_2416), .b(n_3560), .o(n_3561) );
no02f80 g565118 ( .a(n_3751), .b(x_in_41_11), .o(n_3103) );
na02f80 g565119 ( .a(n_4533), .b(x_in_43_4), .o(n_3652) );
na02f80 g565120 ( .a(n_4392), .b(x_in_11_4), .o(n_3977) );
no02f80 g565121 ( .a(n_7048), .b(n_5679), .o(n_3316) );
na02f80 g565122 ( .a(n_2414), .b(n_13241), .o(n_3416) );
na02f80 g565123 ( .a(n_6926), .b(x_in_5_7), .o(n_2710) );
no02f80 g565124 ( .a(n_6926), .b(x_in_5_7), .o(n_2852) );
na02f80 g565125 ( .a(n_3172), .b(x_in_29_5), .o(n_8734) );
no02f80 g565126 ( .a(n_5226), .b(n_2533), .o(n_3370) );
in01f80 g565127 ( .a(n_9132), .o(n_3493) );
na02f80 g565128 ( .a(n_3346), .b(x_in_39_5), .o(n_9132) );
na02f80 g565129 ( .a(n_2544), .b(x_in_29_9), .o(n_8731) );
na02f80 g565130 ( .a(n_4948), .b(n_8957), .o(n_2604) );
in01f80 g565131 ( .a(n_10861), .o(n_3414) );
na02f80 g565132 ( .a(n_2809), .b(x_in_39_11), .o(n_10861) );
in01f80 g565133 ( .a(n_10866), .o(n_4031) );
na02f80 g565134 ( .a(n_12817), .b(x_in_19_13), .o(n_10866) );
in01f80 g565135 ( .a(n_8608), .o(n_4876) );
no02f80 g565136 ( .a(n_3424), .b(x_in_45_1), .o(n_8608) );
na02f80 g565137 ( .a(n_2495), .b(x_in_29_4), .o(n_8728) );
na02f80 g565138 ( .a(n_2827), .b(x_in_35_10), .o(n_9984) );
in01f80 g565139 ( .a(n_3436), .o(n_8722) );
no02f80 g565140 ( .a(n_2876), .b(n_3035), .o(n_3436) );
in01f80 g565141 ( .a(n_3651), .o(n_8725) );
no02f80 g565142 ( .a(n_2865), .b(n_2864), .o(n_3651) );
no02f80 g565143 ( .a(n_3291), .b(x_in_39_4), .o(n_3099) );
in01f80 g565144 ( .a(n_9129), .o(n_3494) );
na02f80 g565145 ( .a(n_4168), .b(x_in_39_8), .o(n_9129) );
in01f80 g565146 ( .a(n_9123), .o(n_3649) );
na02f80 g565147 ( .a(n_3098), .b(x_in_39_7), .o(n_9123) );
no02f80 g565148 ( .a(n_3848), .b(n_2650), .o(n_8655) );
na02f80 g565149 ( .a(n_2584), .b(n_2583), .o(n_2585) );
na02f80 g565150 ( .a(n_2423), .b(n_9329), .o(n_3648) );
na02f80 g565151 ( .a(n_3096), .b(x_in_29_4), .o(n_3097) );
na02f80 g565152 ( .a(n_2598), .b(x_in_45_2), .o(n_3434) );
na02f80 g565153 ( .a(n_2323), .b(n_5388), .o(n_4036) );
na02f80 g565154 ( .a(n_2751), .b(x_in_17_14), .o(n_4714) );
na02f80 g565155 ( .a(n_2623), .b(n_4057), .o(n_4045) );
na02f80 g565156 ( .a(n_2641), .b(n_9327), .o(n_2642) );
in01f80 g565157 ( .a(n_9126), .o(n_4842) );
no02f80 g565158 ( .a(n_3980), .b(x_in_25_11), .o(n_9126) );
no02f80 g565159 ( .a(n_4972), .b(n_8851), .o(n_6884) );
no02f80 g565160 ( .a(n_4030), .b(n_2595), .o(n_8636) );
na02f80 g565161 ( .a(n_3208), .b(n_2321), .o(n_4629) );
na02f80 g565162 ( .a(n_9095), .b(x_in_41_5), .o(n_5688) );
in01f80 g565163 ( .a(n_9969), .o(n_4037) );
na02f80 g565164 ( .a(n_3222), .b(x_in_35_5), .o(n_9969) );
na02f80 g565165 ( .a(n_6892), .b(x_in_57_8), .o(n_2702) );
in01f80 g565166 ( .a(n_9120), .o(n_4028) );
na02f80 g565167 ( .a(n_2750), .b(x_in_39_10), .o(n_9120) );
no02f80 g565168 ( .a(n_2487), .b(x_in_5_9), .o(n_3367) );
na02f80 g565169 ( .a(n_2806), .b(n_5849), .o(n_2807) );
na02f80 g565170 ( .a(n_2296), .b(n_5888), .o(n_3391) );
no02f80 g565171 ( .a(n_6892), .b(x_in_57_8), .o(n_3264) );
in01f80 g565172 ( .a(n_8719), .o(n_4128) );
na02f80 g565173 ( .a(n_3225), .b(x_in_29_10), .o(n_8719) );
na02f80 g565174 ( .a(n_2304), .b(n_4055), .o(n_4056) );
no02f80 g565175 ( .a(n_7650), .b(x_in_21_10), .o(n_3335) );
in01f80 g565176 ( .a(n_6475), .o(n_4867) );
na02f80 g565177 ( .a(n_5046), .b(x_in_29_10), .o(n_6475) );
na02f80 g565178 ( .a(n_6875), .b(n_5291), .o(n_3093) );
in01f80 g565179 ( .a(n_10236), .o(n_3647) );
no02f80 g565180 ( .a(n_2998), .b(x_in_61_1), .o(n_10236) );
na02f80 g565181 ( .a(n_2470), .b(n_5302), .o(n_4064) );
in01f80 g565182 ( .a(n_5844), .o(n_6751) );
no02f80 g565183 ( .a(n_4401), .b(n_5902), .o(n_5844) );
in01f80 g565184 ( .a(n_8647), .o(n_4840) );
na02f80 g565185 ( .a(n_3811), .b(n_2342), .o(n_8647) );
na02f80 g565186 ( .a(n_6817), .b(n_3245), .o(n_3246) );
no02f80 g565187 ( .a(n_8299), .b(x_in_37_6), .o(n_3645) );
na02f80 g565188 ( .a(n_8303), .b(n_3318), .o(n_3319) );
na02f80 g565189 ( .a(n_2837), .b(n_4687), .o(n_2561) );
in01f80 g565190 ( .a(n_9961), .o(n_3644) );
na02f80 g565191 ( .a(n_3233), .b(x_in_35_4), .o(n_9961) );
in01f80 g565192 ( .a(n_4383), .o(n_5786) );
na02f80 g565193 ( .a(n_3643), .b(x_in_41_12), .o(n_4383) );
no02f80 g565194 ( .a(n_2463), .b(x_in_21_8), .o(n_4071) );
in01f80 g565195 ( .a(n_9946), .o(n_3361) );
na02f80 g565196 ( .a(n_3257), .b(x_in_35_7), .o(n_9946) );
no02f80 g565197 ( .a(n_3041), .b(x_in_21_6), .o(n_3092) );
na02f80 g565198 ( .a(n_7690), .b(n_3887), .o(n_3888) );
in01f80 g565199 ( .a(n_9940), .o(n_4070) );
na02f80 g565200 ( .a(n_3255), .b(x_in_35_9), .o(n_9940) );
in01f80 g565201 ( .a(n_4082), .o(n_9958) );
no02f80 g565202 ( .a(n_3366), .b(n_4939), .o(n_4082) );
in01f80 g565203 ( .a(n_9896), .o(n_4078) );
na02f80 g565204 ( .a(n_3784), .b(x_in_35_6), .o(n_9896) );
na02f80 g565205 ( .a(n_2514), .b(n_3409), .o(n_3410) );
na02f80 g565206 ( .a(n_3516), .b(n_3096), .o(n_4765) );
in01f80 g565207 ( .a(n_3360), .o(n_10820) );
no02f80 g565208 ( .a(n_4903), .b(n_3186), .o(n_3360) );
no02f80 g565209 ( .a(n_3839), .b(n_2339), .o(n_8671) );
no02f80 g565210 ( .a(n_4080), .b(n_2325), .o(n_8624) );
no02f80 g565211 ( .a(n_3095), .b(x_in_37_11), .o(n_3091) );
na02f80 g565212 ( .a(n_2367), .b(n_5754), .o(n_3844) );
na02f80 g565213 ( .a(n_2300), .b(n_5754), .o(n_4081) );
na02f80 g565214 ( .a(n_2335), .b(n_5313), .o(n_3640) );
in01f80 g565215 ( .a(n_4032), .o(n_4033) );
no02f80 g565216 ( .a(n_4970), .b(n_8336), .o(n_4032) );
in01f80 g565217 ( .a(n_8664), .o(n_4381) );
na02f80 g565218 ( .a(n_3902), .b(n_2612), .o(n_8664) );
no02f80 g565219 ( .a(n_4402), .b(x_in_53_13), .o(n_3914) );
in01f80 g565220 ( .a(n_9923), .o(n_4023) );
na02f80 g565221 ( .a(n_3090), .b(x_in_35_11), .o(n_9923) );
no02f80 g565222 ( .a(n_6409), .b(n_3263), .o(n_5994) );
no02f80 g565223 ( .a(n_7790), .b(n_3263), .o(n_3089) );
na02f80 g565224 ( .a(n_6409), .b(n_6405), .o(n_5459) );
na02f80 g565225 ( .a(n_7790), .b(n_3263), .o(n_5992) );
no02f80 g565226 ( .a(n_6409), .b(n_6405), .o(n_3280) );
na02f80 g565227 ( .a(n_6409), .b(n_3263), .o(n_3088) );
no02f80 g565228 ( .a(n_3323), .b(n_6405), .o(n_4818) );
na02f80 g565229 ( .a(n_3323), .b(n_6405), .o(n_3087) );
na02f80 g565230 ( .a(n_7790), .b(n_7781), .o(n_3086) );
no02f80 g565231 ( .a(n_7790), .b(n_7781), .o(n_5990) );
no02f80 g565232 ( .a(n_7776), .b(n_7781), .o(n_3179) );
na02f80 g565233 ( .a(n_6797), .b(x_in_3_13), .o(n_3942) );
na02f80 g565234 ( .a(n_3321), .b(x_in_3_13), .o(n_9888) );
na02f80 g565235 ( .a(n_3235), .b(x_in_53_13), .o(n_3236) );
na02f80 g565236 ( .a(n_2542), .b(x_in_51_4), .o(n_3639) );
na02f80 g565237 ( .a(n_3323), .b(n_8336), .o(n_4365) );
no02f80 g565238 ( .a(n_3323), .b(n_8336), .o(n_3085) );
na02f80 g565239 ( .a(n_2454), .b(x_in_17_13), .o(n_3587) );
na02f80 g565240 ( .a(n_3638), .b(x_in_17_13), .o(n_9891) );
in01f80 g565241 ( .a(n_8632), .o(n_4878) );
na02f80 g565242 ( .a(n_3397), .b(n_2600), .o(n_8632) );
na02f80 g565243 ( .a(n_2658), .b(n_3324), .o(n_4727) );
no02f80 g565244 ( .a(n_2602), .b(n_4034), .o(n_5205) );
no02f80 g565245 ( .a(n_3834), .b(n_2369), .o(n_8682) );
in01f80 g565246 ( .a(n_5969), .o(n_5748) );
na02f80 g565247 ( .a(n_3322), .b(n_2578), .o(n_5969) );
in01f80 g565248 ( .a(n_6958), .o(n_6959) );
no02f80 g565249 ( .a(n_3385), .b(n_2497), .o(n_6958) );
in01f80 g565250 ( .a(n_7602), .o(n_3637) );
na02f80 g565251 ( .a(n_3310), .b(n_3325), .o(n_7602) );
no02f80 g565252 ( .a(n_3379), .b(n_3498), .o(n_5200) );
in01f80 g565253 ( .a(n_9594), .o(n_9334) );
na02f80 g565254 ( .a(n_3716), .b(n_2429), .o(n_9594) );
in01f80 g565255 ( .a(n_5157), .o(n_6572) );
no02f80 g565256 ( .a(n_2671), .b(n_3526), .o(n_5157) );
in01f80 g565257 ( .a(n_7571), .o(n_5144) );
na02f80 g565258 ( .a(n_2888), .b(n_2460), .o(n_7571) );
in01f80 g565259 ( .a(n_5867), .o(n_5762) );
na02f80 g565260 ( .a(n_2906), .b(n_2383), .o(n_5867) );
in01f80 g565261 ( .a(n_5706), .o(n_5705) );
na02f80 g565262 ( .a(n_2901), .b(n_2355), .o(n_5706) );
in01f80 g565263 ( .a(n_9604), .o(n_6760) );
na02f80 g565264 ( .a(n_3796), .b(n_2503), .o(n_9604) );
in01f80 g565265 ( .a(n_8489), .o(n_5801) );
na02f80 g565266 ( .a(n_2360), .b(n_3784), .o(n_8489) );
in01f80 g565267 ( .a(n_8092), .o(n_5847) );
no02f80 g565268 ( .a(n_2336), .b(n_3220), .o(n_8092) );
no02f80 g565269 ( .a(n_2519), .b(n_3634), .o(n_3635) );
no02f80 g565270 ( .a(n_3448), .b(n_2346), .o(n_3633) );
in01f80 g565271 ( .a(n_12697), .o(n_10779) );
no02f80 g565272 ( .a(n_2856), .b(n_2499), .o(n_12697) );
in01f80 g565273 ( .a(n_5149), .o(n_8023) );
no02f80 g565274 ( .a(n_2459), .b(n_3543), .o(n_5149) );
in01f80 g565275 ( .a(n_5824), .o(n_9088) );
no02f80 g565276 ( .a(n_3885), .b(n_3298), .o(n_5824) );
in01f80 g565277 ( .a(n_8920), .o(n_4379) );
no02f80 g565278 ( .a(n_2479), .b(n_3782), .o(n_8920) );
in01f80 g565279 ( .a(n_8982), .o(n_3476) );
no02f80 g565280 ( .a(n_3313), .b(n_2406), .o(n_8982) );
no02f80 g565281 ( .a(n_2306), .b(n_2844), .o(n_8618) );
in01f80 g565282 ( .a(n_9007), .o(n_5189) );
na02f80 g565283 ( .a(n_2576), .b(n_3084), .o(n_9007) );
in01f80 g565284 ( .a(n_8086), .o(n_5771) );
na02f80 g565285 ( .a(n_2674), .b(n_3083), .o(n_8086) );
no02f80 g565286 ( .a(n_2455), .b(n_3331), .o(n_5918) );
in01f80 g565287 ( .a(n_8041), .o(n_4069) );
na02f80 g565288 ( .a(n_3223), .b(n_2312), .o(n_8041) );
no02f80 g565289 ( .a(n_2297), .b(n_3248), .o(n_8108) );
na02f80 g565290 ( .a(n_2404), .b(n_3330), .o(n_9010) );
in01f80 g565291 ( .a(n_7211), .o(n_6477) );
no02f80 g565292 ( .a(n_4122), .b(n_4121), .o(n_7211) );
in01f80 g565293 ( .a(n_8089), .o(n_5840) );
no02f80 g565294 ( .a(n_2457), .b(n_3332), .o(n_8089) );
in01f80 g565295 ( .a(n_6457), .o(n_5811) );
no02f80 g565296 ( .a(n_3501), .b(n_3500), .o(n_6457) );
in01f80 g565297 ( .a(n_8103), .o(n_3499) );
na02f80 g565298 ( .a(n_2484), .b(n_3333), .o(n_8103) );
in01f80 g565299 ( .a(n_8157), .o(n_3392) );
no02f80 g565300 ( .a(n_2481), .b(n_2848), .o(n_8157) );
in01f80 g565301 ( .a(n_4748), .o(n_10553) );
no02f80 g565302 ( .a(n_2869), .b(n_2868), .o(n_4748) );
no02f80 g565303 ( .a(n_3082), .b(n_2474), .o(n_5928) );
na02f80 g565304 ( .a(n_2348), .b(n_3875), .o(n_5995) );
in01f80 g565305 ( .a(n_8494), .o(n_5799) );
no02f80 g565306 ( .a(n_2311), .b(n_3449), .o(n_8494) );
no02f80 g565307 ( .a(n_2467), .b(n_3632), .o(n_5978) );
no02f80 g565308 ( .a(n_2469), .b(n_3453), .o(n_6330) );
in01f80 g565309 ( .a(n_8142), .o(n_5828) );
no02f80 g565310 ( .a(n_2638), .b(n_2804), .o(n_8142) );
in01f80 g565311 ( .a(n_8496), .o(n_5797) );
no02f80 g565312 ( .a(n_2399), .b(n_3386), .o(n_8496) );
in01f80 g565313 ( .a(n_8491), .o(n_5780) );
no02f80 g565314 ( .a(n_2375), .b(n_3353), .o(n_8491) );
no02f80 g565315 ( .a(n_2380), .b(n_2728), .o(n_8162) );
in01f80 g565316 ( .a(n_8971), .o(n_4924) );
no02f80 g565317 ( .a(n_2621), .b(n_3081), .o(n_8971) );
in01f80 g565318 ( .a(n_7648), .o(n_4969) );
na02f80 g565319 ( .a(n_2735), .b(n_2734), .o(n_7648) );
in01f80 g565320 ( .a(n_6583), .o(n_5814) );
no02f80 g565321 ( .a(n_3389), .b(n_3388), .o(n_6583) );
oa12f80 g565322 ( .a(n_2320), .b(x_in_13_2), .c(x_in_13_1), .o(n_7197) );
oa12f80 g565323 ( .a(n_7150), .b(n_2603), .c(x_in_63_0), .o(n_4786) );
in01f80 g565324 ( .a(n_6788), .o(n_3266) );
oa12f80 g565325 ( .a(n_9171), .b(x_in_29_3), .c(x_in_29_2), .o(n_6788) );
in01f80 g565326 ( .a(n_4953), .o(n_8019) );
no02f80 g565327 ( .a(n_3366), .b(n_2341), .o(n_4953) );
na03f80 g565328 ( .a(x_in_5_0), .b(n_2413), .c(x_in_5_1), .o(n_10937) );
oa12f80 g565329 ( .a(n_6504), .b(n_2618), .c(x_in_55_0), .o(n_4788) );
oa12f80 g565330 ( .a(n_7156), .b(n_2646), .c(x_in_23_0), .o(n_4790) );
no02f80 g565331 ( .a(n_2592), .b(n_3358), .o(n_5993) );
in01f80 g565332 ( .a(n_9167), .o(n_10489) );
oa12f80 g565333 ( .a(n_2753), .b(n_5365), .c(n_2747), .o(n_9167) );
ao12f80 g565334 ( .a(n_2209), .b(x_in_5_15), .c(x_in_4_13), .o(n_24032) );
na02f80 g565335 ( .a(n_2397), .b(n_3691), .o(n_5123) );
in01f80 g565336 ( .a(n_4952), .o(n_4775) );
ao12f80 g565337 ( .a(n_3872), .b(x_in_15_14), .c(x_in_15_13), .o(n_4952) );
in01f80 g565338 ( .a(n_9163), .o(n_10421) );
oa12f80 g565339 ( .a(n_3131), .b(n_5336), .c(n_3079), .o(n_9163) );
in01f80 g565340 ( .a(n_8650), .o(n_3378) );
na02f80 g565341 ( .a(n_3078), .b(n_2449), .o(n_8650) );
oa12f80 g565342 ( .a(n_7162), .b(n_2593), .c(x_in_15_0), .o(n_4785) );
na02f80 g565343 ( .a(n_2666), .b(n_3368), .o(n_5991) );
oa12f80 g565344 ( .a(n_7166), .b(n_2707), .c(x_in_13_0), .o(n_6296) );
oa12f80 g565345 ( .a(n_7153), .b(n_2660), .c(x_in_31_0), .o(n_4787) );
in01f80 g565346 ( .a(n_9157), .o(n_10455) );
oa12f80 g565347 ( .a(n_3293), .b(n_5373), .c(n_2721), .o(n_9157) );
in01f80 g565348 ( .a(n_9852), .o(n_6671) );
oa12f80 g565349 ( .a(n_2223), .b(x_in_13_3), .c(x_in_13_2), .o(n_9852) );
in01f80 g565350 ( .a(n_7396), .o(n_10529) );
oa12f80 g565351 ( .a(n_3076), .b(n_5430), .c(n_3075), .o(n_7396) );
in01f80 g565352 ( .a(n_3646), .o(n_2299) );
no03m80 g565353 ( .a(x_in_13_0), .b(x_in_13_2), .c(x_in_13_1), .o(n_3646) );
no02f80 g565354 ( .a(n_4432), .b(n_3803), .o(n_4253) );
in01f80 g565355 ( .a(n_4916), .o(n_4562) );
ao12f80 g565356 ( .a(n_7924), .b(x_in_49_4), .c(x_in_49_2), .o(n_4916) );
in01f80 g565357 ( .a(n_10385), .o(n_10387) );
oa12f80 g565358 ( .a(n_2781), .b(n_4946), .c(n_2780), .o(n_10385) );
in01f80 g565359 ( .a(n_2793), .o(n_5328) );
ao12f80 g565360 ( .a(n_4759), .b(x_in_13_4), .c(x_in_13_2), .o(n_2793) );
oa12f80 g565361 ( .a(n_3758), .b(x_in_9_4), .c(x_in_9_1), .o(n_4020) );
in01f80 g565362 ( .a(n_5852), .o(n_5851) );
oa12f80 g565363 ( .a(n_5034), .b(n_2230), .c(x_in_9_3), .o(n_5852) );
in01f80 g565364 ( .a(n_4288), .o(n_3441) );
oa12f80 g565365 ( .a(n_7076), .b(n_2445), .c(x_in_59_0), .o(n_4288) );
in01f80 g565366 ( .a(n_6507), .o(n_5808) );
no02f80 g565367 ( .a(n_3438), .b(n_3437), .o(n_6507) );
in01f80 g565368 ( .a(n_4965), .o(n_4394) );
ao12f80 g565369 ( .a(n_3870), .b(x_in_47_14), .c(x_in_47_13), .o(n_4965) );
in01f80 g565370 ( .a(n_4018), .o(n_3074) );
oa12f80 g565371 ( .a(n_4144), .b(x_in_25_3), .c(x_in_25_1), .o(n_4018) );
in01f80 g565372 ( .a(n_3439), .o(n_3440) );
ao12f80 g565373 ( .a(n_2817), .b(n_2419), .c(n_3241), .o(n_3439) );
ao12f80 g565374 ( .a(n_4013), .b(x_in_49_3), .c(x_in_49_1), .o(n_4016) );
oa12f80 g565375 ( .a(x_in_19_0), .b(x_in_19_2), .c(x_in_19_1), .o(n_2102) );
oa12f80 g565376 ( .a(n_7159), .b(n_2616), .c(x_in_47_0), .o(n_4789) );
in01f80 g565377 ( .a(n_9160), .o(n_10434) );
oa12f80 g565378 ( .a(n_3289), .b(n_5351), .c(n_2828), .o(n_9160) );
ao12f80 g565379 ( .a(n_4250), .b(x_in_29_3), .c(x_in_29_1), .o(n_4828) );
in01f80 g565380 ( .a(n_7598), .o(n_5385) );
oa12f80 g565381 ( .a(n_2599), .b(x_in_29_13), .c(x_in_29_11), .o(n_7598) );
in01f80 g565382 ( .a(n_9066), .o(n_4123) );
no02f80 g565383 ( .a(n_2370), .b(n_3334), .o(n_9066) );
in01f80 g565384 ( .a(n_5349), .o(n_4780) );
ao12f80 g565385 ( .a(n_3504), .b(x_in_63_14), .c(x_in_63_13), .o(n_5349) );
no02f80 g565386 ( .a(n_3629), .b(n_2560), .o(n_7639) );
ao12f80 g565387 ( .a(n_2148), .b(x_in_59_1), .c(x_in_59_0), .o(n_4771) );
in01f80 g565388 ( .a(n_8376), .o(n_3628) );
oa12f80 g565389 ( .a(n_3292), .b(n_2607), .c(x_in_39_0), .o(n_8376) );
oa12f80 g565390 ( .a(n_7237), .b(n_1042), .c(FE_OFN56_n_27012), .o(n_7356) );
oa12f80 g565391 ( .a(n_7237), .b(n_1821), .c(n_27449), .o(n_7233) );
oa12f80 g565392 ( .a(n_7237), .b(n_1418), .c(FE_OFN324_n_4860), .o(n_7238) );
oa12f80 g565393 ( .a(n_7239), .b(n_1330), .c(FE_OFN63_n_27012), .o(n_7240) );
oa12f80 g565394 ( .a(n_8188), .b(n_1801), .c(FE_OFN326_n_4860), .o(n_7243) );
oa12f80 g565395 ( .a(n_8204), .b(n_809), .c(FE_OFN136_n_27449), .o(n_7252) );
oa12f80 g565396 ( .a(FE_OFN144_n_7361), .b(n_1328), .c(FE_OFN78_n_27012), .o(n_7249) );
oa12f80 g565397 ( .a(n_7250), .b(n_1497), .c(FE_OFN68_n_27012), .o(n_7251) );
oa12f80 g565398 ( .a(n_4349), .b(n_1229), .c(FE_OFN1118_rst), .o(n_5775) );
oa12f80 g565399 ( .a(n_6481), .b(n_685), .c(FE_OFN1115_rst), .o(n_6482) );
oa12f80 g565400 ( .a(FE_OFN144_n_7361), .b(n_1652), .c(FE_OFN1121_rst), .o(n_5776) );
oa12f80 g565401 ( .a(n_7239), .b(n_1262), .c(FE_OFN1108_rst), .o(n_6480) );
oa12f80 g565402 ( .a(n_7254), .b(n_1499), .c(FE_OFN94_n_27449), .o(n_7255) );
oa12f80 g565403 ( .a(n_7250), .b(n_1210), .c(n_27449), .o(n_7257) );
oa12f80 g565404 ( .a(n_7261), .b(n_1435), .c(FE_OFN358_n_4860), .o(n_7256) );
oa12f80 g565405 ( .a(n_2799), .b(n_1074), .c(FE_OFN89_n_27449), .o(n_7258) );
oa12f80 g565406 ( .a(n_8204), .b(n_1422), .c(FE_OFN136_n_27449), .o(n_7259) );
oa12f80 g565407 ( .a(n_7261), .b(n_1427), .c(FE_OFN142_n_27449), .o(n_7262) );
oa12f80 g565408 ( .a(n_7283), .b(n_431), .c(FE_OFN100_n_27449), .o(n_7284) );
oa12f80 g565409 ( .a(n_4319), .b(n_300), .c(FE_OFN74_n_27012), .o(n_7293) );
oa12f80 g565410 ( .a(n_8198), .b(n_1684), .c(FE_OFN99_n_27449), .o(n_7306) );
oa12f80 g565411 ( .a(n_7330), .b(n_1728), .c(FE_OFN134_n_27449), .o(n_7331) );
oa12f80 g565412 ( .a(n_7283), .b(n_1938), .c(FE_OFN363_n_4860), .o(n_7345) );
oa12f80 g565413 ( .a(n_7330), .b(n_1747), .c(FE_OFN69_n_27012), .o(n_7344) );
oa12f80 g565414 ( .a(n_7347), .b(n_1665), .c(FE_OFN324_n_4860), .o(n_7348) );
oa12f80 g565415 ( .a(n_4307), .b(n_226), .c(FE_OFN358_n_4860), .o(n_7358) );
oa12f80 g565416 ( .a(n_7239), .b(n_1337), .c(FE_OFN336_n_4860), .o(n_7357) );
oa12f80 g565417 ( .a(FE_OFN144_n_7361), .b(n_1393), .c(FE_OFN141_n_27449), .o(n_7362) );
oa12f80 g565418 ( .a(n_7359), .b(n_1837), .c(FE_OFN64_n_27012), .o(n_7360) );
oa12f80 g565419 ( .a(n_4299), .b(n_1101), .c(FE_OFN104_n_27449), .o(n_7363) );
oa12f80 g565420 ( .a(n_7254), .b(n_1026), .c(FE_OFN94_n_27449), .o(n_7366) );
oa12f80 g565421 ( .a(n_4881), .b(n_1698), .c(FE_OFN133_n_27449), .o(n_7367) );
oa12f80 g565422 ( .a(n_2776), .b(n_26), .c(FE_OFN74_n_27012), .o(n_7368) );
oa12f80 g565423 ( .a(n_8188), .b(n_1219), .c(FE_OFN91_n_27449), .o(n_7369) );
oa12f80 g565424 ( .a(n_7359), .b(n_471), .c(n_29104), .o(n_7378) );
oa12f80 g565425 ( .a(n_4221), .b(n_1948), .c(FE_OFN1112_rst), .o(n_5785) );
oa12f80 g565426 ( .a(n_2821), .b(n_575), .c(FE_OFN126_n_27449), .o(n_7355) );
oa12f80 g565427 ( .a(n_8056), .b(n_360), .c(FE_OFN1112_rst), .o(n_5787) );
oa12f80 g565428 ( .a(n_4201), .b(n_102), .c(FE_OFN76_n_27012), .o(n_7375) );
oa12f80 g565429 ( .a(n_2859), .b(n_1970), .c(FE_OFN74_n_27012), .o(n_7374) );
oa12f80 g565430 ( .a(n_3348), .b(n_132), .c(FE_OFN138_n_27449), .o(n_7376) );
oa12f80 g565431 ( .a(n_4305), .b(n_645), .c(n_29261), .o(n_7377) );
oa12f80 g565432 ( .a(n_4295), .b(n_744), .c(FE_OFN94_n_27449), .o(n_7379) );
oa12f80 g565433 ( .a(n_2823), .b(n_101), .c(FE_OFN72_n_27012), .o(n_7388) );
oa12f80 g565434 ( .a(n_4194), .b(n_1541), .c(FE_OFN72_n_27012), .o(n_7392) );
oa12f80 g565435 ( .a(n_7406), .b(n_1334), .c(FE_OFN125_n_27449), .o(n_7393) );
oa12f80 g565436 ( .a(n_7261), .b(n_918), .c(FE_OFN1124_rst), .o(n_5952) );
oa12f80 g565437 ( .a(n_8198), .b(n_135), .c(FE_OFN1112_rst), .o(n_5971) );
oa12f80 g565438 ( .a(n_4311), .b(n_1234), .c(FE_OFN122_n_27449), .o(n_7354) );
oa12f80 g565439 ( .a(n_4233), .b(n_120), .c(FE_OFN74_n_27012), .o(n_7401) );
oa12f80 g565440 ( .a(n_7406), .b(n_325), .c(FE_OFN125_n_27449), .o(n_7407) );
oa12f80 g565441 ( .a(n_7406), .b(n_1344), .c(FE_OFN1112_rst), .o(n_6094) );
oa12f80 g565442 ( .a(n_8188), .b(n_1169), .c(n_29068), .o(n_5733) );
oa12f80 g565443 ( .a(n_6737), .b(n_494), .c(FE_OFN1108_rst), .o(n_6738) );
oa12f80 g565444 ( .a(n_7424), .b(n_1049), .c(FE_OFN347_n_4860), .o(n_7425) );
oa12f80 g565445 ( .a(n_7446), .b(n_1671), .c(FE_OFN335_n_4860), .o(n_7447) );
oa12f80 g565446 ( .a(n_7575), .b(n_648), .c(FE_OFN336_n_4860), .o(n_7576) );
oa12f80 g565447 ( .a(n_7575), .b(n_709), .c(FE_OFN336_n_4860), .o(n_7574) );
oa12f80 g565448 ( .a(n_7364), .b(n_128), .c(FE_OFN68_n_27012), .o(n_7588) );
oa12f80 g565449 ( .a(n_6737), .b(n_1223), .c(FE_OFN134_n_27449), .o(n_7628) );
oa12f80 g565450 ( .a(n_7347), .b(n_15), .c(n_27449), .o(n_7394) );
oa12f80 g565451 ( .a(n_7575), .b(n_1097), .c(n_29068), .o(n_6408) );
oa12f80 g565452 ( .a(n_4887), .b(n_1394), .c(FE_OFN122_n_27449), .o(n_7353) );
oa12f80 g565453 ( .a(n_4192), .b(n_143), .c(FE_OFN99_n_27449), .o(n_8005) );
oa12f80 g565454 ( .a(n_2986), .b(n_1522), .c(FE_OFN352_n_4860), .o(n_8002) );
oa12f80 g565455 ( .a(n_4315), .b(n_35), .c(FE_OFN357_n_4860), .o(n_8007) );
oa12f80 g565456 ( .a(FE_OFN282_n_7349), .b(n_765), .c(FE_OFN78_n_27012), .o(n_8018) );
oa12f80 g565457 ( .a(n_4301), .b(n_769), .c(FE_OFN364_n_4860), .o(n_8009) );
oa12f80 g565458 ( .a(n_4211), .b(n_705), .c(FE_OFN1182_rst), .o(n_6401) );
oa12f80 g565459 ( .a(n_4141), .b(n_737), .c(FE_OFN122_n_27449), .o(n_7352) );
oa12f80 g565460 ( .a(n_8198), .b(n_1280), .c(FE_OFN64_n_27012), .o(n_8199) );
oa12f80 g565461 ( .a(n_7446), .b(n_171), .c(FE_OFN335_n_4860), .o(n_8028) );
oa12f80 g565462 ( .a(n_4293), .b(n_1120), .c(FE_OFN95_n_27449), .o(n_8038) );
oa12f80 g565463 ( .a(n_8056), .b(n_1378), .c(FE_OFN125_n_27449), .o(n_8057) );
oa12f80 g565464 ( .a(n_6481), .b(n_1083), .c(FE_OFN324_n_4860), .o(n_8060) );
oa12f80 g565465 ( .a(n_8188), .b(n_1757), .c(FE_OFN1110_rst), .o(n_6428) );
oa12f80 g565466 ( .a(n_4297), .b(n_626), .c(FE_OFN68_n_27012), .o(n_7351) );
oa12f80 g565467 ( .a(n_8188), .b(n_702), .c(FE_OFN91_n_27449), .o(n_8189) );
oa12f80 g565468 ( .a(n_8056), .b(n_952), .c(FE_OFN1112_rst), .o(n_6430) );
oa12f80 g565469 ( .a(FE_OFN282_n_7349), .b(n_1758), .c(FE_OFN1119_rst), .o(n_6431) );
oa12f80 g565470 ( .a(FE_OFN282_n_7349), .b(n_222), .c(FE_OFN138_n_27449), .o(n_7350) );
oa12f80 g565471 ( .a(n_7364), .b(n_1812), .c(n_27449), .o(n_7365) );
oa12f80 g565472 ( .a(FE_OFN282_n_7349), .b(n_484), .c(n_27709), .o(n_7260) );
oa12f80 g565473 ( .a(n_2796), .b(n_1663), .c(FE_OFN1140_n_27012), .o(n_8203) );
oa12f80 g565474 ( .a(n_8204), .b(n_1887), .c(FE_OFN136_n_27449), .o(n_8205) );
in01f80 g565475 ( .a(n_5907), .o(n_4782) );
oa12f80 g565476 ( .a(n_2672), .b(x_in_53_2), .c(x_in_53_1), .o(n_5907) );
in01f80 g565477 ( .a(n_6285), .o(n_2843) );
oa12f80 g565478 ( .a(n_4099), .b(x_in_13_13), .c(x_in_13_11), .o(n_6285) );
oa12f80 g565479 ( .a(x_in_33_0), .b(x_in_33_2), .c(x_in_33_1), .o(n_2116) );
oa12f80 g565480 ( .a(n_2330), .b(x_in_59_3), .c(x_in_59_2), .o(n_2331) );
in01f80 g565481 ( .a(n_5850), .o(n_3612) );
na02f80 g565482 ( .a(n_2215), .b(n_3234), .o(n_5850) );
in01f80 g565483 ( .a(n_8541), .o(n_6359) );
ao12f80 g565484 ( .a(n_5723), .b(x_in_49_15), .c(x_in_49_12), .o(n_8541) );
ao12f80 g565485 ( .a(n_4317), .b(x_in_33_3), .c(x_in_33_1), .o(n_5215) );
in01f80 g565486 ( .a(n_9302), .o(n_8497) );
oa12f80 g565487 ( .a(n_2676), .b(x_in_35_14), .c(x_in_35_11), .o(n_9302) );
in01f80 g565488 ( .a(n_3496), .o(n_5923) );
ao12f80 g565489 ( .a(n_2763), .b(n_2762), .c(n_3193), .o(n_3496) );
in01f80 g565490 ( .a(n_7086), .o(n_3068) );
oa12f80 g565491 ( .a(n_3978), .b(x_in_35_13), .c(x_in_35_10), .o(n_7086) );
oa12f80 g565492 ( .a(n_5267), .b(x_in_57_3), .c(x_in_57_2), .o(n_2557) );
oa12f80 g565493 ( .a(n_2556), .b(x_in_25_5), .c(x_in_25_3), .o(n_5701) );
oa12f80 g565494 ( .a(x_in_49_10), .b(x_in_49_13), .c(x_in_49_12), .o(n_2237) );
in01f80 g565495 ( .a(n_3765), .o(n_3766) );
ao12f80 g565496 ( .a(n_2832), .b(n_23944), .c(n_3169), .o(n_3765) );
in01f80 g565497 ( .a(n_12606), .o(n_11320) );
oa12f80 g565498 ( .a(n_2555), .b(x_in_21_13), .c(x_in_21_10), .o(n_12606) );
oa12f80 g565499 ( .a(x_in_49_7), .b(x_in_49_10), .c(x_in_49_9), .o(n_2204) );
oa12f80 g565500 ( .a(x_in_49_6), .b(x_in_49_9), .c(x_in_49_8), .o(n_2284) );
oa12f80 g565501 ( .a(n_3354), .b(n_2539), .c(x_in_5_3), .o(n_2729) );
ao12f80 g565502 ( .a(n_7835), .b(x_in_61_3), .c(x_in_61_1), .o(n_7147) );
ao12f80 g565503 ( .a(n_2350), .b(n_5387), .c(n_2430), .o(n_2351) );
in01f80 g565504 ( .a(n_5853), .o(n_3611) );
na02f80 g565505 ( .a(n_2115), .b(n_2837), .o(n_5853) );
ao12f80 g565506 ( .a(n_2352), .b(x_in_19_12), .c(x_in_19_11), .o(n_8846) );
in01f80 g565507 ( .a(n_6750), .o(n_5443) );
ao12f80 g565508 ( .a(n_5838), .b(x_in_33_4), .c(x_in_33_2), .o(n_6750) );
oa12f80 g565509 ( .a(x_in_53_4), .b(x_in_53_7), .c(x_in_53_6), .o(n_2294) );
oa12f80 g565510 ( .a(x_in_53_6), .b(x_in_53_9), .c(x_in_53_8), .o(n_2081) );
oa12f80 g565511 ( .a(n_6945), .b(x_in_45_4), .c(x_in_45_1), .o(n_2740) );
oa12f80 g565512 ( .a(x_in_53_5), .b(x_in_53_8), .c(x_in_53_7), .o(n_2137) );
oa12f80 g565513 ( .a(x_in_53_7), .b(x_in_53_10), .c(x_in_53_9), .o(n_2203) );
oa12f80 g565514 ( .a(x_in_53_9), .b(x_in_53_12), .c(x_in_53_11), .o(n_2202) );
oa12f80 g565515 ( .a(x_in_53_8), .b(x_in_53_11), .c(x_in_53_10), .o(n_2069) );
oa12f80 g565516 ( .a(x_in_53_3), .b(x_in_53_6), .c(x_in_53_5), .o(n_2292) );
oa12f80 g565518 ( .a(n_2765), .b(x_in_59_5), .c(x_in_59_4), .o(n_2766) );
in01f80 g565519 ( .a(n_10053), .o(n_2754) );
oa12f80 g565520 ( .a(n_4707), .b(n_2554), .c(x_in_25_2), .o(n_10053) );
oa12f80 g565521 ( .a(x_in_53_10), .b(x_in_53_13), .c(x_in_53_12), .o(n_2079) );
in01f80 g565522 ( .a(n_7847), .o(n_3382) );
oa12f80 g565523 ( .a(n_2700), .b(n_2699), .c(x_in_7_0), .o(n_7847) );
ao12f80 g565524 ( .a(x_in_45_1), .b(n_2442), .c(x_in_45_0), .o(n_2328) );
ao12f80 g565526 ( .a(x_in_11_1), .b(n_5387), .c(n_2332), .o(n_2333) );
ao12f80 g565527 ( .a(n_5048), .b(n_4687), .c(x_in_17_0), .o(n_4772) );
in01f80 g565528 ( .a(n_4895), .o(n_5210) );
oa12f80 g565529 ( .a(n_5161), .b(n_8957), .c(x_in_9_9), .o(n_4895) );
ao12f80 g565530 ( .a(x_in_11_2), .b(n_2431), .c(n_2430), .o(n_2432) );
oa12f80 g565531 ( .a(n_4742), .b(x_in_51_5), .c(x_in_51_4), .o(n_3064) );
ao12f80 g565532 ( .a(x_in_27_1), .b(n_5679), .c(n_2478), .o(n_2553) );
ao12f80 g565533 ( .a(x_in_43_2), .b(n_2541), .c(n_3176), .o(n_2412) );
ao12f80 g565534 ( .a(n_2789), .b(x_in_21_3), .c(x_in_21_0), .o(n_2790) );
ao12f80 g565535 ( .a(x_in_43_1), .b(n_5293), .c(n_2349), .o(n_2552) );
ao12f80 g565536 ( .a(x_in_11_5), .b(n_5309), .c(n_5352), .o(n_2551) );
ao12f80 g565537 ( .a(n_3063), .b(n_5244), .c(x_in_19_15), .o(n_10048) );
in01f80 g565538 ( .a(n_10045), .o(n_2895) );
oa12f80 g565539 ( .a(n_2372), .b(n_3038), .c(x_in_53_2), .o(n_10045) );
ao12f80 g565540 ( .a(x_in_9_11), .b(n_8957), .c(x_in_9_15), .o(n_2441) );
oa12f80 g565541 ( .a(n_2611), .b(x_in_25_14), .c(x_in_25_12), .o(n_2820) );
ao12f80 g565542 ( .a(x_in_11_3), .b(n_5387), .c(n_5309), .o(n_2435) );
ao12f80 g565543 ( .a(n_2058), .b(x_in_61_6), .c(x_in_61_3), .o(n_4197) );
ao12f80 g565544 ( .a(x_in_27_2), .b(n_2421), .c(n_3747), .o(n_2402) );
in01f80 g565545 ( .a(n_10036), .o(n_2779) );
oa12f80 g565546 ( .a(n_3399), .b(n_2651), .c(x_in_53_4), .o(n_10036) );
in01f80 g565547 ( .a(n_10027), .o(n_3062) );
oa12f80 g565548 ( .a(n_3535), .b(n_2525), .c(x_in_53_5), .o(n_10027) );
in01f80 g565549 ( .a(n_10033), .o(n_2853) );
oa12f80 g565550 ( .a(n_3530), .b(n_2654), .c(x_in_53_6), .o(n_10033) );
ao12f80 g565551 ( .a(x_in_59_1), .b(n_5271), .c(n_2445), .o(n_2446) );
in01f80 g565552 ( .a(n_10030), .o(n_2836) );
oa12f80 g565553 ( .a(n_3963), .b(n_2653), .c(x_in_53_8), .o(n_10030) );
in01f80 g565554 ( .a(n_3607), .o(n_7813) );
oa12f80 g565555 ( .a(n_3516), .b(n_2409), .c(x_in_29_0), .o(n_3607) );
oa12f80 g565556 ( .a(n_6945), .b(n_2385), .c(x_in_45_0), .o(n_4891) );
in01f80 g565557 ( .a(n_10013), .o(n_3061) );
oa12f80 g565558 ( .a(n_3968), .b(n_2626), .c(x_in_53_3), .o(n_10013) );
in01f80 g565559 ( .a(n_10024), .o(n_3059) );
oa12f80 g565560 ( .a(n_3545), .b(n_2550), .c(x_in_53_7), .o(n_10024) );
in01f80 g565561 ( .a(n_10020), .o(n_2863) );
oa12f80 g565562 ( .a(n_4004), .b(n_4593), .c(x_in_25_3), .o(n_10020) );
ao12f80 g565563 ( .a(x_in_49_15), .b(n_2737), .c(x_in_49_14), .o(n_3966) );
in01f80 g565564 ( .a(n_10010), .o(n_2847) );
oa12f80 g565565 ( .a(n_3946), .b(n_3771), .c(x_in_25_4), .o(n_10010) );
ao12f80 g565566 ( .a(x_in_43_3), .b(n_5293), .c(n_5327), .o(n_2489) );
in01f80 g565567 ( .a(n_3488), .o(n_6576) );
oa12f80 g565568 ( .a(n_3387), .b(n_6726), .c(x_in_9_10), .o(n_3488) );
ao12f80 g565569 ( .a(n_4000), .b(n_8537), .c(x_in_29_12), .o(n_4706) );
in01f80 g565570 ( .a(n_5743), .o(n_5821) );
na02f80 g565571 ( .a(n_7757), .b(n_2246), .o(n_5743) );
in01f80 g565572 ( .a(n_10007), .o(n_3058) );
oa12f80 g565573 ( .a(n_3464), .b(n_3132), .c(x_in_25_5), .o(n_10007) );
in01f80 g565574 ( .a(n_4230), .o(n_4108) );
ao12f80 g565575 ( .a(n_4148), .b(n_7434), .c(x_in_21_0), .o(n_4230) );
oa12f80 g565576 ( .a(n_2504), .b(n_2214), .c(x_in_41_12), .o(n_7419) );
oa12f80 g565577 ( .a(n_3949), .b(n_5317), .c(x_in_25_10), .o(n_8747) );
ao12f80 g565578 ( .a(x_in_21_1), .b(n_7434), .c(n_8557), .o(n_2502) );
oa12f80 g565579 ( .a(n_3777), .b(x_in_35_5), .c(x_in_35_4), .o(n_2873) );
oa12f80 g565580 ( .a(n_3954), .b(n_2548), .c(x_in_53_10), .o(n_8360) );
in01f80 g565581 ( .a(n_10001), .o(n_3057) );
oa12f80 g565582 ( .a(n_3943), .b(n_3129), .c(x_in_25_6), .o(n_10001) );
oa12f80 g565583 ( .a(n_7434), .b(x_in_21_5), .c(x_in_21_3), .o(n_2199) );
in01f80 g565584 ( .a(n_9995), .o(n_2899) );
oa12f80 g565585 ( .a(n_3472), .b(n_2581), .c(x_in_25_7), .o(n_9995) );
in01f80 g565586 ( .a(n_9989), .o(n_2916) );
oa12f80 g565587 ( .a(n_3563), .b(n_2743), .c(x_in_25_8), .o(n_9989) );
in01f80 g565588 ( .a(n_9992), .o(n_2926) );
oa12f80 g565589 ( .a(n_3927), .b(n_3189), .c(x_in_25_9), .o(n_9992) );
in01f80 g565590 ( .a(n_5823), .o(n_8704) );
oa12f80 g565591 ( .a(n_4205), .b(n_2376), .c(x_in_9_13), .o(n_5823) );
in01f80 g565592 ( .a(n_4182), .o(n_3605) );
oa12f80 g565593 ( .a(n_2948), .b(n_2535), .c(x_in_25_3), .o(n_4182) );
in01f80 g565594 ( .a(n_3553), .o(n_6563) );
oa12f80 g565595 ( .a(n_4894), .b(n_2488), .c(x_in_9_8), .o(n_3553) );
in01f80 g565596 ( .a(n_9949), .o(n_3276) );
oa12f80 g565597 ( .a(n_4138), .b(n_2870), .c(x_in_53_9), .o(n_9949) );
ao12f80 g565598 ( .a(n_4725), .b(n_5825), .c(x_in_3_1), .o(n_2999) );
ao12f80 g565599 ( .a(n_4958), .b(n_2527), .c(x_in_45_11), .o(n_6216) );
ao12f80 g565600 ( .a(n_4659), .b(n_2528), .c(x_in_45_10), .o(n_6219) );
oa12f80 g565601 ( .a(x_in_35_12), .b(n_2652), .c(x_in_35_13), .o(n_9926) );
ao12f80 g565602 ( .a(n_2991), .b(n_2643), .c(x_in_9_14), .o(n_4206) );
in01f80 g565603 ( .a(n_5892), .o(n_5891) );
oa12f80 g565604 ( .a(n_3773), .b(n_3736), .c(x_in_29_13), .o(n_5892) );
oa12f80 g565605 ( .a(n_2680), .b(n_4057), .c(x_in_19_15), .o(n_5146) );
ao12f80 g565606 ( .a(n_4639), .b(n_3011), .c(x_in_37_0), .o(n_4655) );
in01f80 g565607 ( .a(n_8561), .o(n_8546) );
oa12f80 g565608 ( .a(n_2950), .b(n_4825), .c(x_in_53_0), .o(n_8561) );
ao12f80 g565609 ( .a(n_3022), .b(n_7765), .c(x_in_19_13), .o(n_4700) );
in01f80 g565610 ( .a(n_5826), .o(n_5830) );
ao12f80 g565611 ( .a(n_7748), .b(n_5931), .c(x_in_3_2), .o(n_5826) );
ao12f80 g565612 ( .a(n_2842), .b(n_5418), .c(x_in_17_14), .o(n_5489) );
in01f80 g565613 ( .a(n_3601), .o(n_6577) );
oa12f80 g565614 ( .a(n_4645), .b(n_2289), .c(x_in_9_4), .o(n_3601) );
in01f80 g565615 ( .a(n_9338), .o(n_3631) );
oa12f80 g565616 ( .a(n_8693), .b(n_5872), .c(x_in_21_14), .o(n_9338) );
in01f80 g565617 ( .a(n_5925), .o(n_3630) );
oa12f80 g565618 ( .a(n_3827), .b(n_3077), .c(x_in_13_13), .o(n_5925) );
in01f80 g565619 ( .a(n_12197), .o(n_11201) );
no02f80 g565620 ( .a(n_7734), .b(n_2232), .o(n_12197) );
in01f80 g565621 ( .a(n_7499), .o(n_7498) );
oa12f80 g565622 ( .a(n_3025), .b(n_5926), .c(x_in_13_11), .o(n_7499) );
oa12f80 g565623 ( .a(n_5271), .b(n_3260), .c(x_in_59_2), .o(n_5268) );
in01f80 g565624 ( .a(n_5859), .o(n_5858) );
ao12f80 g565625 ( .a(n_3108), .b(n_5537), .c(x_in_19_11), .o(n_5859) );
oa12f80 g565626 ( .a(n_3980), .b(n_5317), .c(x_in_25_15), .o(n_3600) );
in01f80 g565627 ( .a(n_7519), .o(n_5795) );
ao12f80 g565628 ( .a(n_6935), .b(n_5415), .c(x_in_17_14), .o(n_7519) );
oa12f80 g565629 ( .a(n_3054), .b(n_5679), .c(x_in_27_1), .o(n_3055) );
in01f80 g565630 ( .a(n_7556), .o(n_5140) );
ao12f80 g565631 ( .a(n_6932), .b(n_5247), .c(x_in_3_14), .o(n_7556) );
oa12f80 g565632 ( .a(n_4636), .b(n_2588), .c(x_in_49_4), .o(n_4160) );
in01f80 g565633 ( .a(n_8477), .o(n_7581) );
na02f80 g565634 ( .a(n_4903), .b(n_2125), .o(n_8477) );
in01f80 g565635 ( .a(n_6416), .o(n_5970) );
oa12f80 g565636 ( .a(n_3027), .b(n_2737), .c(x_in_49_11), .o(n_6416) );
in01f80 g565637 ( .a(n_9287), .o(n_5135) );
oa12f80 g565638 ( .a(n_6921), .b(n_2752), .c(x_in_35_12), .o(n_9287) );
in01f80 g565639 ( .a(n_4646), .o(n_5212) );
oa12f80 g565640 ( .a(n_4980), .b(n_2060), .c(x_in_9_5), .o(n_4646) );
in01f80 g565641 ( .a(n_3580), .o(n_3581) );
oa12f80 g565642 ( .a(n_2808), .b(n_2673), .c(x_in_13_11), .o(n_3580) );
in01f80 g565643 ( .a(n_4251), .o(n_3599) );
oa12f80 g565644 ( .a(n_5790), .b(n_3724), .c(x_in_29_2), .o(n_4251) );
oa12f80 g565645 ( .a(n_2563), .b(n_2583), .c(x_in_41_6), .o(n_5482) );
ao12f80 g565646 ( .a(n_4027), .b(n_2597), .c(x_in_29_11), .o(n_4183) );
in01f80 g565647 ( .a(n_5889), .o(n_5476) );
ao12f80 g565648 ( .a(n_3845), .b(n_2875), .c(x_in_29_12), .o(n_5889) );
in01f80 g565649 ( .a(n_4833), .o(n_5191) );
no02f80 g565650 ( .a(n_2857), .b(n_2128), .o(n_4833) );
in01f80 g565651 ( .a(n_5436), .o(n_4960) );
no02f80 g565652 ( .a(n_9095), .b(n_2168), .o(n_5436) );
oa12f80 g565653 ( .a(n_2663), .b(n_2636), .c(x_in_33_2), .o(n_4052) );
in01f80 g565654 ( .a(n_5956), .o(n_4124) );
oa12f80 g565655 ( .a(n_3305), .b(n_5905), .c(x_in_3_11), .o(n_5956) );
in01f80 g565656 ( .a(n_7475), .o(n_7474) );
oa12f80 g565657 ( .a(n_2880), .b(n_9608), .c(x_in_41_11), .o(n_7475) );
in01f80 g565658 ( .a(n_5893), .o(n_4024) );
ao12f80 g565659 ( .a(n_3239), .b(n_5939), .c(x_in_19_6), .o(n_5893) );
in01f80 g565660 ( .a(n_5855), .o(n_3598) );
na02f80 g565661 ( .a(n_4213), .b(n_2075), .o(n_5855) );
oa12f80 g565662 ( .a(n_2334), .b(n_5415), .c(x_in_17_11), .o(n_3051) );
oa12f80 g565663 ( .a(n_3050), .b(n_10477), .c(x_in_17_10), .o(n_4998) );
ao12f80 g565664 ( .a(n_4258), .b(n_4738), .c(x_in_31_2), .o(n_3049) );
ao12f80 g565665 ( .a(n_4582), .b(n_4737), .c(x_in_47_2), .o(n_3048) );
in01f80 g565666 ( .a(n_5936), .o(n_5937) );
oa12f80 g565667 ( .a(n_3047), .b(n_5244), .c(x_in_19_10), .o(n_5936) );
in01f80 g565668 ( .a(n_6213), .o(n_4959) );
oa12f80 g565669 ( .a(n_4997), .b(n_10486), .c(x_in_45_9), .o(n_6213) );
oa12f80 g565670 ( .a(n_3046), .b(n_5360), .c(x_in_17_5), .o(n_5478) );
in01f80 g565671 ( .a(n_5727), .o(n_5728) );
oa12f80 g565672 ( .a(n_7380), .b(n_5931), .c(x_in_3_6), .o(n_5727) );
ao12f80 g565673 ( .a(n_2530), .b(n_2870), .c(x_in_53_15), .o(n_6573) );
in01f80 g565674 ( .a(n_4634), .o(n_3597) );
oa12f80 g565675 ( .a(n_4642), .b(n_3186), .c(x_in_49_9), .o(n_4634) );
in01f80 g565676 ( .a(n_4347), .o(n_5163) );
ao12f80 g565677 ( .a(n_6766), .b(n_5849), .c(x_in_37_10), .o(n_4347) );
ao12f80 g565678 ( .a(n_3045), .b(n_2438), .c(x_in_45_8), .o(n_6209) );
ao12f80 g565679 ( .a(n_4220), .b(n_2442), .c(x_in_45_7), .o(n_6437) );
in01f80 g565680 ( .a(n_10224), .o(n_10226) );
no02f80 g565681 ( .a(n_4857), .b(n_2071), .o(n_10224) );
in01f80 g565682 ( .a(n_5915), .o(n_5989) );
no02f80 g565683 ( .a(n_2791), .b(n_2282), .o(n_5915) );
ao12f80 g565684 ( .a(n_3879), .b(n_3187), .c(x_in_49_12), .o(n_4643) );
in01f80 g565685 ( .a(n_5873), .o(n_5087) );
oa12f80 g565686 ( .a(n_3044), .b(n_3043), .c(x_in_21_13), .o(n_5873) );
in01f80 g565687 ( .a(n_4739), .o(n_5831) );
ao12f80 g565688 ( .a(n_10793), .b(n_3560), .c(x_in_57_14), .o(n_4739) );
in01f80 g565689 ( .a(n_5740), .o(n_3596) );
na02f80 g565690 ( .a(n_8303), .b(n_2253), .o(n_5740) );
oa12f80 g565691 ( .a(n_4172), .b(n_8537), .c(x_in_29_8), .o(n_4236) );
in01f80 g565692 ( .a(n_10220), .o(n_10222) );
no02f80 g565693 ( .a(n_2095), .b(n_3042), .o(n_10220) );
ao12f80 g565694 ( .a(n_4146), .b(n_2513), .c(x_in_45_9), .o(n_6204) );
in01f80 g565695 ( .a(n_5885), .o(n_5886) );
ao12f80 g565696 ( .a(n_8305), .b(n_4180), .c(x_in_37_9), .o(n_5885) );
in01f80 g565697 ( .a(n_8295), .o(n_8297) );
na02f80 g565698 ( .a(n_2898), .b(n_2082), .o(n_8295) );
in01f80 g565699 ( .a(n_5751), .o(n_3595) );
oa12f80 g565700 ( .a(n_7710), .b(n_5860), .c(x_in_21_10), .o(n_5751) );
in01f80 g565701 ( .a(n_4341), .o(n_5837) );
no02f80 g565702 ( .a(n_3041), .b(n_2118), .o(n_4341) );
in01f80 g565703 ( .a(n_5749), .o(n_5750) );
ao12f80 g565704 ( .a(n_3040), .b(n_5881), .c(x_in_37_6), .o(n_5749) );
in01f80 g565705 ( .a(n_5639), .o(n_4109) );
oa12f80 g565706 ( .a(n_3039), .b(n_9610), .c(x_in_41_7), .o(n_5639) );
oa12f80 g565707 ( .a(n_2387), .b(n_7915), .c(x_in_41_11), .o(n_5645) );
oa12f80 g565708 ( .a(n_3326), .b(n_9329), .c(x_in_41_10), .o(n_5685) );
in01f80 g565709 ( .a(n_10218), .o(n_10216) );
oa12f80 g565710 ( .a(n_5633), .b(n_3038), .c(x_in_53_5), .o(n_10218) );
in01f80 g565711 ( .a(n_5922), .o(n_3430) );
oa12f80 g565712 ( .a(n_7687), .b(n_8557), .c(x_in_21_6), .o(n_5922) );
in01f80 g565713 ( .a(n_5752), .o(n_5753) );
ao12f80 g565714 ( .a(n_7693), .b(n_5872), .c(x_in_21_9), .o(n_5752) );
in01f80 g565715 ( .a(n_5861), .o(n_5887) );
ao12f80 g565716 ( .a(n_3037), .b(n_3036), .c(x_in_21_5), .o(n_5861) );
in01f80 g565717 ( .a(n_10212), .o(n_10214) );
na02f80 g565718 ( .a(n_6374), .b(n_2108), .o(n_10212) );
in01f80 g565719 ( .a(n_4554), .o(n_3475) );
ao12f80 g565720 ( .a(n_4159), .b(n_3238), .c(x_in_49_5), .o(n_4554) );
in01f80 g565721 ( .a(n_3593), .o(n_5468) );
oa12f80 g565722 ( .a(n_2841), .b(n_9651), .c(x_in_17_4), .o(n_3593) );
in01f80 g565723 ( .a(n_5121), .o(n_4367) );
ao12f80 g565724 ( .a(n_3592), .b(n_3591), .c(x_in_29_5), .o(n_5121) );
ao12f80 g565725 ( .a(n_4226), .b(n_3035), .c(x_in_29_9), .o(n_4615) );
in01f80 g565726 ( .a(n_3589), .o(n_5464) );
oa12f80 g565727 ( .a(n_3336), .b(n_9654), .c(x_in_17_6), .o(n_3589) );
ao12f80 g565728 ( .a(n_5789), .b(n_3724), .c(x_in_29_6), .o(n_5116) );
in01f80 g565729 ( .a(n_5932), .o(n_5933) );
ao12f80 g565730 ( .a(n_3034), .b(n_3174), .c(x_in_19_7), .o(n_5932) );
oa12f80 g565731 ( .a(n_7683), .b(n_5869), .c(x_in_21_12), .o(n_5943) );
in01f80 g565732 ( .a(n_5874), .o(n_3588) );
oa12f80 g565733 ( .a(n_7697), .b(n_5963), .c(x_in_3_7), .o(n_5874) );
in01f80 g565734 ( .a(n_5411), .o(n_5062) );
no02f80 g565735 ( .a(n_2109), .b(n_7681), .o(n_5411) );
in01f80 g565736 ( .a(n_5880), .o(n_4053) );
oa12f80 g565737 ( .a(n_7679), .b(n_5742), .c(x_in_37_7), .o(n_5880) );
in01f80 g565738 ( .a(n_5882), .o(n_5883) );
ao12f80 g565739 ( .a(n_3095), .b(n_5962), .c(x_in_37_7), .o(n_5882) );
oa12f80 g565740 ( .a(n_3200), .b(n_5415), .c(x_in_17_9), .o(n_5611) );
ao12f80 g565741 ( .a(n_7675), .b(n_2548), .c(x_in_53_14), .o(n_6200) );
in01f80 g565742 ( .a(n_3586), .o(n_5460) );
oa12f80 g565743 ( .a(n_2830), .b(n_5418), .c(x_in_17_8), .o(n_3586) );
oa22f80 g565744 ( .a(n_1711), .b(FE_OFN133_n_27449), .c(n_4280), .d(n_8513), .o(n_7342) );
oa22f80 g565745 ( .a(n_0), .b(FE_OFN108_n_27449), .c(FE_OFN416_n_28303), .d(n_7340), .o(n_7341) );
oa22f80 g565746 ( .a(n_1009), .b(FE_OFN94_n_27449), .c(FE_OFN307_n_3069), .d(n_7338), .o(n_7339) );
oa12f80 g565747 ( .a(n_2301), .b(n_3191), .c(x_in_49_7), .o(n_4606) );
oa22f80 g565748 ( .a(n_435), .b(FE_OFN77_n_27012), .c(FE_OFN296_n_3069), .d(n_7336), .o(n_7337) );
oa22f80 g565749 ( .a(n_922), .b(FE_OFN355_n_4860), .c(FE_OFN260_n_4280), .d(n_7334), .o(n_7335) );
oa22f80 g565750 ( .a(n_970), .b(FE_OFN1119_rst), .c(FE_OFN404_n_28303), .d(n_11041), .o(n_6456) );
oa22f80 g565751 ( .a(n_978), .b(FE_OFN357_n_4860), .c(FE_OFN234_n_4162), .d(n_5679), .o(n_7223) );
in01f80 g565752 ( .a(n_3909), .o(n_2730) );
oa12f80 g565753 ( .a(n_2029), .b(x_in_57_2), .c(x_in_57_0), .o(n_3909) );
in01f80 g565754 ( .a(n_3562), .o(n_5774) );
ao12f80 g565755 ( .a(n_3859), .b(n_7216), .c(x_in_45_14), .o(n_3562) );
in01f80 g565756 ( .a(n_11168), .o(n_8502) );
no02f80 g565757 ( .a(n_2279), .b(n_6382), .o(n_11168) );
oa22f80 g565758 ( .a(n_1744), .b(FE_OFN104_n_27449), .c(FE_OFN258_n_4280), .d(n_7332), .o(n_7333) );
in01f80 g565759 ( .a(n_5877), .o(n_5876) );
ao12f80 g565760 ( .a(n_3033), .b(n_5940), .c(x_in_19_9), .o(n_5877) );
in01f80 g565761 ( .a(n_3582), .o(n_6571) );
oa12f80 g565762 ( .a(n_4608), .b(n_2248), .c(x_in_9_6), .o(n_3582) );
oa22f80 g565763 ( .a(n_468), .b(FE_OFN336_n_4860), .c(FE_OFN1167_n_4162), .d(n_5272), .o(n_7329) );
oa22f80 g565764 ( .a(n_60), .b(FE_OFN331_n_4860), .c(FE_OFN404_n_28303), .d(n_5677), .o(n_7328) );
oa22f80 g565765 ( .a(n_768), .b(FE_OFN78_n_27012), .c(FE_OFN294_n_3069), .d(n_7417), .o(n_7418) );
oa22f80 g565766 ( .a(x_in_32_15), .b(x_in_33_15), .c(n_2538), .d(n_1383), .o(n_29187) );
in01f80 g565767 ( .a(n_11148), .o(n_8503) );
no02f80 g565768 ( .a(n_2070), .b(n_6369), .o(n_11148) );
oa22f80 g565769 ( .a(n_466), .b(FE_OFN101_n_27449), .c(FE_OFN230_n_4162), .d(n_3742), .o(n_7327) );
oa22f80 g565770 ( .a(n_857), .b(FE_OFN63_n_27012), .c(FE_OFN400_n_28303), .d(n_7325), .o(n_7326) );
ao12f80 g565771 ( .a(n_5107), .b(n_5095), .c(x_in_49_7), .o(n_4638) );
oa22f80 g565772 ( .a(n_1921), .b(FE_OFN1119_rst), .c(FE_OFN203_n_28771), .d(n_3075), .o(n_6498) );
oa22f80 g565773 ( .a(n_146), .b(n_29068), .c(n_29664), .d(n_6496), .o(n_6497) );
in01f80 g565774 ( .a(n_5930), .o(n_3381) );
oa12f80 g565775 ( .a(n_3031), .b(n_5825), .c(x_in_3_5), .o(n_5930) );
oa22f80 g565776 ( .a(n_320), .b(FE_OFN74_n_27012), .c(FE_OFN294_n_3069), .d(n_7323), .o(n_7324) );
oa22f80 g565777 ( .a(n_1780), .b(FE_OFN133_n_27449), .c(n_4280), .d(n_7229), .o(n_7230) );
oa22f80 g565778 ( .a(n_1196), .b(FE_OFN91_n_27449), .c(FE_OFN308_n_3069), .d(n_5501), .o(n_7253) );
ao22s80 g565779 ( .a(n_2413), .b(n_742), .c(x_in_5_2), .d(x_in_5_0), .o(n_3542) );
oa22f80 g565780 ( .a(n_346), .b(FE_OFN1108_rst), .c(FE_OFN256_n_4280), .d(n_6494), .o(n_6495) );
in01f80 g565781 ( .a(n_4609), .o(n_5218) );
oa12f80 g565782 ( .a(n_5130), .b(n_2285), .c(x_in_9_7), .o(n_4609) );
oa22f80 g565783 ( .a(n_1191), .b(FE_OFN324_n_4860), .c(FE_OFN293_n_3069), .d(n_2828), .o(n_7322) );
oa22f80 g565784 ( .a(n_580), .b(FE_OFN102_n_27449), .c(FE_OFN230_n_4162), .d(n_7320), .o(n_7321) );
oa22f80 g565785 ( .a(n_1839), .b(FE_OFN96_n_27449), .c(n_27933), .d(n_3107), .o(n_7319) );
oa22f80 g565786 ( .a(n_42), .b(FE_OFN56_n_27012), .c(FE_OFN184_n_29402), .d(n_7317), .o(n_7318) );
oa22f80 g565787 ( .a(n_285), .b(FE_OFN352_n_4860), .c(FE_OFN230_n_4162), .d(n_7315), .o(n_7316) );
oa22f80 g565788 ( .a(n_1402), .b(FE_OFN125_n_27449), .c(FE_OFN306_n_3069), .d(n_2780), .o(n_7314) );
oa22f80 g565789 ( .a(n_75), .b(n_27449), .c(n_22960), .d(n_7311), .o(n_7312) );
oa22f80 g565790 ( .a(n_1799), .b(FE_OFN102_n_27449), .c(FE_OFN402_n_28303), .d(n_5256), .o(n_7310) );
oa22f80 g565791 ( .a(n_525), .b(n_27449), .c(n_28597), .d(n_7308), .o(n_7309) );
ao12f80 g565792 ( .a(n_1994), .b(x_in_57_3), .c(x_in_57_1), .o(n_3618) );
oa22f80 g565793 ( .a(x_in_57_15), .b(x_in_56_15), .c(n_3641), .d(n_818), .o(n_28813) );
oa22f80 g565794 ( .a(n_1591), .b(FE_OFN60_n_27012), .c(FE_OFN267_n_4280), .d(n_5327), .o(n_7307) );
in01f80 g565795 ( .a(n_5953), .o(n_5959) );
ao12f80 g565796 ( .a(n_2801), .b(n_5247), .c(x_in_3_10), .o(n_5953) );
oa22f80 g565797 ( .a(n_1008), .b(FE_OFN102_n_27449), .c(FE_OFN296_n_3069), .d(n_7304), .o(n_7305) );
oa22f80 g565798 ( .a(n_1247), .b(FE_OFN60_n_27012), .c(FE_OFN267_n_4280), .d(n_5519), .o(n_7303) );
oa22f80 g565799 ( .a(n_1150), .b(FE_OFN1112_rst), .c(FE_OFN307_n_3069), .d(n_6492), .o(n_6493) );
oa22f80 g565800 ( .a(n_1548), .b(FE_OFN1110_rst), .c(FE_OFN267_n_4280), .d(n_3176), .o(n_6491) );
oa22f80 g565801 ( .a(x_in_25_15), .b(x_in_24_15), .c(n_2546), .d(n_2545), .o(n_28801) );
oa22f80 g565802 ( .a(n_920), .b(FE_OFN136_n_27449), .c(FE_OFN299_n_3069), .d(n_6689), .o(n_7302) );
oa22f80 g565803 ( .a(n_1151), .b(FE_OFN94_n_27449), .c(FE_OFN306_n_3069), .d(n_2747), .o(n_7234) );
oa22f80 g565804 ( .a(n_870), .b(FE_OFN94_n_27449), .c(FE_OFN264_n_4280), .d(n_3445), .o(n_7235) );
oa22f80 g565805 ( .a(n_1204), .b(FE_OFN72_n_27012), .c(FE_OFN236_n_4162), .d(n_6683), .o(n_7236) );
oa22f80 g565806 ( .a(n_1468), .b(FE_OFN64_n_27012), .c(n_26454), .d(n_7241), .o(n_7242) );
oa22f80 g565807 ( .a(n_807), .b(FE_OFN64_n_27012), .c(FE_OFN409_n_28303), .d(n_11034), .o(n_7244) );
oa22f80 g565808 ( .a(n_1322), .b(FE_OFN94_n_27449), .c(FE_OFN307_n_3069), .d(n_7245), .o(n_7246) );
oa22f80 g565809 ( .a(n_7), .b(FE_OFN94_n_27449), .c(FE_OFN236_n_4162), .d(n_7247), .o(n_7248) );
oa22f80 g565810 ( .a(n_1233), .b(FE_OFN1112_rst), .c(FE_OFN409_n_28303), .d(n_2558), .o(n_6490) );
oa22f80 g565811 ( .a(n_1352), .b(FE_OFN1119_rst), .c(FE_OFN404_n_28303), .d(n_6488), .o(n_6489) );
oa22f80 g565812 ( .a(n_410), .b(FE_OFN1112_rst), .c(FE_OFN260_n_4280), .d(n_3482), .o(n_6499) );
oa12f80 g565813 ( .a(n_2025), .b(x_in_16_15), .c(x_in_17_15), .o(n_29201) );
in01f80 g565814 ( .a(n_5732), .o(n_3575) );
oa12f80 g565815 ( .a(n_2997), .b(n_5757), .c(x_in_3_9), .o(n_5732) );
in01f80 g565816 ( .a(n_11166), .o(n_8485) );
no02f80 g565817 ( .a(n_2085), .b(n_6362), .o(n_11166) );
oa22f80 g565818 ( .a(n_1216), .b(FE_OFN102_n_27449), .c(FE_OFN256_n_4280), .d(n_5968), .o(n_7301) );
in01f80 g565819 ( .a(n_5942), .o(n_5941) );
oa12f80 g565820 ( .a(n_3021), .b(n_3020), .c(x_in_19_8), .o(n_5942) );
oa12f80 g565821 ( .a(n_3026), .b(n_5554), .c(x_in_19_6), .o(n_5934) );
oa22f80 g565822 ( .a(n_1915), .b(FE_OFN56_n_27012), .c(n_29664), .d(n_3739), .o(n_7300) );
oa22f80 g565823 ( .a(n_98), .b(FE_OFN63_n_27012), .c(FE_OFN266_n_4280), .d(n_11698), .o(n_7313) );
oa22f80 g565824 ( .a(n_891), .b(n_27449), .c(n_22019), .d(n_7298), .o(n_7299) );
oa22f80 g565825 ( .a(n_656), .b(FE_OFN68_n_27012), .c(FE_OFN198_n_29637), .d(n_2606), .o(n_7343) );
oa12f80 g565826 ( .a(n_2806), .b(n_5881), .c(x_in_37_10), .o(n_5409) );
oa22f80 g565827 ( .a(n_1946), .b(FE_OFN95_n_27449), .c(FE_OFN292_n_3069), .d(n_2537), .o(n_7346) );
oa22f80 g565828 ( .a(n_1973), .b(FE_OFN100_n_27449), .c(FE_OFN299_n_3069), .d(n_7296), .o(n_7297) );
oa22f80 g565829 ( .a(n_1087), .b(FE_OFN68_n_27012), .c(n_28303), .d(n_11696), .o(n_7295) );
oa12f80 g565830 ( .a(n_3345), .b(n_5359), .c(x_in_17_7), .o(n_5616) );
oa22f80 g565831 ( .a(n_178), .b(FE_OFN1182_rst), .c(n_26184), .d(n_6753), .o(n_6487) );
oa22f80 g565832 ( .a(n_252), .b(FE_OFN1108_rst), .c(FE_OFN303_n_3069), .d(n_6500), .o(n_6501) );
oa22f80 g565833 ( .a(n_1809), .b(FE_OFN1117_rst), .c(FE_OFN292_n_3069), .d(n_3079), .o(n_6486) );
in01f80 g565834 ( .a(n_5756), .o(n_5758) );
oa12f80 g565835 ( .a(n_7645), .b(n_5524), .c(x_in_3_10), .o(n_5756) );
in01f80 g565836 ( .a(n_3573), .o(n_5109) );
ao12f80 g565837 ( .a(n_5125), .b(n_3188), .c(x_in_49_10), .o(n_3573) );
oa22f80 g565838 ( .a(n_958), .b(FE_OFN76_n_27012), .c(FE_OFN307_n_3069), .d(n_11037), .o(n_7294) );
oa22f80 g565839 ( .a(n_376), .b(FE_OFN345_n_4860), .c(FE_OFN266_n_4280), .d(n_7291), .o(n_7292) );
oa22f80 g565840 ( .a(n_1365), .b(FE_OFN355_n_4860), .c(FE_OFN260_n_4280), .d(n_6687), .o(n_7370) );
oa22f80 g565841 ( .a(n_841), .b(FE_OFN133_n_27449), .c(FE_OFN404_n_28303), .d(n_7402), .o(n_7403) );
oa22f80 g565842 ( .a(n_1582), .b(FE_OFN347_n_4860), .c(FE_OFN300_n_3069), .d(n_2036), .o(n_7371) );
oa22f80 g565843 ( .a(n_1796), .b(FE_OFN63_n_27012), .c(n_23291), .d(n_7289), .o(n_7290) );
oa12f80 g565844 ( .a(n_2013), .b(x_in_0_15), .c(x_in_1_15), .o(n_26552) );
oa22f80 g565845 ( .a(n_1356), .b(FE_OFN355_n_4860), .c(FE_OFN307_n_3069), .d(n_2574), .o(n_7372) );
oa22f80 g565846 ( .a(n_1263), .b(FE_OFN101_n_27449), .c(n_4280), .d(n_7287), .o(n_7288) );
ao12f80 g565847 ( .a(n_4089), .b(n_3390), .c(x_in_29_8), .o(n_4598) );
in01f80 g565848 ( .a(n_5862), .o(n_5864) );
ao12f80 g565849 ( .a(n_3024), .b(n_5216), .c(x_in_9_5), .o(n_5862) );
oa22f80 g565850 ( .a(n_12), .b(FE_OFN108_n_27449), .c(FE_OFN416_n_28303), .d(n_7285), .o(n_7286) );
oa22f80 g565851 ( .a(x_in_9_15), .b(x_in_8_15), .c(n_2643), .d(n_1942), .o(n_28765) );
oa22f80 g565852 ( .a(n_1865), .b(FE_OFN1109_rst), .c(FE_OFN404_n_28303), .d(n_5680), .o(n_6485) );
oa22f80 g565853 ( .a(n_1662), .b(FE_OFN104_n_27449), .c(FE_OFN230_n_4162), .d(n_11040), .o(n_7282) );
oa22f80 g565854 ( .a(n_388), .b(FE_OFN122_n_27449), .c(FE_OFN311_n_3069), .d(n_8522), .o(n_7281) );
oa12f80 g565855 ( .a(n_3019), .b(n_9612), .c(x_in_41_9), .o(n_5642) );
oa12f80 g565856 ( .a(n_3252), .b(n_9327), .c(x_in_41_8), .o(n_5916) );
oa22f80 g565857 ( .a(n_1892), .b(n_29266), .c(n_27933), .d(n_6483), .o(n_6484) );
in01f80 g565858 ( .a(n_5111), .o(n_4852) );
oa12f80 g565859 ( .a(n_4336), .b(n_3035), .c(x_in_29_5), .o(n_5111) );
oa22f80 g565860 ( .a(n_1417), .b(FE_OFN68_n_27012), .c(FE_OFN258_n_4280), .d(n_6685), .o(n_7280) );
oa22f80 g565861 ( .a(n_457), .b(FE_OFN138_n_27449), .c(FE_OFN297_n_3069), .d(n_7278), .o(n_7279) );
in01f80 g565862 ( .a(n_5870), .o(n_5903) );
ao12f80 g565863 ( .a(n_3211), .b(n_3887), .c(x_in_21_7), .o(n_5870) );
in01f80 g565864 ( .a(n_5039), .o(n_3018) );
oa22f80 g565865 ( .a(x_in_39_2), .b(x_in_39_1), .c(n_2037), .d(n_2607), .o(n_5039) );
ao22s80 g565866 ( .a(n_23944), .b(n_2608), .c(x_in_4_15), .d(x_in_5_15), .o(n_25702) );
oa22f80 g565867 ( .a(n_541), .b(FE_OFN101_n_27449), .c(n_16028), .d(n_3747), .o(n_7277) );
oa22f80 g565868 ( .a(n_1974), .b(FE_OFN63_n_27012), .c(FE_OFN235_n_4162), .d(n_8133), .o(n_8134) );
oa22f80 g565869 ( .a(n_1034), .b(FE_OFN102_n_27449), .c(FE_OFN256_n_4280), .d(n_8165), .o(n_8166) );
oa22f80 g565870 ( .a(n_1458), .b(FE_OFN122_n_27449), .c(FE_OFN303_n_3069), .d(n_8200), .o(n_8201) );
oa22f80 g565871 ( .a(n_1732), .b(FE_OFN129_n_27449), .c(n_29496), .d(n_2721), .o(n_8202) );
in01f80 g565872 ( .a(n_4599), .o(n_3495) );
oa12f80 g565873 ( .a(n_2883), .b(n_3188), .c(x_in_49_6), .o(n_4599) );
oa22f80 g565874 ( .a(n_980), .b(FE_OFN350_n_4860), .c(FE_OFN253_n_4280), .d(n_3744), .o(n_7276) );
oa22f80 g565875 ( .a(n_1597), .b(FE_OFN68_n_27012), .c(n_29698), .d(n_8206), .o(n_8207) );
oa22f80 g565876 ( .a(n_931), .b(FE_OFN1118_rst), .c(FE_OFN219_n_23315), .d(n_7213), .o(n_7214) );
oa12f80 g565877 ( .a(n_1997), .b(x_in_49_15), .c(x_in_48_15), .o(n_29456) );
oa22f80 g565878 ( .a(n_520), .b(FE_OFN1106_rst), .c(n_29496), .d(n_3737), .o(n_6479) );
oa22f80 g565879 ( .a(n_1630), .b(FE_OFN60_n_27012), .c(FE_OFN412_n_28303), .d(n_7274), .o(n_7275) );
oa22f80 g565880 ( .a(n_1108), .b(FE_OFN74_n_27012), .c(n_29691), .d(n_7272), .o(n_7273) );
oa22f80 g565881 ( .a(n_1852), .b(FE_OFN350_n_4860), .c(FE_OFN404_n_28303), .d(n_7270), .o(n_7271) );
oa22f80 g565882 ( .a(n_627), .b(FE_OFN326_n_4860), .c(FE_OFN267_n_4280), .d(n_7268), .o(n_7269) );
in01f80 g565883 ( .a(n_5901), .o(n_5890) );
ao12f80 g565884 ( .a(n_7650), .b(n_5860), .c(x_in_21_6), .o(n_5901) );
oa22f80 g565885 ( .a(n_1460), .b(n_27449), .c(n_22019), .d(n_6711), .o(n_7267) );
in01f80 g565886 ( .a(n_5958), .o(n_5957) );
oa12f80 g565887 ( .a(n_7655), .b(n_5515), .c(x_in_3_8), .o(n_5958) );
oa22f80 g565888 ( .a(n_538), .b(FE_OFN90_n_27449), .c(FE_OFN308_n_3069), .d(n_8443), .o(n_7266) );
oa12f80 g565889 ( .a(n_1992), .b(x_in_41_15), .c(x_in_40_15), .o(n_29537) );
oa22f80 g565890 ( .a(n_1459), .b(n_27449), .c(FE_OFN400_n_28303), .d(n_8851), .o(n_7265) );
in01f80 g565891 ( .a(n_5913), .o(n_3357) );
no02f80 g565892 ( .a(n_4604), .b(n_2065), .o(n_5913) );
in01f80 g565893 ( .a(n_5026), .o(n_5024) );
oa12f80 g565894 ( .a(n_1979), .b(x_in_11_15), .c(x_in_11_14), .o(n_5026) );
oa22f80 g565895 ( .a(n_237), .b(FE_OFN89_n_27449), .c(n_29683), .d(n_7263), .o(n_7264) );
oa22f80 g565896 ( .a(n_1421), .b(FE_OFN104_n_27449), .c(n_29496), .d(n_7231), .o(n_7232) );
oa12f80 g565897 ( .a(n_2003), .b(x_in_9_4), .c(x_in_9_0), .o(n_3566) );
ao22s80 g565898 ( .a(n_2395), .b(n_2434), .c(x_in_1_1), .d(x_in_0_1), .o(n_3533) );
ao22s80 g565899 ( .a(n_2326), .b(n_1720), .c(x_in_45_15), .d(x_in_45_14), .o(n_3860) );
oa22f80 g565900 ( .a(x_in_29_15), .b(x_in_29_14), .c(n_2327), .d(n_3736), .o(n_3774) );
oa22f80 g565901 ( .a(x_in_13_15), .b(x_in_13_14), .c(n_3077), .d(n_2354), .o(n_3828) );
in01f80 g565902 ( .a(FE_OFN458_n_5621), .o(n_4908) );
oa22f80 g565903 ( .a(x_in_3_15), .b(x_in_3_14), .c(n_123), .d(n_2317), .o(n_5621) );
in01f80 g565904 ( .a(n_3013), .o(n_3014) );
oa22f80 g565905 ( .a(x_in_51_15), .b(x_in_51_14), .c(n_558), .d(n_2269), .o(n_3013) );
in01f80 g565906 ( .a(n_3989), .o(n_4767) );
oa22f80 g565907 ( .a(x_in_3_2), .b(x_in_3_0), .c(n_2272), .d(n_2139), .o(n_3989) );
in01f80 g565908 ( .a(n_5251), .o(n_5253) );
oa22f80 g565909 ( .a(x_in_19_2), .b(x_in_19_0), .c(n_2440), .d(n_2039), .o(n_5251) );
ao22s80 g565910 ( .a(n_2540), .b(n_2539), .c(x_in_5_3), .d(x_in_5_1), .o(n_3355) );
in01f80 g565911 ( .a(FE_OFN726_n_5240), .o(n_5241) );
ao22s80 g565912 ( .a(n_2538), .b(n_2052), .c(x_in_33_15), .d(x_in_33_14), .o(n_5240) );
in01f80 g565913 ( .a(n_5338), .o(n_3012) );
oa22f80 g565914 ( .a(x_in_13_15), .b(x_in_13_12), .c(n_5926), .d(n_2354), .o(n_5338) );
in01f80 g565915 ( .a(n_4694), .o(n_6779) );
oa22f80 g565916 ( .a(x_in_39_4), .b(x_in_39_3), .c(n_3107), .d(n_2537), .o(n_4694) );
in01f80 g565917 ( .a(n_5278), .o(n_5279) );
oa22f80 g565918 ( .a(x_in_27_15), .b(x_in_27_14), .c(n_2536), .d(n_14997), .o(n_5278) );
ao22s80 g565919 ( .a(n_5296), .b(n_2567), .c(x_in_5_5), .d(x_in_4_1), .o(n_3975) );
ao22s80 g565920 ( .a(n_2428), .b(n_2134), .c(x_in_45_10), .d(x_in_45_9), .o(n_6086) );
oa22f80 g565921 ( .a(n_1021), .b(x_in_25_2), .c(n_2535), .d(x_in_25_0), .o(n_5277) );
in01f80 g565922 ( .a(FE_OFN612_n_5698), .o(n_5243) );
oa22f80 g565923 ( .a(x_in_19_15), .b(x_in_19_14), .c(n_149), .d(n_4057), .o(n_5698) );
in01f80 g565924 ( .a(n_5273), .o(n_5274) );
oa22f80 g565925 ( .a(x_in_43_15), .b(x_in_43_14), .c(n_2394), .d(n_7311), .o(n_5273) );
in01f80 g565926 ( .a(FE_OFN765_n_5707), .o(n_5031) );
oa22f80 g565927 ( .a(x_in_35_15), .b(x_in_35_14), .c(n_1388), .d(n_2752), .o(n_5707) );
in01f80 g565928 ( .a(n_3008), .o(n_3009) );
oa22f80 g565929 ( .a(x_in_21_15), .b(x_in_21_14), .c(n_3043), .d(n_2309), .o(n_3008) );
oa22f80 g565930 ( .a(x_in_5_15), .b(x_in_4_14), .c(n_23944), .d(n_2403), .o(n_24652) );
oa22f80 g565931 ( .a(x_in_41_15), .b(x_in_41_14), .c(n_1175), .d(n_8032), .o(n_4979) );
ao22s80 g565932 ( .a(n_4592), .b(n_2409), .c(x_in_29_2), .d(x_in_29_1), .o(n_4015) );
in01f80 g565933 ( .a(n_2785), .o(n_2786) );
ao22s80 g565934 ( .a(n_4946), .b(n_2593), .c(x_in_15_2), .d(x_in_15_1), .o(n_2785) );
in01f80 g565935 ( .a(n_3006), .o(n_3007) );
ao22s80 g565936 ( .a(n_5365), .b(n_2616), .c(x_in_47_2), .d(x_in_47_1), .o(n_3006) );
in01f80 g565937 ( .a(n_5297), .o(n_5295) );
oa22f80 g565938 ( .a(x_in_5_4), .b(x_in_5_2), .c(n_2517), .d(n_2413), .o(n_5297) );
in01f80 g565939 ( .a(n_2697), .o(n_2698) );
ao22s80 g565940 ( .a(n_5336), .b(n_2618), .c(x_in_55_2), .d(x_in_55_1), .o(n_2697) );
oa22f80 g565941 ( .a(x_in_31_2), .b(x_in_31_1), .c(n_5373), .d(n_2660), .o(n_9044) );
in01f80 g565942 ( .a(n_3004), .o(n_3005) );
ao22s80 g565943 ( .a(n_5351), .b(n_2603), .c(x_in_63_2), .d(x_in_63_1), .o(n_3004) );
in01f80 g565944 ( .a(n_3002), .o(n_3003) );
ao22s80 g565945 ( .a(n_5430), .b(n_2646), .c(x_in_23_2), .d(x_in_23_1), .o(n_3002) );
in01f80 g565946 ( .a(n_7490), .o(n_3001) );
oa22f80 g565947 ( .a(x_in_39_13), .b(x_in_39_11), .c(n_7317), .d(n_7213), .o(n_7490) );
in01f80 g565948 ( .a(n_4991), .o(n_2819) );
ao22s80 g565949 ( .a(n_4409), .b(n_2422), .c(x_in_59_15), .d(x_in_59_14), .o(n_4991) );
oa22f80 g565950 ( .a(n_2534), .b(x_in_41_1), .c(n_533), .d(x_in_41_0), .o(n_6081) );
oa22f80 g565951 ( .a(n_2235), .b(x_in_1_1), .c(n_2395), .d(x_in_1_0), .o(n_4808) );
in01f80 g565952 ( .a(n_9032), .o(n_9038) );
ao22s80 g565953 ( .a(n_2433), .b(n_2505), .c(x_in_13_5), .d(x_in_13_4), .o(n_9032) );
in01f80 g565954 ( .a(n_10390), .o(n_3000) );
oa22f80 g565955 ( .a(x_in_45_9), .b(x_in_45_8), .c(n_2527), .d(n_2428), .o(n_10390) );
in01f80 g565956 ( .a(n_5374), .o(n_5375) );
oa22f80 g565957 ( .a(x_in_7_15), .b(x_in_7_14), .c(n_15590), .d(n_2624), .o(n_5374) );
in01f80 g565958 ( .a(n_10405), .o(n_2829) );
ao22s80 g565959 ( .a(n_5986), .b(n_2439), .c(x_in_45_3), .d(x_in_45_2), .o(n_10405) );
in01f80 g565960 ( .a(n_10406), .o(n_2831) );
oa22f80 g565961 ( .a(x_in_45_4), .b(x_in_45_3), .c(n_2442), .d(n_2439), .o(n_10406) );
oa22f80 g565962 ( .a(x_in_11_13), .b(x_in_11_10), .c(n_3229), .d(n_2681), .o(n_3934) );
in01f80 g565963 ( .a(FE_OFN544_n_9030), .o(n_9034) );
oa22f80 g565964 ( .a(x_in_13_4), .b(x_in_13_3), .c(n_2433), .d(n_2516), .o(n_9030) );
oa22f80 g565965 ( .a(x_in_9_12), .b(x_in_9_11), .c(n_8957), .d(n_2488), .o(n_3938) );
in01f80 g565966 ( .a(FE_OFN546_n_9036), .o(n_9042) );
oa22f80 g565967 ( .a(x_in_13_6), .b(x_in_13_5), .c(n_2506), .d(n_2505), .o(n_9036) );
in01f80 g565968 ( .a(n_9480), .o(n_11700) );
oa22f80 g565969 ( .a(x_in_13_8), .b(x_in_13_7), .c(n_2657), .d(n_2522), .o(n_9480) );
in01f80 g565970 ( .a(FE_OFN548_n_10452), .o(n_9638) );
oa22f80 g565971 ( .a(x_in_13_7), .b(x_in_13_6), .c(n_2506), .d(n_2657), .o(n_10452) );
in01f80 g565972 ( .a(n_10413), .o(n_10392) );
oa22f80 g565973 ( .a(x_in_45_7), .b(x_in_45_6), .c(n_2513), .d(n_2528), .o(n_10413) );
in01f80 g565974 ( .a(FE_OFN801_n_6782), .o(n_4717) );
oa22f80 g565975 ( .a(x_in_39_6), .b(x_in_39_5), .c(n_4338), .d(n_6500), .o(n_6782) );
in01f80 g565976 ( .a(FE_OFN552_n_9482), .o(n_4603) );
oa22f80 g565977 ( .a(x_in_13_9), .b(x_in_13_8), .c(n_2522), .d(n_2521), .o(n_9482) );
in01f80 g565978 ( .a(n_10351), .o(n_9458) );
oa22f80 g565979 ( .a(x_in_45_8), .b(x_in_45_7), .c(n_2528), .d(n_2527), .o(n_10351) );
in01f80 g565980 ( .a(n_5307), .o(n_4669) );
oa22f80 g565981 ( .a(x_in_57_4), .b(x_in_57_2), .c(n_2601), .d(n_2222), .o(n_5307) );
in01f80 g565982 ( .a(FE_OFN1256_n_10520), .o(n_3010) );
oa22f80 g565983 ( .a(x_in_55_4), .b(x_in_55_3), .c(n_3742), .d(n_3079), .o(n_10520) );
in01f80 g565984 ( .a(n_10550), .o(n_9514) );
oa22f80 g565985 ( .a(x_in_15_4), .b(x_in_15_3), .c(n_3482), .d(n_2780), .o(n_10550) );
in01f80 g565986 ( .a(FE_OFN1238_n_10491), .o(n_2749) );
oa22f80 g565987 ( .a(x_in_47_4), .b(x_in_47_3), .c(n_3445), .d(n_2747), .o(n_10491) );
in01f80 g565988 ( .a(n_9024), .o(n_10418) );
oa22f80 g565989 ( .a(x_in_23_4), .b(x_in_23_3), .c(n_3744), .d(n_3075), .o(n_9024) );
in01f80 g565990 ( .a(n_5358), .o(n_5357) );
oa22f80 g565991 ( .a(x_in_17_15), .b(x_in_17_14), .c(n_4794), .d(n_2549), .o(n_5358) );
in01f80 g565992 ( .a(FE_OFN1208_n_10456), .o(n_3023) );
oa22f80 g565993 ( .a(x_in_31_4), .b(x_in_31_3), .c(n_3739), .d(n_2721), .o(n_10456) );
in01f80 g565994 ( .a(n_10435), .o(n_2996) );
oa22f80 g565995 ( .a(x_in_63_4), .b(x_in_63_3), .c(n_3737), .d(n_2828), .o(n_10435) );
in01f80 g565996 ( .a(n_5176), .o(n_7449) );
oa22f80 g565997 ( .a(x_in_39_9), .b(x_in_39_8), .c(n_8133), .d(n_4514), .o(n_5176) );
in01f80 g565998 ( .a(n_5170), .o(n_7553) );
oa22f80 g565999 ( .a(x_in_39_5), .b(x_in_39_4), .c(n_3107), .d(n_4338), .o(n_5170) );
ao22s80 g566000 ( .a(n_2864), .b(n_2597), .c(x_in_29_9), .d(x_in_29_8), .o(n_6715) );
in01f80 g566001 ( .a(n_5159), .o(n_7503) );
oa22f80 g566002 ( .a(x_in_39_7), .b(x_in_39_6), .c(n_6500), .d(n_7325), .o(n_5159) );
in01f80 g566003 ( .a(n_3518), .o(n_3270) );
ao22s80 g566004 ( .a(n_8957), .b(n_2643), .c(x_in_9_15), .d(x_in_9_12), .o(n_3518) );
in01f80 g566005 ( .a(n_7002), .o(n_8449) );
oa22f80 g566006 ( .a(x_in_11_14), .b(x_in_11_11), .c(n_7818), .d(n_2124), .o(n_7002) );
in01f80 g566007 ( .a(FE_OFN554_n_9468), .o(n_12366) );
oa22f80 g566008 ( .a(x_in_13_10), .b(x_in_13_9), .c(n_2521), .d(n_2673), .o(n_9468) );
ao22s80 g566009 ( .a(n_3591), .b(n_3724), .c(x_in_29_4), .d(x_in_29_3), .o(n_6708) );
in01f80 g566010 ( .a(FE_OFN843_n_10412), .o(n_3192) );
ao22s80 g566011 ( .a(n_2513), .b(n_2438), .c(x_in_45_6), .d(x_in_45_5), .o(n_10412) );
in01f80 g566012 ( .a(n_4677), .o(n_6744) );
oa22f80 g566013 ( .a(x_in_29_7), .b(x_in_29_6), .c(n_3390), .d(n_3035), .o(n_4677) );
in01f80 g566014 ( .a(n_6749), .o(n_2995) );
oa22f80 g566015 ( .a(x_in_29_8), .b(x_in_29_7), .c(n_3035), .d(n_2864), .o(n_6749) );
in01f80 g566016 ( .a(n_5166), .o(n_7466) );
oa22f80 g566017 ( .a(x_in_39_8), .b(x_in_39_7), .c(n_7325), .d(n_8133), .o(n_5166) );
in01f80 g566018 ( .a(n_6713), .o(n_2994) );
oa22f80 g566019 ( .a(x_in_29_6), .b(x_in_29_5), .c(n_3470), .d(n_3390), .o(n_6713) );
in01f80 g566020 ( .a(FE_OFN576_n_10136), .o(n_10138) );
oa22f80 g566021 ( .a(x_in_15_13), .b(x_in_15_11), .c(n_7334), .d(n_2575), .o(n_10136) );
ao22s80 g566022 ( .a(n_4847), .b(n_2655), .c(x_in_61_15), .d(x_in_61_14), .o(n_5391) );
in01f80 g566023 ( .a(n_10133), .o(n_10135) );
oa22f80 g566024 ( .a(x_in_47_13), .b(x_in_47_11), .c(n_7245), .d(n_2448), .o(n_10133) );
in01f80 g566025 ( .a(n_11028), .o(n_11030) );
oa22f80 g566026 ( .a(x_in_63_13), .b(x_in_63_11), .c(n_7308), .d(n_2523), .o(n_11028) );
in01f80 g566027 ( .a(n_9072), .o(n_2993) );
ao22s80 g566028 ( .a(n_7336), .b(n_2624), .c(x_in_7_15), .d(x_in_7_11), .o(n_9072) );
in01f80 g566029 ( .a(FE_OFN803_n_6771), .o(n_4674) );
oa22f80 g566030 ( .a(x_in_39_10), .b(x_in_39_9), .c(n_4514), .d(n_8851), .o(n_6771) );
in01f80 g566031 ( .a(n_5068), .o(n_6727) );
oa22f80 g566032 ( .a(x_in_29_10), .b(x_in_29_9), .c(n_2597), .d(n_8537), .o(n_5068) );
ao22s80 g566033 ( .a(n_3724), .b(n_3470), .c(x_in_29_5), .d(x_in_29_4), .o(n_6709) );
in01f80 g566034 ( .a(n_10400), .o(n_2992) );
oa22f80 g566035 ( .a(x_in_45_5), .b(x_in_45_4), .c(n_2438), .d(n_2442), .o(n_10400) );
in01f80 g566036 ( .a(n_8861), .o(n_3278) );
oa22f80 g566037 ( .a(x_in_45_2), .b(x_in_45_1), .c(n_2385), .d(n_5986), .o(n_8861) );
in01f80 g566038 ( .a(n_8532), .o(n_4613) );
oa22f80 g566039 ( .a(x_in_57_14), .b(x_in_57_11), .c(n_5313), .d(n_442), .o(n_8532) );
in01f80 g566040 ( .a(n_10139), .o(n_10141) );
oa22f80 g566041 ( .a(x_in_55_13), .b(x_in_55_11), .c(n_7332), .d(n_7231), .o(n_10139) );
in01f80 g566042 ( .a(n_10145), .o(n_10147) );
oa22f80 g566043 ( .a(x_in_23_13), .b(x_in_23_11), .c(n_7296), .d(n_6488), .o(n_10145) );
in01f80 g566044 ( .a(n_11031), .o(n_11033) );
oa22f80 g566045 ( .a(x_in_31_13), .b(x_in_31_11), .c(n_7298), .d(n_7291), .o(n_11031) );
in01f80 g566046 ( .a(n_10544), .o(n_9461) );
oa22f80 g566047 ( .a(x_in_55_5), .b(x_in_55_4), .c(n_3742), .d(n_4329), .o(n_10544) );
in01f80 g566048 ( .a(n_10396), .o(n_9454) );
oa22f80 g566049 ( .a(x_in_15_5), .b(x_in_15_4), .c(n_3482), .d(n_4746), .o(n_10396) );
in01f80 g566050 ( .a(n_9054), .o(n_10430) );
oa22f80 g566051 ( .a(x_in_23_5), .b(x_in_23_4), .c(n_3744), .d(n_4744), .o(n_9054) );
in01f80 g566052 ( .a(n_5392), .o(n_2990) );
ao22s80 g566053 ( .a(n_3568), .b(n_5291), .c(x_in_5_8), .d(x_in_5_6), .o(n_5392) );
ao22s80 g566054 ( .a(n_2517), .b(n_3568), .c(x_in_5_6), .d(x_in_5_4), .o(n_5036) );
in01f80 g566055 ( .a(n_10437), .o(n_2989) );
ao22s80 g566056 ( .a(n_3737), .b(n_4745), .c(x_in_63_5), .d(x_in_63_4), .o(n_10437) );
oa22f80 g566057 ( .a(x_in_17_15), .b(x_in_17_12), .c(n_5415), .d(n_2549), .o(n_6230) );
in01f80 g566058 ( .a(FE_OFN1089_n_8985), .o(n_3016) );
ao22s80 g566059 ( .a(n_4529), .b(n_2655), .c(x_in_61_15), .d(x_in_61_11), .o(n_8985) );
in01f80 g566060 ( .a(n_3376), .o(n_5674) );
oa22f80 g566061 ( .a(x_in_61_4), .b(x_in_61_0), .c(n_8929), .d(n_2605), .o(n_3376) );
oa22f80 g566062 ( .a(x_in_59_13), .b(x_in_59_10), .c(n_2668), .d(n_2635), .o(n_3571) );
in01f80 g566063 ( .a(n_5294), .o(n_2988) );
oa22f80 g566064 ( .a(x_in_5_5), .b(x_in_5_3), .c(n_2540), .d(n_5296), .o(n_5294) );
in01f80 g566065 ( .a(FE_OFN1210_n_10458), .o(n_2985) );
ao22s80 g566066 ( .a(n_4738), .b(n_3739), .c(x_in_31_5), .d(x_in_31_4), .o(n_10458) );
in01f80 g566067 ( .a(FE_OFN861_n_10492), .o(n_2984) );
ao22s80 g566068 ( .a(n_4737), .b(n_3445), .c(x_in_47_5), .d(x_in_47_4), .o(n_10492) );
in01f80 g566069 ( .a(n_5389), .o(n_2983) );
oa22f80 g566070 ( .a(x_in_5_9), .b(x_in_5_7), .c(n_2645), .d(n_6000), .o(n_5389) );
in01f80 g566071 ( .a(n_9678), .o(n_10548) );
oa22f80 g566072 ( .a(x_in_55_9), .b(x_in_55_8), .c(n_7315), .d(n_10915), .o(n_9678) );
in01f80 g566073 ( .a(FE_OFN1240_n_10499), .o(n_9493) );
oa22f80 g566074 ( .a(x_in_47_7), .b(x_in_47_6), .c(n_7901), .d(n_6683), .o(n_10499) );
in01f80 g566075 ( .a(n_10355), .o(n_9473) );
oa22f80 g566076 ( .a(x_in_63_9), .b(x_in_63_8), .c(n_7272), .d(n_10916), .o(n_10355) );
in01f80 g566077 ( .a(n_10547), .o(n_9517) );
oa22f80 g566078 ( .a(x_in_55_6), .b(x_in_55_5), .c(n_4329), .d(n_6685), .o(n_10547) );
in01f80 g566079 ( .a(n_10525), .o(n_9502) );
oa22f80 g566080 ( .a(x_in_55_7), .b(x_in_55_6), .c(n_7905), .d(n_6685), .o(n_10525) );
in01f80 g566081 ( .a(FE_OFN658_n_10424), .o(n_2982) );
ao22s80 g566082 ( .a(n_7270), .b(n_10918), .c(x_in_23_9), .d(x_in_23_8), .o(n_10424) );
in01f80 g566083 ( .a(n_5288), .o(n_2981) );
oa22f80 g566084 ( .a(x_in_5_12), .b(x_in_5_10), .c(n_5388), .d(n_5888), .o(n_5288) );
in01f80 g566085 ( .a(FE_OFN869_n_10506), .o(n_9499) );
oa22f80 g566086 ( .a(x_in_47_9), .b(x_in_47_8), .c(n_7241), .d(n_10913), .o(n_10506) );
in01f80 g566087 ( .a(FE_OFN865_n_10501), .o(n_9496) );
oa22f80 g566088 ( .a(x_in_47_8), .b(x_in_47_7), .c(n_7901), .d(n_7241), .o(n_10501) );
in01f80 g566089 ( .a(n_10398), .o(n_9506) );
oa22f80 g566090 ( .a(x_in_23_7), .b(x_in_23_6), .c(n_7906), .d(n_6689), .o(n_10398) );
in01f80 g566091 ( .a(n_9673), .o(n_10537) );
oa22f80 g566092 ( .a(x_in_15_6), .b(x_in_15_5), .c(n_4746), .d(n_6687), .o(n_9673) );
in01f80 g566093 ( .a(n_10442), .o(n_9470) );
oa22f80 g566094 ( .a(x_in_63_8), .b(x_in_63_7), .c(n_7903), .d(n_7272), .o(n_10442) );
in01f80 g566095 ( .a(n_10472), .o(n_9477) );
oa22f80 g566096 ( .a(x_in_31_9), .b(x_in_31_8), .c(n_8200), .d(n_10914), .o(n_10472) );
in01f80 g566097 ( .a(n_5290), .o(n_2980) );
oa22f80 g566098 ( .a(x_in_5_10), .b(x_in_5_8), .c(n_5291), .d(n_5388), .o(n_5290) );
in01f80 g566099 ( .a(n_10367), .o(n_2979) );
oa22f80 g566100 ( .a(x_in_63_6), .b(x_in_63_5), .c(n_4745), .d(n_6711), .o(n_10367) );
in01f80 g566101 ( .a(FE_OFN656_n_10503), .o(n_3299) );
oa22f80 g566102 ( .a(x_in_23_6), .b(x_in_23_5), .c(n_4744), .d(n_6689), .o(n_10503) );
in01f80 g566103 ( .a(FE_OFN1214_n_10469), .o(n_2978) );
oa22f80 g566104 ( .a(x_in_31_8), .b(x_in_31_7), .c(n_7902), .d(n_8200), .o(n_10469) );
in01f80 g566105 ( .a(n_8991), .o(n_10513) );
oa22f80 g566106 ( .a(x_in_15_8), .b(x_in_15_7), .c(n_7904), .d(n_6492), .o(n_8991) );
in01f80 g566107 ( .a(n_10526), .o(n_9451) );
oa22f80 g566108 ( .a(x_in_55_8), .b(x_in_55_7), .c(n_7905), .d(n_7315), .o(n_10526) );
in01f80 g566109 ( .a(n_10370), .o(n_9523) );
oa22f80 g566110 ( .a(x_in_63_7), .b(x_in_63_6), .c(n_7903), .d(n_6711), .o(n_10370) );
in01f80 g566111 ( .a(n_9063), .o(n_10555) );
oa22f80 g566112 ( .a(x_in_15_7), .b(x_in_15_6), .c(n_7904), .d(n_6687), .o(n_9063) );
in01f80 g566113 ( .a(n_10535), .o(n_9509) );
oa22f80 g566114 ( .a(x_in_23_8), .b(x_in_23_7), .c(n_7906), .d(n_7270), .o(n_10535) );
in01f80 g566115 ( .a(FE_OFN1212_n_10465), .o(n_2977) );
ao22s80 g566116 ( .a(n_7902), .b(n_6483), .c(x_in_31_7), .d(x_in_31_6), .o(n_10465) );
in01f80 g566117 ( .a(n_9079), .o(n_10516) );
oa22f80 g566118 ( .a(x_in_15_9), .b(x_in_15_8), .c(n_6492), .d(n_10917), .o(n_9079) );
oa22f80 g566119 ( .a(x_in_37_13), .b(x_in_37_10), .c(n_5745), .d(n_4343), .o(n_3577) );
ao22s80 g566120 ( .a(n_2526), .b(n_4668), .c(x_in_57_5), .d(x_in_57_3), .o(n_5306) );
ao22s80 g566121 ( .a(n_4668), .b(n_2601), .c(x_in_57_5), .d(x_in_57_4), .o(n_4132) );
in01f80 g566122 ( .a(n_5361), .o(n_2976) );
oa22f80 g566123 ( .a(x_in_57_6), .b(x_in_57_4), .c(n_2601), .d(n_2512), .o(n_5361) );
in01f80 g566124 ( .a(FE_OFN704_n_10462), .o(n_2975) );
oa22f80 g566125 ( .a(x_in_31_6), .b(x_in_31_5), .c(n_4738), .d(n_6483), .o(n_10462) );
oa22f80 g566126 ( .a(x_in_19_13), .b(x_in_19_10), .c(n_3020), .d(n_5556), .o(n_3620) );
in01f80 g566127 ( .a(FE_OFN863_n_10495), .o(n_2973) );
oa22f80 g566128 ( .a(x_in_47_6), .b(x_in_47_5), .c(n_4737), .d(n_6683), .o(n_10495) );
in01f80 g566129 ( .a(n_3866), .o(n_2972) );
ao22s80 g566130 ( .a(n_4180), .b(n_2419), .c(x_in_37_11), .d(x_in_37_14), .o(n_3866) );
in01f80 g566131 ( .a(n_8848), .o(n_7879) );
oa22f80 g566132 ( .a(x_in_59_14), .b(x_in_59_11), .c(n_8482), .d(n_2422), .o(n_8848) );
in01f80 g566133 ( .a(n_2970), .o(n_2971) );
oa22f80 g566134 ( .a(x_in_43_13), .b(x_in_43_10), .c(n_6496), .d(n_7274), .o(n_2970) );
in01f80 g566135 ( .a(n_2968), .o(n_2969) );
oa22f80 g566136 ( .a(x_in_27_13), .b(x_in_27_10), .c(n_7417), .d(n_7229), .o(n_2968) );
in01f80 g566137 ( .a(n_5292), .o(n_2966) );
oa22f80 g566138 ( .a(x_in_5_7), .b(x_in_5_5), .c(n_5296), .d(n_2645), .o(n_5292) );
in01f80 g566139 ( .a(n_6963), .o(n_8506) );
oa22f80 g566140 ( .a(x_in_3_14), .b(x_in_3_11), .c(n_6380), .d(n_2317), .o(n_6963) );
ao22s80 g566141 ( .a(n_4668), .b(n_4055), .c(x_in_57_7), .d(x_in_57_5), .o(n_5305) );
in01f80 g566142 ( .a(n_5304), .o(n_2965) );
oa22f80 g566143 ( .a(x_in_57_9), .b(x_in_57_7), .c(n_4055), .d(n_3245), .o(n_5304) );
in01f80 g566144 ( .a(n_5298), .o(n_2964) );
oa22f80 g566145 ( .a(x_in_57_8), .b(x_in_57_6), .c(n_2512), .d(n_2627), .o(n_5298) );
in01f80 g566146 ( .a(n_6970), .o(n_8504) );
oa22f80 g566147 ( .a(x_in_27_14), .b(x_in_27_11), .c(n_8513), .d(n_14997), .o(n_6970) );
in01f80 g566148 ( .a(n_2962), .o(n_2963) );
oa22f80 g566149 ( .a(x_in_61_13), .b(x_in_61_10), .c(n_3833), .d(n_2518), .o(n_2962) );
in01f80 g566150 ( .a(n_9622), .o(n_2961) );
oa22f80 g566151 ( .a(x_in_7_14), .b(x_in_7_11), .c(n_7336), .d(n_15590), .o(n_9622) );
in01f80 g566152 ( .a(n_2959), .o(n_2960) );
oa22f80 g566153 ( .a(x_in_7_13), .b(x_in_7_10), .c(n_8165), .d(n_7285), .o(n_2959) );
in01f80 g566154 ( .a(n_5314), .o(n_2958) );
oa22f80 g566155 ( .a(x_in_57_10), .b(x_in_57_8), .c(n_2627), .d(n_3409), .o(n_5314) );
in01f80 g566156 ( .a(n_5276), .o(n_2957) );
oa22f80 g566157 ( .a(x_in_57_12), .b(x_in_57_10), .c(n_3409), .d(n_5302), .o(n_5276) );
in01f80 g566158 ( .a(n_3899), .o(n_8530) );
oa22f80 g566159 ( .a(x_in_5_14), .b(x_in_5_11), .c(n_5754), .d(n_3169), .o(n_3899) );
in01f80 g566160 ( .a(n_5485), .o(n_2956) );
ao22s80 g566161 ( .a(n_2548), .b(n_3193), .c(x_in_53_15), .d(x_in_53_12), .o(n_5485) );
in01f80 g566162 ( .a(n_5289), .o(n_2955) );
oa22f80 g566163 ( .a(x_in_5_11), .b(x_in_5_9), .c(n_6000), .d(n_5754), .o(n_5289) );
in01f80 g566164 ( .a(n_6464), .o(n_8445) );
oa22f80 g566165 ( .a(x_in_43_14), .b(x_in_43_11), .c(n_8443), .d(n_7311), .o(n_6464) );
in01f80 g566166 ( .a(n_4640), .o(n_4101) );
no02f80 g566167 ( .a(n_2138), .b(n_2023), .o(n_4640) );
oa22f80 g566168 ( .a(x_in_53_6), .b(x_in_53_4), .c(n_3038), .d(n_2651), .o(n_3400) );
oa22f80 g566169 ( .a(x_in_53_8), .b(x_in_53_6), .c(n_2654), .d(n_2651), .o(n_3531) );
oa22f80 g566170 ( .a(x_in_53_9), .b(x_in_53_7), .c(n_2550), .d(n_2525), .o(n_3546) );
in01f80 g566171 ( .a(n_10475), .o(n_9484) );
oa22f80 g566172 ( .a(x_in_31_10), .b(x_in_31_9), .c(n_10914), .d(n_11698), .o(n_10475) );
in01f80 g566173 ( .a(n_10507), .o(n_9487) );
oa22f80 g566174 ( .a(x_in_47_10), .b(x_in_47_9), .c(n_10913), .d(n_11034), .o(n_10507) );
in01f80 g566175 ( .a(n_10557), .o(n_10510) );
oa22f80 g566176 ( .a(x_in_15_10), .b(x_in_15_9), .c(n_10917), .d(n_11037), .o(n_10557) );
in01f80 g566177 ( .a(n_10444), .o(n_9490) );
oa22f80 g566178 ( .a(x_in_63_10), .b(x_in_63_9), .c(n_10916), .d(n_11696), .o(n_10444) );
in01f80 g566179 ( .a(n_10539), .o(n_10517) );
oa22f80 g566180 ( .a(x_in_55_10), .b(x_in_55_9), .c(n_10915), .d(n_11040), .o(n_10539) );
in01f80 g566181 ( .a(n_10541), .o(n_10531) );
oa22f80 g566182 ( .a(x_in_23_10), .b(x_in_23_9), .c(n_10918), .d(n_11041), .o(n_10541) );
in01f80 g566183 ( .a(n_5303), .o(n_2954) );
oa22f80 g566184 ( .a(x_in_57_11), .b(x_in_57_9), .c(n_3245), .d(n_5313), .o(n_5303) );
oa22f80 g566185 ( .a(x_in_53_11), .b(x_in_53_9), .c(n_2870), .d(n_2550), .o(n_4139) );
ao22s80 g566186 ( .a(n_5827), .b(n_4825), .c(x_in_53_3), .d(x_in_53_1), .o(n_4327) );
oa22f80 g566187 ( .a(x_in_53_7), .b(x_in_53_5), .c(n_2626), .d(n_2525), .o(n_3536) );
in01f80 g566188 ( .a(FE_OFN1272_n_9600), .o(n_2953) );
ao22s80 g566189 ( .a(n_4529), .b(n_4847), .c(x_in_61_14), .d(x_in_61_11), .o(n_9600) );
oa22f80 g566190 ( .a(x_in_51_13), .b(x_in_51_10), .c(n_5283), .d(n_5689), .o(n_3486) );
in01f80 g566191 ( .a(n_6947), .o(n_8486) );
oa22f80 g566192 ( .a(x_in_19_14), .b(x_in_19_11), .c(n_7765), .d(n_4057), .o(n_6947) );
oa22f80 g566193 ( .a(x_in_53_10), .b(x_in_53_8), .c(n_2654), .d(n_2653), .o(n_3964) );
oa22f80 g566194 ( .a(x_in_25_6), .b(x_in_25_4), .c(n_2554), .d(n_3771), .o(n_3947) );
oa22f80 g566195 ( .a(x_in_53_12), .b(x_in_53_10), .c(n_2653), .d(n_2548), .o(n_3955) );
oa22f80 g566196 ( .a(x_in_3_13), .b(x_in_3_10), .c(n_5666), .d(n_6746), .o(n_3922) );
in01f80 g566197 ( .a(n_5280), .o(n_2952) );
ao22s80 g566198 ( .a(n_5247), .b(n_6380), .c(x_in_3_12), .d(x_in_3_11), .o(n_5280) );
in01f80 g566199 ( .a(n_5669), .o(n_2951) );
oa22f80 g566200 ( .a(x_in_17_4), .b(x_in_17_2), .c(n_4021), .d(n_4687), .o(n_5669) );
oa22f80 g566201 ( .a(x_in_25_7), .b(x_in_25_5), .c(n_3132), .d(n_4593), .o(n_3465) );
oa22f80 g566202 ( .a(x_in_35_12), .b(x_in_35_11), .c(n_8524), .d(n_5032), .o(n_3961) );
in01f80 g566203 ( .a(n_4812), .o(n_3317) );
ao22s80 g566204 ( .a(n_9651), .b(n_9646), .c(x_in_17_7), .d(x_in_17_5), .o(n_4812) );
in01f80 g566205 ( .a(n_4819), .o(n_2745) );
oa22f80 g566206 ( .a(x_in_25_15), .b(x_in_25_12), .c(n_5317), .d(n_2546), .o(n_4819) );
ao22s80 g566207 ( .a(n_2870), .b(n_5988), .c(x_in_53_13), .d(x_in_53_11), .o(n_3624) );
oa22f80 g566208 ( .a(x_in_53_5), .b(x_in_53_3), .c(n_2626), .d(n_5827), .o(n_3969) );
in01f80 g566209 ( .a(n_4871), .o(n_3180) );
oa22f80 g566210 ( .a(x_in_17_12), .b(x_in_17_10), .c(n_5415), .d(n_5359), .o(n_4871) );
in01f80 g566211 ( .a(n_4811), .o(n_2947) );
oa22f80 g566212 ( .a(x_in_17_9), .b(x_in_17_7), .c(n_9654), .d(n_9651), .o(n_4811) );
oa22f80 g566213 ( .a(x_in_25_8), .b(x_in_25_6), .c(n_3129), .d(n_3771), .o(n_3944) );
in01f80 g566214 ( .a(n_5356), .o(n_2946) );
ao22s80 g566215 ( .a(n_5415), .b(n_5418), .c(x_in_17_12), .d(x_in_17_11), .o(n_5356) );
oa22f80 g566216 ( .a(x_in_25_9), .b(x_in_25_7), .c(n_3132), .d(n_2581), .o(n_3473) );
oa22f80 g566217 ( .a(x_in_25_10), .b(x_in_25_8), .c(n_3129), .d(n_2743), .o(n_3564) );
in01f80 g566218 ( .a(n_4816), .o(n_2774) );
oa22f80 g566219 ( .a(x_in_17_10), .b(x_in_17_8), .c(n_5360), .d(n_5359), .o(n_4816) );
in01f80 g566220 ( .a(n_4815), .o(n_3032) );
oa22f80 g566221 ( .a(x_in_17_11), .b(x_in_17_9), .c(n_5418), .d(n_9654), .o(n_4815) );
oa22f80 g566222 ( .a(x_in_25_11), .b(x_in_25_9), .c(n_2581), .d(n_3189), .o(n_3928) );
oa22f80 g566223 ( .a(x_in_25_12), .b(x_in_25_10), .c(n_2743), .d(n_5317), .o(n_3950) );
in01f80 g566224 ( .a(n_4868), .o(n_3240) );
oa22f80 g566225 ( .a(x_in_17_6), .b(x_in_17_4), .c(n_4021), .d(n_5362), .o(n_4868) );
in01f80 g566226 ( .a(n_4869), .o(n_3067) );
oa22f80 g566227 ( .a(x_in_17_8), .b(x_in_17_6), .c(n_5360), .d(n_5362), .o(n_4869) );
in01f80 g566228 ( .a(n_5384), .o(n_2945) );
oa22f80 g566229 ( .a(n_7213), .b(x_in_39_14), .c(n_2343), .d(x_in_39_13), .o(n_5384) );
in01f80 g566230 ( .a(n_5364), .o(n_2944) );
oa22f80 g566231 ( .a(n_2616), .b(x_in_47_5), .c(n_4737), .d(x_in_47_1), .o(n_5364) );
ao22s80 g566232 ( .a(n_2558), .b(x_in_47_11), .c(n_7245), .d(x_in_47_14), .o(n_6157) );
in01f80 g566233 ( .a(n_5372), .o(n_2692) );
oa22f80 g566234 ( .a(n_2660), .b(x_in_31_5), .c(n_4738), .d(x_in_31_1), .o(n_5372) );
ao22s80 g566235 ( .a(n_2606), .b(x_in_63_11), .c(n_7308), .d(x_in_63_14), .o(n_6116) );
ao22s80 g566236 ( .a(n_2574), .b(x_in_15_11), .c(n_7334), .d(x_in_15_14), .o(n_6424) );
ao22s80 g566237 ( .a(n_1624), .b(x_in_49_14), .c(n_9118), .d(x_in_49_15), .o(n_3462) );
in01f80 g566238 ( .a(n_4945), .o(n_2943) );
oa22f80 g566239 ( .a(n_2593), .b(x_in_15_5), .c(n_4746), .d(x_in_15_1), .o(n_4945) );
in01f80 g566240 ( .a(n_5380), .o(n_3228) );
oa22f80 g566241 ( .a(n_2646), .b(x_in_23_5), .c(n_4744), .d(x_in_23_1), .o(n_5380) );
in01f80 g566242 ( .a(n_5350), .o(n_2942) );
oa22f80 g566243 ( .a(n_2603), .b(x_in_63_5), .c(n_4745), .d(x_in_63_1), .o(n_5350) );
in01f80 g566244 ( .a(n_5335), .o(n_2941) );
oa22f80 g566245 ( .a(n_2618), .b(x_in_55_5), .c(n_4329), .d(x_in_55_1), .o(n_5335) );
ao22s80 g566246 ( .a(n_2549), .b(x_in_17_13), .c(n_10477), .d(x_in_17_15), .o(n_4176) );
in01f80 g566247 ( .a(n_5270), .o(n_2861) );
oa22f80 g566248 ( .a(n_2509), .b(x_in_59_3), .c(n_3260), .d(x_in_59_1), .o(n_5270) );
in01f80 g566249 ( .a(n_2802), .o(n_2803) );
oa22f80 g566250 ( .a(n_2408), .b(x_in_7_5), .c(n_5256), .d(x_in_7_1), .o(n_2802) );
oa22f80 g566251 ( .a(n_2349), .b(x_in_43_4), .c(n_5293), .d(x_in_43_2), .o(n_3959) );
oa22f80 g566252 ( .a(n_2478), .b(x_in_27_4), .c(n_5679), .d(x_in_27_2), .o(n_3930) );
in01f80 g566253 ( .a(n_5318), .o(n_2940) );
ao22s80 g566254 ( .a(n_2492), .b(x_in_25_11), .c(n_3189), .d(x_in_25_14), .o(n_5318) );
ao22s80 g566255 ( .a(n_16158), .b(x_in_23_11), .c(n_7296), .d(x_in_23_14), .o(n_6169) );
ao22s80 g566256 ( .a(n_16156), .b(x_in_55_11), .c(n_7332), .d(x_in_55_14), .o(n_6181) );
ao22s80 g566257 ( .a(n_16154), .b(x_in_31_11), .c(n_7298), .d(x_in_31_14), .o(n_6089) );
oa22f80 g566258 ( .a(n_2332), .b(x_in_11_4), .c(n_5387), .d(x_in_11_2), .o(n_3554) );
in01f80 g566259 ( .a(n_5284), .o(n_2937) );
oa22f80 g566260 ( .a(n_2664), .b(x_in_43_3), .c(n_2541), .d(x_in_43_1), .o(n_5284) );
in01f80 g566261 ( .a(n_5386), .o(n_2936) );
oa22f80 g566262 ( .a(n_2365), .b(x_in_11_3), .c(n_2431), .d(x_in_11_1), .o(n_5386) );
oa22f80 g566263 ( .a(n_3186), .b(x_in_49_13), .c(n_2691), .d(x_in_49_11), .o(n_3880) );
in01f80 g566264 ( .a(n_8612), .o(n_4777) );
oa22f80 g566265 ( .a(n_1164), .b(x_in_29_15), .c(n_2327), .d(x_in_29_12), .o(n_8612) );
in01f80 g566266 ( .a(n_3510), .o(n_2935) );
oa22f80 g566267 ( .a(n_1913), .b(x_in_49_3), .c(n_3238), .d(x_in_49_2), .o(n_3510) );
ao22s80 g566268 ( .a(n_2448), .b(x_in_47_10), .c(n_11034), .d(x_in_47_13), .o(n_6095) );
ao22s80 g566269 ( .a(n_2523), .b(x_in_63_10), .c(n_11696), .d(x_in_63_13), .o(n_6119) );
in01f80 g566270 ( .a(n_5320), .o(n_4683) );
oa22f80 g566271 ( .a(n_2329), .b(x_in_33_4), .c(n_5281), .d(x_in_33_3), .o(n_5320) );
ao22s80 g566272 ( .a(n_2575), .b(x_in_15_10), .c(n_11037), .d(x_in_15_13), .o(n_5763) );
in01f80 g566273 ( .a(n_5322), .o(n_2934) );
oa22f80 g566274 ( .a(n_2488), .b(x_in_9_14), .c(n_2376), .d(x_in_9_11), .o(n_5322) );
ao22s80 g566275 ( .a(n_2533), .b(x_in_33_11), .c(n_12178), .d(x_in_33_13), .o(n_4793) );
in01f80 g566276 ( .a(FE_OFN676_n_6824), .o(n_2775) );
ao22s80 g566277 ( .a(n_2492), .b(x_in_25_13), .c(n_5311), .d(x_in_25_14), .o(n_6824) );
ao22s80 g566278 ( .a(n_2533), .b(x_in_33_12), .c(n_12635), .d(x_in_33_13), .o(n_3636) );
in01f80 g566279 ( .a(n_5377), .o(n_4627) );
oa22f80 g566280 ( .a(n_6488), .b(x_in_23_14), .c(n_16158), .d(x_in_23_13), .o(n_5377) );
in01f80 g566281 ( .a(n_4919), .o(n_4624) );
oa22f80 g566282 ( .a(n_7231), .b(x_in_55_14), .c(n_16156), .d(x_in_55_13), .o(n_4919) );
in01f80 g566283 ( .a(FE_OFN646_n_6732), .o(n_4630) );
oa22f80 g566284 ( .a(n_2310), .b(x_in_21_15), .c(n_2309), .d(x_in_21_13), .o(n_6732) );
in01f80 g566285 ( .a(n_5299), .o(n_3435) );
no02f80 g566286 ( .a(n_2140), .b(n_2067), .o(n_5299) );
in01f80 g566287 ( .a(n_5353), .o(n_4248) );
oa22f80 g566288 ( .a(n_7291), .b(x_in_31_14), .c(n_16154), .d(x_in_31_13), .o(n_5353) );
oa22f80 g566289 ( .a(n_2445), .b(x_in_59_4), .c(n_5271), .d(x_in_59_2), .o(n_3457) );
in01f80 g566290 ( .a(n_3602), .o(n_2812) );
oa22f80 g566291 ( .a(n_2061), .b(x_in_35_4), .c(n_5987), .d(x_in_35_2), .o(n_3602) );
in01f80 g566292 ( .a(FE_OFN1202_n_5312), .o(n_2818) );
ao22s80 g566293 ( .a(n_2421), .b(x_in_27_1), .c(n_2420), .d(x_in_27_3), .o(n_5312) );
ao22s80 g566294 ( .a(n_4687), .b(x_in_17_1), .c(n_3363), .d(x_in_17_2), .o(n_8287) );
in01f80 g566295 ( .a(n_4823), .o(n_2933) );
oa22f80 g566296 ( .a(n_2424), .b(x_in_41_5), .c(n_2583), .d(x_in_41_3), .o(n_4823) );
oa22f80 g566297 ( .a(n_2699), .b(x_in_7_4), .c(n_8522), .d(x_in_7_2), .o(n_3952) );
oa22f80 g566298 ( .a(n_2520), .b(x_in_17_6), .c(n_5362), .d(x_in_17_3), .o(n_5453) );
in01f80 g566299 ( .a(n_5261), .o(n_5260) );
oa22f80 g566300 ( .a(n_2440), .b(x_in_19_4), .c(n_5939), .d(x_in_19_2), .o(n_5261) );
oa22f80 g566301 ( .a(n_11041), .b(x_in_23_13), .c(n_6488), .d(x_in_23_10), .o(n_6064) );
ao22s80 g566302 ( .a(n_7291), .b(x_in_31_10), .c(n_11698), .d(x_in_31_13), .o(n_6133) );
ao22s80 g566303 ( .a(n_7231), .b(x_in_55_10), .c(n_11040), .d(x_in_55_13), .o(n_5720) );
in01f80 g566304 ( .a(n_3425), .o(n_6390) );
oa22f80 g566305 ( .a(n_4343), .b(x_in_37_15), .c(n_3241), .d(x_in_37_13), .o(n_3425) );
ao22s80 g566306 ( .a(n_2691), .b(x_in_49_12), .c(n_2737), .d(x_in_49_13), .o(n_3912) );
ao22s80 g566307 ( .a(n_2452), .b(x_in_33_0), .c(n_2636), .d(x_in_33_1), .o(n_3527) );
ao22s80 g566308 ( .a(n_6483), .b(x_in_31_3), .c(n_2721), .d(x_in_31_6), .o(n_6317) );
oa22f80 g566309 ( .a(n_3075), .b(x_in_23_6), .c(n_6689), .d(x_in_23_3), .o(n_5450) );
oa22f80 g566310 ( .a(n_2828), .b(x_in_63_6), .c(n_6711), .d(x_in_63_3), .o(n_5447) );
oa22f80 g566311 ( .a(n_3079), .b(x_in_55_6), .c(n_6685), .d(x_in_55_3), .o(n_4905) );
ao22s80 g566312 ( .a(n_6683), .b(x_in_47_3), .c(n_2747), .d(x_in_47_6), .o(n_5777) );
oa22f80 g566313 ( .a(n_2780), .b(x_in_15_6), .c(n_6687), .d(x_in_15_3), .o(n_5456) );
ao22s80 g566314 ( .a(n_23944), .b(x_in_5_13), .c(n_13241), .d(x_in_5_15), .o(n_6701) );
in01f80 g566315 ( .a(n_4040), .o(n_4041) );
na02f80 g566316 ( .a(n_2041), .b(n_2120), .o(n_4040) );
in01f80 g566317 ( .a(n_6740), .o(n_3017) );
ao22s80 g566318 ( .a(n_3193), .b(x_in_53_13), .c(n_5988), .d(x_in_53_15), .o(n_6740) );
in01f80 g566319 ( .a(n_5417), .o(n_3550) );
na02f80 g566320 ( .a(n_2271), .b(n_2270), .o(n_5417) );
in01f80 g566321 ( .a(n_10431), .o(n_10426) );
oa22f80 g566322 ( .a(n_2673), .b(x_in_13_14), .c(n_3077), .d(x_in_13_10), .o(n_10431) );
in01f80 g566323 ( .a(n_5871), .o(n_3606) );
na02f80 g566324 ( .a(n_2101), .b(n_2093), .o(n_5871) );
oa22f80 g566325 ( .a(n_2541), .b(x_in_43_5), .c(n_3176), .d(x_in_43_3), .o(n_3502) );
oa22f80 g566326 ( .a(n_4042), .b(x_in_53_2), .c(n_2231), .d(x_in_53_0), .o(n_3918) );
oa22f80 g566327 ( .a(n_4143), .b(x_in_61_4), .c(n_8929), .d(x_in_61_2), .o(n_3907) );
in01f80 g566328 ( .a(n_3793), .o(n_2932) );
ao22s80 g566329 ( .a(n_5979), .b(x_in_51_2), .c(n_2490), .d(x_in_51_4), .o(n_3793) );
ao22s80 g566330 ( .a(n_2635), .b(x_in_59_12), .c(n_4992), .d(x_in_59_13), .o(n_3889) );
oa22f80 g566331 ( .a(n_5387), .b(x_in_11_6), .c(n_5309), .d(x_in_11_4), .o(n_3513) );
oa22f80 g566332 ( .a(n_5872), .b(x_in_21_12), .c(n_5977), .d(x_in_21_11), .o(n_5425) );
oa22f80 g566333 ( .a(n_2431), .b(x_in_11_5), .c(n_2430), .d(x_in_11_3), .o(n_3936) );
in01f80 g566334 ( .a(n_8569), .o(n_4977) );
no02f80 g566335 ( .a(n_2286), .b(n_2242), .o(n_8569) );
in01f80 g566336 ( .a(FE_OFN845_n_7616), .o(n_3181) );
oa22f80 g566337 ( .a(n_2049), .b(x_in_45_14), .c(n_2326), .d(x_in_45_11), .o(n_7616) );
ao22s80 g566338 ( .a(n_11041), .b(x_in_23_7), .c(n_7906), .d(x_in_23_10), .o(n_6187) );
ao22s80 g566339 ( .a(n_11040), .b(x_in_55_7), .c(n_7905), .d(x_in_55_10), .o(n_6178) );
ao22s80 g566340 ( .a(n_11698), .b(x_in_31_7), .c(n_7902), .d(x_in_31_10), .o(n_6017) );
ao22s80 g566341 ( .a(n_11034), .b(x_in_47_7), .c(n_7901), .d(x_in_47_10), .o(n_6052) );
ao22s80 g566342 ( .a(n_11696), .b(x_in_63_7), .c(n_7903), .d(x_in_63_10), .o(n_6110) );
ao22s80 g566343 ( .a(n_11037), .b(x_in_15_7), .c(n_7904), .d(x_in_15_10), .o(n_6184) );
oa22f80 g566344 ( .a(n_5390), .b(x_in_35_5), .c(n_2377), .d(x_in_35_3), .o(n_4956) );
in01f80 g566345 ( .a(n_2930), .o(n_2931) );
oa22f80 g566346 ( .a(n_2363), .b(x_in_59_11), .c(n_8482), .d(x_in_59_9), .o(n_2930) );
in01f80 g566347 ( .a(FE_OFN674_n_6720), .o(n_2929) );
ao22s80 g566348 ( .a(n_2546), .b(x_in_25_11), .c(n_3189), .d(x_in_25_15), .o(n_6720) );
in01f80 g566349 ( .a(n_5286), .o(n_5287) );
oa22f80 g566350 ( .a(n_5987), .b(x_in_35_6), .c(n_5369), .d(x_in_35_4), .o(n_5286) );
oa22f80 g566351 ( .a(n_5271), .b(x_in_59_6), .c(n_5275), .d(x_in_59_4), .o(n_3418) );
ao22s80 g566352 ( .a(n_3641), .b(x_in_57_13), .c(n_3560), .d(x_in_57_15), .o(n_6707) );
in01f80 g566353 ( .a(n_3538), .o(n_2731) );
oa22f80 g566354 ( .a(n_5302), .b(x_in_57_13), .c(n_3560), .d(x_in_57_12), .o(n_3538) );
in01f80 g566355 ( .a(FE_OFN1274_n_8977), .o(n_4652) );
ao22s80 g566356 ( .a(n_2518), .b(x_in_61_12), .c(n_2353), .d(x_in_61_13), .o(n_8977) );
ao22s80 g566357 ( .a(n_6420), .b(x_in_51_11), .c(n_8420), .d(x_in_51_12), .o(n_4950) );
in01f80 g566358 ( .a(n_3213), .o(n_3214) );
oa22f80 g566359 ( .a(n_3229), .b(x_in_11_12), .c(n_5025), .d(x_in_11_10), .o(n_3213) );
oa22f80 g566360 ( .a(n_2522), .b(x_in_13_10), .c(n_2673), .d(x_in_13_8), .o(n_6373) );
oa22f80 g566361 ( .a(n_3833), .b(x_in_61_12), .c(n_2353), .d(x_in_61_10), .o(n_3894) );
in01f80 g566362 ( .a(FE_OFN1091_n_8621), .o(n_4915) );
ao22s80 g566363 ( .a(n_2353), .b(x_in_61_11), .c(n_4529), .d(x_in_61_12), .o(n_8621) );
oa22f80 g566364 ( .a(n_4180), .b(x_in_37_12), .c(n_5849), .d(x_in_37_11), .o(n_3932) );
in01f80 g566365 ( .a(n_6435), .o(n_5132) );
oa22f80 g566366 ( .a(n_4825), .b(x_in_53_5), .c(n_2626), .d(x_in_53_1), .o(n_6435) );
oa22f80 g566367 ( .a(n_2421), .b(x_in_27_5), .c(n_3747), .d(x_in_27_3), .o(n_3940) );
in01f80 g566368 ( .a(n_2927), .o(n_2928) );
oa22f80 g566369 ( .a(n_5256), .b(x_in_7_7), .c(n_6494), .d(x_in_7_5), .o(n_2927) );
in01f80 g566370 ( .a(n_5345), .o(n_5347) );
oa22f80 g566371 ( .a(n_5252), .b(x_in_19_5), .c(n_3174), .d(x_in_19_3), .o(n_5345) );
in01f80 g566372 ( .a(n_3226), .o(n_3227) );
oa22f80 g566373 ( .a(n_5310), .b(x_in_11_11), .c(n_7818), .d(x_in_11_9), .o(n_3226) );
oa22f80 g566374 ( .a(n_2521), .b(x_in_13_11), .c(n_482), .d(x_in_13_9), .o(n_6136) );
ao22s80 g566375 ( .a(n_2506), .b(x_in_13_4), .c(n_2433), .d(x_in_13_6), .o(n_6122) );
oa22f80 g566376 ( .a(n_2540), .b(x_in_5_4), .c(n_2517), .d(x_in_5_3), .o(n_6826) );
oa22f80 g566377 ( .a(n_8482), .b(x_in_59_12), .c(n_4992), .d(x_in_59_11), .o(n_4364) );
ao22s80 g566378 ( .a(n_8482), .b(x_in_59_10), .c(n_2668), .d(x_in_59_11), .o(n_4817) );
in01f80 g566379 ( .a(n_4941), .o(n_4940) );
oa22f80 g566380 ( .a(n_5098), .b(x_in_35_11), .c(n_8524), .d(x_in_35_9), .o(n_4941) );
in01f80 g566381 ( .a(n_4594), .o(n_3290) );
oa22f80 g566382 ( .a(n_2554), .b(x_in_25_7), .c(n_3132), .d(x_in_25_4), .o(n_4594) );
ao22s80 g566383 ( .a(n_3186), .b(x_in_49_10), .c(n_3187), .d(x_in_49_11), .o(n_3653) );
in01f80 g566384 ( .a(n_9520), .o(n_4702) );
oa22f80 g566385 ( .a(n_7340), .b(x_in_7_13), .c(n_7285), .d(x_in_7_12), .o(n_9520) );
ao22s80 g566386 ( .a(n_8557), .b(x_in_21_3), .c(n_6781), .d(x_in_21_4), .o(n_7641) );
in01f80 g566387 ( .a(n_3998), .o(n_3205) );
oa22f80 g566388 ( .a(n_2516), .b(x_in_13_5), .c(n_2505), .d(x_in_13_3), .o(n_3998) );
in01f80 g566389 ( .a(FE_OFN1188_n_5249), .o(n_5248) );
oa22f80 g566390 ( .a(n_2699), .b(x_in_7_3), .c(n_5272), .d(x_in_7_2), .o(n_5249) );
in01f80 g566391 ( .a(n_8021), .o(n_4660) );
oa22f80 g566392 ( .a(n_5988), .b(x_in_53_14), .c(n_2762), .d(x_in_53_13), .o(n_8021) );
oa22f80 g566393 ( .a(n_2673), .b(x_in_13_12), .c(n_5926), .d(x_in_13_10), .o(n_6139) );
ao22s80 g566394 ( .a(n_4654), .b(x_in_37_2), .c(n_3011), .d(x_in_37_3), .o(n_4862) );
in01f80 g566395 ( .a(n_5329), .o(n_5330) );
ao22s80 g566396 ( .a(n_3792), .b(x_in_51_3), .c(n_5180), .d(x_in_51_5), .o(n_5329) );
in01f80 g566397 ( .a(n_3548), .o(n_3337) );
oa22f80 g566398 ( .a(n_5313), .b(x_in_57_12), .c(n_5302), .d(x_in_57_11), .o(n_3548) );
in01f80 g566399 ( .a(n_8029), .o(n_4264) );
oa22f80 g566400 ( .a(n_5317), .b(x_in_25_13), .c(n_5311), .d(x_in_25_12), .o(n_8029) );
in01f80 g566401 ( .a(n_5057), .o(n_2925) );
ao22s80 g566402 ( .a(n_3129), .b(x_in_25_5), .c(n_4593), .d(x_in_25_8), .o(n_5057) );
in01f80 g566403 ( .a(n_2923), .o(n_2924) );
oa22f80 g566404 ( .a(n_3237), .b(x_in_61_5), .c(n_5242), .d(x_in_61_1), .o(n_2923) );
oa22f80 g566405 ( .a(n_2517), .b(x_in_5_5), .c(n_5296), .d(x_in_5_4), .o(n_4872) );
oa22f80 g566406 ( .a(n_5679), .b(x_in_27_6), .c(n_5677), .d(x_in_27_4), .o(n_3778) );
oa22f80 g566407 ( .a(n_2452), .b(x_in_33_2), .c(n_2451), .d(x_in_33_1), .o(n_6828) );
oa22f80 g566408 ( .a(n_2451), .b(x_in_33_3), .c(n_2329), .d(x_in_33_2), .o(n_4820) );
in01f80 g566409 ( .a(FE_OFN973_n_6822), .o(n_4902) );
ao22s80 g566410 ( .a(n_5988), .b(x_in_53_12), .c(n_2548), .d(x_in_53_13), .o(n_6822) );
in01f80 g566411 ( .a(n_4841), .o(n_3347) );
oa22f80 g566412 ( .a(n_5332), .b(x_in_51_11), .c(n_8420), .d(x_in_51_9), .o(n_4841) );
in01f80 g566413 ( .a(n_2890), .o(n_2891) );
oa22f80 g566414 ( .a(n_7417), .b(x_in_27_12), .c(n_7402), .d(x_in_27_10), .o(n_2890) );
in01f80 g566415 ( .a(n_2920), .o(n_2921) );
oa22f80 g566416 ( .a(n_6496), .b(x_in_43_12), .c(n_7263), .d(x_in_43_10), .o(n_2920) );
in01f80 g566417 ( .a(n_5099), .o(n_2919) );
ao22s80 g566418 ( .a(n_5032), .b(x_in_35_10), .c(n_2652), .d(x_in_35_12), .o(n_5099) );
ao22s80 g566419 ( .a(n_7905), .b(x_in_55_4), .c(n_3742), .d(x_in_55_7), .o(n_6175) );
ao22s80 g566420 ( .a(n_7904), .b(x_in_15_4), .c(n_3482), .d(x_in_15_7), .o(n_6438) );
ao22s80 g566421 ( .a(n_7903), .b(x_in_63_4), .c(n_3737), .d(x_in_63_7), .o(n_6098) );
ao22s80 g566422 ( .a(n_7901), .b(x_in_47_4), .c(n_3445), .d(x_in_47_7), .o(n_6172) );
ao22s80 g566423 ( .a(n_7902), .b(x_in_31_4), .c(n_3739), .d(x_in_31_7), .o(n_6193) );
oa22f80 g566424 ( .a(n_3744), .b(x_in_23_7), .c(n_7906), .d(x_in_23_4), .o(n_6190) );
in01f80 g566425 ( .a(n_2917), .o(n_2918) );
oa22f80 g566426 ( .a(n_2430), .b(x_in_11_7), .c(n_5089), .d(x_in_11_5), .o(n_2917) );
oa22f80 g566427 ( .a(n_5293), .b(x_in_43_6), .c(n_5327), .d(x_in_43_4), .o(n_3920) );
in01f80 g566428 ( .a(n_8454), .o(n_8880) );
oa22f80 g566429 ( .a(n_4593), .b(x_in_25_6), .c(n_3771), .d(x_in_25_5), .o(n_8454) );
in01f80 g566430 ( .a(n_2787), .o(n_2788) );
oa22f80 g566431 ( .a(n_7289), .b(x_in_27_11), .c(n_8513), .d(x_in_27_9), .o(n_2787) );
in01f80 g566432 ( .a(n_2756), .o(n_2757) );
oa22f80 g566433 ( .a(n_7268), .b(x_in_43_11), .c(n_8443), .d(x_in_43_9), .o(n_2756) );
oa22f80 g566434 ( .a(n_2657), .b(x_in_13_9), .c(n_2521), .d(x_in_13_7), .o(n_6125) );
oa22f80 g566435 ( .a(n_2505), .b(x_in_13_7), .c(n_2657), .d(x_in_13_5), .o(n_6058) );
ao22s80 g566436 ( .a(n_2522), .b(x_in_13_6), .c(n_2506), .d(x_in_13_8), .o(n_6072) );
in01f80 g566437 ( .a(n_3981), .o(n_2782) );
oa22f80 g566438 ( .a(n_3409), .b(x_in_57_11), .c(n_5313), .d(x_in_57_10), .o(n_3981) );
in01f80 g566439 ( .a(n_7477), .o(n_2736) );
ao22s80 g566440 ( .a(n_2546), .b(x_in_25_13), .c(n_5311), .d(x_in_25_15), .o(n_7477) );
in01f80 g566441 ( .a(n_2783), .o(n_2784) );
oa22f80 g566442 ( .a(n_7320), .b(x_in_7_11), .c(n_7336), .d(x_in_7_9), .o(n_2783) );
in01f80 g566443 ( .a(n_5285), .o(n_2915) );
ao22s80 g566444 ( .a(n_5311), .b(x_in_25_10), .c(n_2743), .d(x_in_25_13), .o(n_5285) );
ao22s80 g566445 ( .a(n_7332), .b(x_in_55_8), .c(n_7315), .d(x_in_55_11), .o(n_6083) );
ao22s80 g566446 ( .a(n_7334), .b(x_in_15_8), .c(n_6492), .d(x_in_15_11), .o(n_6164) );
in01f80 g566447 ( .a(n_2913), .o(n_2914) );
oa22f80 g566448 ( .a(n_7298), .b(x_in_31_12), .c(n_6753), .d(x_in_31_11), .o(n_2913) );
oa22f80 g566449 ( .a(n_8200), .b(x_in_31_11), .c(n_7298), .d(x_in_31_8), .o(n_6075) );
in01f80 g566450 ( .a(n_2825), .o(n_2826) );
oa22f80 g566451 ( .a(n_7334), .b(x_in_15_12), .c(n_7338), .d(x_in_15_11), .o(n_2825) );
ao22s80 g566452 ( .a(n_8200), .b(x_in_31_5), .c(n_4738), .d(x_in_31_8), .o(n_6128) );
in01f80 g566453 ( .a(n_2911), .o(n_2912) );
oa22f80 g566454 ( .a(n_7308), .b(x_in_63_12), .c(n_8206), .d(x_in_63_11), .o(n_2911) );
ao22s80 g566455 ( .a(n_7241), .b(x_in_47_5), .c(n_4737), .d(x_in_47_8), .o(n_6145) );
ao22s80 g566456 ( .a(n_7296), .b(x_in_23_8), .c(n_7270), .d(x_in_23_11), .o(n_6161) );
in01f80 g566457 ( .a(n_2909), .o(n_2910) );
oa22f80 g566458 ( .a(n_7296), .b(x_in_23_12), .c(n_7323), .d(x_in_23_11), .o(n_2909) );
ao22s80 g566459 ( .a(n_7245), .b(x_in_47_8), .c(n_7241), .d(x_in_47_11), .o(n_6151) );
in01f80 g566460 ( .a(n_2711), .o(n_2712) );
oa22f80 g566461 ( .a(n_7245), .b(x_in_47_12), .c(n_7247), .d(x_in_47_11), .o(n_2711) );
ao22s80 g566462 ( .a(n_7308), .b(x_in_63_8), .c(n_7272), .d(x_in_63_11), .o(n_6113) );
in01f80 g566463 ( .a(n_3303), .o(n_3304) );
oa22f80 g566464 ( .a(n_7332), .b(x_in_55_12), .c(n_7278), .d(x_in_55_11), .o(n_3303) );
in01f80 g566465 ( .a(n_6856), .o(n_5246) );
ao22s80 g566466 ( .a(n_2870), .b(x_in_53_10), .c(n_2653), .d(x_in_53_11), .o(n_6856) );
in01f80 g566467 ( .a(FE_OFN1254_n_12186), .o(n_3053) );
ao22s80 g566468 ( .a(n_2762), .b(x_in_53_10), .c(n_2653), .d(x_in_53_14), .o(n_12186) );
in01f80 g566469 ( .a(n_4944), .o(n_4943) );
oa22f80 g566470 ( .a(n_4939), .b(x_in_35_10), .c(n_2652), .d(x_in_35_8), .o(n_4944) );
in01f80 g566471 ( .a(n_2907), .o(n_2908) );
oa22f80 g566472 ( .a(n_3259), .b(x_in_59_7), .c(n_5699), .d(x_in_59_5), .o(n_2907) );
oa22f80 g566474 ( .a(n_4143), .b(x_in_61_3), .c(n_3608), .d(x_in_61_2), .o(n_6399) );
oa22f80 g566475 ( .a(n_5275), .b(x_in_59_8), .c(n_5691), .d(x_in_59_6), .o(n_3824) );
in01f80 g566476 ( .a(n_2726), .o(n_2727) );
oa22f80 g566477 ( .a(n_3176), .b(x_in_43_7), .c(n_5519), .d(x_in_43_5), .o(n_2726) );
in01f80 g566478 ( .a(n_3983), .o(n_3216) );
oa22f80 g566479 ( .a(n_3245), .b(x_in_57_10), .c(n_3409), .d(x_in_57_9), .o(n_3983) );
in01f80 g566480 ( .a(n_3183), .o(n_3184) );
oa22f80 g566481 ( .a(n_5691), .b(x_in_59_10), .c(n_2668), .d(x_in_59_8), .o(n_3183) );
in01f80 g566482 ( .a(n_4936), .o(n_3182) );
oa22f80 g566483 ( .a(n_5979), .b(x_in_51_6), .c(n_6350), .d(x_in_51_4), .o(n_4936) );
in01f80 g566484 ( .a(FE_OFN1250_n_5334), .o(n_5333) );
oa22f80 g566485 ( .a(n_5283), .b(x_in_51_12), .c(n_6420), .d(x_in_51_10), .o(n_5334) );
oa22f80 g566486 ( .a(n_5677), .b(x_in_27_8), .c(n_7287), .d(x_in_27_6), .o(n_3897) );
in01f80 g566487 ( .a(n_5367), .o(n_2905) );
ao22s80 g566488 ( .a(n_4942), .b(x_in_35_5), .c(n_2377), .d(x_in_35_7), .o(n_5367) );
oa22f80 g566489 ( .a(n_3260), .b(x_in_59_5), .c(n_3259), .d(x_in_59_3), .o(n_5269) );
in01f80 g566490 ( .a(n_2849), .o(n_2850) );
oa22f80 g566491 ( .a(n_5519), .b(x_in_43_9), .c(n_7268), .d(x_in_43_7), .o(n_2849) );
in01f80 g566492 ( .a(n_5704), .o(n_4662) );
oa22f80 g566493 ( .a(n_2554), .b(x_in_25_5), .c(n_4593), .d(x_in_25_4), .o(n_5704) );
in01f80 g566494 ( .a(n_5366), .o(n_2904) );
oa22f80 g566495 ( .a(n_2385), .b(x_in_45_5), .c(n_2438), .d(x_in_45_1), .o(n_5366) );
oa22f80 g566496 ( .a(n_5309), .b(x_in_11_8), .c(n_5352), .d(x_in_11_6), .o(n_4084) );
in01f80 g566497 ( .a(n_2902), .o(n_2903) );
oa22f80 g566498 ( .a(n_5352), .b(x_in_11_10), .c(n_3229), .d(x_in_11_8), .o(n_2902) );
in01f80 g566499 ( .a(n_2717), .o(n_2718) );
oa22f80 g566500 ( .a(n_5089), .b(x_in_11_9), .c(n_5310), .d(x_in_11_7), .o(n_2717) );
ao22s80 g566501 ( .a(n_4180), .b(x_in_37_10), .c(n_5745), .d(x_in_37_11), .o(n_3622) );
in01f80 g566502 ( .a(n_8674), .o(n_3320) );
ao22s80 g566503 ( .a(n_7340), .b(x_in_7_11), .c(n_7336), .d(x_in_7_12), .o(n_8674) );
in01f80 g566504 ( .a(FE_OFN971_n_6854), .o(n_5239) );
ao22s80 g566505 ( .a(n_2548), .b(x_in_53_11), .c(n_2870), .d(x_in_53_12), .o(n_6854) );
oa22f80 g566506 ( .a(n_8165), .b(x_in_7_11), .c(n_7336), .d(x_in_7_10), .o(n_9082) );
in01f80 g566507 ( .a(n_3217), .o(n_3218) );
oa22f80 g566508 ( .a(n_3747), .b(x_in_27_7), .c(n_5680), .d(x_in_27_5), .o(n_3217) );
ao22s80 g566509 ( .a(n_12178), .b(x_in_33_10), .c(n_12634), .d(x_in_33_11), .o(n_3891) );
ao22s80 g566510 ( .a(n_7247), .b(x_in_47_9), .c(n_10913), .d(x_in_47_12), .o(n_6154) );
ao22s80 g566511 ( .a(n_6492), .b(x_in_15_5), .c(n_4746), .d(x_in_15_8), .o(n_6142) );
ao22s80 g566512 ( .a(n_10918), .b(x_in_23_6), .c(n_6689), .d(x_in_23_9), .o(n_6055) );
ao22s80 g566513 ( .a(n_3191), .b(x_in_49_8), .c(n_3188), .d(x_in_49_9), .o(n_3726) );
ao22s80 g566514 ( .a(n_7278), .b(x_in_55_9), .c(n_10915), .d(x_in_55_12), .o(n_6197) );
ao22s80 g566515 ( .a(n_7315), .b(x_in_55_5), .c(n_4329), .d(x_in_55_8), .o(n_6061) );
ao22s80 g566516 ( .a(n_6753), .b(x_in_31_9), .c(n_10914), .d(x_in_31_12), .o(n_6444) );
ao22s80 g566517 ( .a(n_7272), .b(x_in_63_5), .c(n_4745), .d(x_in_63_8), .o(n_6101) );
ao22s80 g566518 ( .a(n_7323), .b(x_in_23_9), .c(n_10918), .d(x_in_23_12), .o(n_6078) );
ao22s80 g566519 ( .a(n_8206), .b(x_in_63_9), .c(n_10916), .d(x_in_63_12), .o(n_6104) );
ao22s80 g566520 ( .a(n_7270), .b(x_in_23_5), .c(n_4744), .d(x_in_23_8), .o(n_5713) );
ao22s80 g566521 ( .a(n_10917), .b(x_in_15_6), .c(n_6687), .d(x_in_15_9), .o(n_6026) );
ao22s80 g566522 ( .a(n_2588), .b(x_in_49_5), .c(n_5095), .d(x_in_49_6), .o(n_3613) );
ao22s80 g566523 ( .a(n_2589), .b(x_in_49_6), .c(n_2588), .d(x_in_49_7), .o(n_3925) );
oa22f80 g566524 ( .a(n_6711), .b(x_in_63_9), .c(n_10916), .d(x_in_63_6), .o(n_6107) );
ao22s80 g566525 ( .a(n_7338), .b(x_in_15_9), .c(n_10917), .d(x_in_15_12), .o(n_6049) );
in01f80 g566526 ( .a(n_3250), .o(n_3251) );
oa22f80 g566527 ( .a(n_2589), .b(x_in_49_8), .c(n_3188), .d(x_in_49_7), .o(n_3250) );
ao22s80 g566528 ( .a(n_10915), .b(x_in_55_6), .c(n_6685), .d(x_in_55_9), .o(n_6067) );
in01f80 g566529 ( .a(n_3916), .o(n_6820) );
oa22f80 g566530 ( .a(n_2526), .b(x_in_57_4), .c(n_2601), .d(x_in_57_3), .o(n_3916) );
ao22s80 g566531 ( .a(n_3187), .b(x_in_49_9), .c(n_3191), .d(x_in_49_10), .o(n_3584) );
oa22f80 g566532 ( .a(n_6483), .b(x_in_31_9), .c(n_10914), .d(x_in_31_6), .o(n_6315) );
oa22f80 g566533 ( .a(n_6683), .b(x_in_47_9), .c(n_10913), .d(x_in_47_6), .o(n_6148) );
in01f80 g566534 ( .a(n_8036), .o(n_4289) );
oa22f80 g566535 ( .a(n_2743), .b(x_in_25_11), .c(n_3189), .d(x_in_25_10), .o(n_8036) );
oa22f80 g566536 ( .a(n_3129), .b(x_in_25_11), .c(n_3189), .d(x_in_25_8), .o(n_4821) );
in01f80 g566537 ( .a(n_4909), .o(n_2974) );
ao22s80 g566538 ( .a(n_5317), .b(x_in_25_9), .c(n_2581), .d(x_in_25_12), .o(n_4909) );
in01f80 g566539 ( .a(n_3164), .o(n_3165) );
oa22f80 g566540 ( .a(n_5699), .b(x_in_59_9), .c(n_2363), .d(x_in_59_7), .o(n_3164) );
oa22f80 g566541 ( .a(n_4668), .b(x_in_57_6), .c(n_2512), .d(x_in_57_5), .o(n_3911) );
in01f80 g566542 ( .a(n_3985), .o(n_2872) );
oa22f80 g566543 ( .a(n_2512), .b(x_in_57_7), .c(n_4055), .d(x_in_57_6), .o(n_3985) );
in01f80 g566544 ( .a(n_3522), .o(n_2897) );
oa22f80 g566545 ( .a(n_2627), .b(x_in_57_9), .c(n_3245), .d(x_in_57_8), .o(n_3522) );
in01f80 g566546 ( .a(n_3524), .o(n_2896) );
oa22f80 g566547 ( .a(n_4055), .b(x_in_57_8), .c(n_2627), .d(x_in_57_7), .o(n_3524) );
oa22f80 g566548 ( .a(n_4914), .b(x_in_61_11), .c(n_4529), .d(x_in_61_9), .o(n_3626) );
oa22f80 g566549 ( .a(n_4937), .b(x_in_61_10), .c(n_3833), .d(x_in_61_8), .o(n_3455) );
in01f80 g566550 ( .a(n_5028), .o(n_5027) );
oa22f80 g566551 ( .a(n_4942), .b(x_in_35_9), .c(n_5098), .d(x_in_35_7), .o(n_5028) );
oa22f80 g566552 ( .a(n_2668), .b(x_in_59_12), .c(n_4992), .d(x_in_59_10), .o(n_3814) );
oa22f80 g566553 ( .a(n_5369), .b(x_in_35_8), .c(n_4939), .d(x_in_35_6), .o(n_5076) );
in01f80 g566554 ( .a(n_8065), .o(n_4755) );
oa22f80 g566555 ( .a(n_3771), .b(x_in_25_7), .c(n_3132), .d(x_in_25_6), .o(n_8065) );
in01f80 g566556 ( .a(FE_OFN1246_n_4900), .o(n_4901) );
ao22s80 g566557 ( .a(n_5331), .b(x_in_51_5), .c(n_3792), .d(x_in_51_7), .o(n_4900) );
in01f80 g566558 ( .a(n_5315), .o(n_3028) );
ao22s80 g566559 ( .a(n_2581), .b(x_in_25_6), .c(n_3771), .d(x_in_25_9), .o(n_5315) );
in01f80 g566560 ( .a(n_2893), .o(n_2894) );
oa22f80 g566561 ( .a(n_8165), .b(x_in_7_12), .c(n_7340), .d(x_in_7_10), .o(n_2893) );
oa22f80 g566562 ( .a(n_5327), .b(x_in_43_8), .c(n_5501), .d(x_in_43_6), .o(n_4025) );
in01f80 g566563 ( .a(n_3029), .o(n_3030) );
oa22f80 g566564 ( .a(n_5501), .b(x_in_43_10), .c(n_6496), .d(x_in_43_8), .o(n_3029) );
in01f80 g566565 ( .a(n_3343), .o(n_3344) );
oa22f80 g566566 ( .a(n_5680), .b(x_in_27_9), .c(n_7289), .d(x_in_27_7), .o(n_3343) );
in01f80 g566567 ( .a(n_3231), .o(n_3232) );
oa22f80 g566568 ( .a(n_7287), .b(x_in_27_10), .c(n_7417), .d(x_in_27_8), .o(n_3231) );
ao22s80 g566569 ( .a(n_12175), .b(x_in_33_7), .c(n_8885), .d(x_in_33_8), .o(n_3604) );
ao22s80 g566570 ( .a(n_8885), .b(x_in_33_6), .c(n_12172), .d(x_in_33_7), .o(n_3896) );
ao22s80 g566571 ( .a(n_8884), .b(x_in_33_8), .c(n_12175), .d(x_in_33_9), .o(n_3359) );
in01f80 g566572 ( .a(n_4927), .o(n_3159) );
oa22f80 g566573 ( .a(n_6350), .b(x_in_51_8), .c(n_6351), .d(x_in_51_6), .o(n_4927) );
in01f80 g566574 ( .a(n_5325), .o(n_5324) );
oa22f80 g566575 ( .a(n_6351), .b(x_in_51_10), .c(n_5283), .d(x_in_51_8), .o(n_5325) );
in01f80 g566576 ( .a(FE_OFN1087_n_8974), .o(n_4938) );
ao22s80 g566577 ( .a(n_4529), .b(x_in_61_10), .c(n_3833), .d(x_in_61_11), .o(n_8974) );
ao22s80 g566578 ( .a(n_12634), .b(x_in_33_9), .c(n_8884), .d(x_in_33_10), .o(n_3403) );
in01f80 g566579 ( .a(n_3551), .o(n_8047) );
oa22f80 g566580 ( .a(n_3132), .b(x_in_25_8), .c(n_3129), .d(x_in_25_7), .o(n_3551) );
in01f80 g566581 ( .a(n_3957), .o(n_8042) );
oa22f80 g566582 ( .a(n_2581), .b(x_in_25_10), .c(n_2743), .d(x_in_25_9), .o(n_3957) );
in01f80 g566583 ( .a(n_8044), .o(n_4358) );
oa22f80 g566584 ( .a(n_3129), .b(x_in_25_9), .c(n_2581), .d(x_in_25_8), .o(n_8044) );
in01f80 g566585 ( .a(FE_OFN931_n_4898), .o(n_4899) );
ao22s80 g566586 ( .a(n_5332), .b(x_in_51_7), .c(n_5331), .d(x_in_51_9), .o(n_4898) );
in01f80 g566587 ( .a(n_5316), .o(n_2725) );
ao22s80 g566588 ( .a(n_2743), .b(x_in_25_7), .c(n_3132), .d(x_in_25_10), .o(n_5316) );
in01f80 g566589 ( .a(n_8034), .o(n_4688) );
oa22f80 g566590 ( .a(n_3189), .b(x_in_25_12), .c(n_5317), .d(x_in_25_11), .o(n_8034) );
na02f80 g566591 ( .a(x_in_5_9), .b(x_in_4_5), .o(n_3224) );
na02f80 g566592 ( .a(x_in_55_0), .b(x_in_55_3), .o(n_7980) );
na02f80 g566593 ( .a(x_in_1_12), .b(x_in_0_12), .o(n_3060) );
na02f80 g566594 ( .a(x_in_15_0), .b(x_in_15_3), .o(n_7991) );
na02f80 g566595 ( .a(x_in_1_5), .b(x_in_0_5), .o(n_3153) );
na02f80 g566596 ( .a(x_in_9_3), .b(x_in_9_0), .o(n_7195) );
in01f80 g566597 ( .a(n_2196), .o(n_2197) );
no02f80 g566598 ( .a(x_in_57_15), .b(x_in_56_14), .o(n_2196) );
in01f80 g566599 ( .a(n_2194), .o(n_2195) );
no02f80 g566600 ( .a(x_in_5_12), .b(x_in_4_8), .o(n_2194) );
na02f80 g566601 ( .a(x_in_5_12), .b(x_in_4_8), .o(n_2874) );
na02f80 g566602 ( .a(x_in_41_15), .b(x_in_40_14), .o(n_2709) );
in01f80 g566603 ( .a(n_2192), .o(n_2193) );
no02f80 g566604 ( .a(x_in_5_7), .b(x_in_4_3), .o(n_2192) );
na02f80 g566605 ( .a(x_in_1_4), .b(x_in_0_4), .o(n_2704) );
na02f80 g566606 ( .a(x_in_5_14), .b(x_in_4_10), .o(n_3230) );
in01f80 g566607 ( .a(n_2190), .o(n_2191) );
no02f80 g566608 ( .a(x_in_5_11), .b(x_in_4_7), .o(n_2190) );
na02f80 g566609 ( .a(x_in_5_13), .b(x_in_4_9), .o(n_2748) );
na02f80 g566610 ( .a(x_in_25_0), .b(x_in_25_2), .o(n_4017) );
na02f80 g566611 ( .a(x_in_31_0), .b(x_in_31_3), .o(n_7978) );
in01f80 g566612 ( .a(n_2188), .o(n_2189) );
no02f80 g566613 ( .a(x_in_1_4), .b(x_in_0_4), .o(n_2188) );
na02f80 g566614 ( .a(x_in_4_0), .b(x_in_5_4), .o(n_7099) );
na02f80 g566615 ( .a(x_in_5_8), .b(x_in_4_4), .o(n_3271) );
in01f80 g566616 ( .a(n_2186), .o(n_2187) );
no02f80 g566617 ( .a(x_in_1_3), .b(x_in_0_3), .o(n_2186) );
na02f80 g566618 ( .a(n_2517), .b(n_63), .o(n_2185) );
in01f80 g566619 ( .a(n_2183), .o(n_2184) );
no02f80 g566620 ( .a(x_in_1_7), .b(x_in_0_7), .o(n_2183) );
in01f80 g566621 ( .a(n_2181), .o(n_2182) );
no02f80 g566622 ( .a(x_in_5_8), .b(x_in_4_4), .o(n_2181) );
in01f80 g566623 ( .a(n_2179), .o(n_2180) );
no02f80 g566624 ( .a(x_in_5_14), .b(x_in_4_10), .o(n_2179) );
in01f80 g566625 ( .a(n_2250), .o(n_2251) );
no02f80 g566626 ( .a(x_in_1_11), .b(x_in_0_11), .o(n_2250) );
na02f80 g566627 ( .a(x_in_0_0), .b(x_in_1_0), .o(n_7102) );
in01f80 g566628 ( .a(n_2177), .o(n_2178) );
no02f80 g566629 ( .a(x_in_1_10), .b(x_in_0_10), .o(n_2177) );
in01f80 g566630 ( .a(n_2175), .o(n_2176) );
no02f80 g566631 ( .a(x_in_1_14), .b(x_in_0_14), .o(n_2175) );
in01f80 g566632 ( .a(n_2173), .o(n_2174) );
no02f80 g566633 ( .a(x_in_1_5), .b(x_in_0_5), .o(n_2173) );
na02f80 g566634 ( .a(x_in_0_15), .b(x_in_1_15), .o(n_2013) );
no02f80 g566635 ( .a(x_in_57_15), .b(x_in_56_13), .o(n_3267) );
na02f80 g566636 ( .a(x_in_5_15), .b(x_in_4_11), .o(n_3249) );
na02f80 g566637 ( .a(x_in_13_2), .b(x_in_13_0), .o(n_7987) );
in01f80 g566638 ( .a(n_2171), .o(n_2172) );
na02f80 g566639 ( .a(x_in_5_6), .b(x_in_4_2), .o(n_2171) );
in01f80 g566640 ( .a(n_2169), .o(n_2170) );
no02f80 g566641 ( .a(x_in_5_10), .b(x_in_4_6), .o(n_2169) );
in01f80 g566642 ( .a(n_2227), .o(n_2228) );
no02f80 g566643 ( .a(x_in_25_15), .b(x_in_24_14), .o(n_2227) );
na02f80 g566644 ( .a(x_in_63_0), .b(x_in_63_3), .o(n_7985) );
na02f80 g566645 ( .a(x_in_57_15), .b(x_in_56_14), .o(n_3247) );
in01f80 g566646 ( .a(n_2257), .o(n_2258) );
no02f80 g566647 ( .a(x_in_1_8), .b(x_in_0_8), .o(n_2257) );
na02f80 g566648 ( .a(x_in_1_14), .b(x_in_0_14), .o(n_2703) );
na02f80 g566649 ( .a(x_in_23_0), .b(x_in_23_3), .o(n_7995) );
in01f80 g566650 ( .a(n_2166), .o(n_2167) );
no02f80 g566651 ( .a(x_in_1_9), .b(x_in_0_9), .o(n_2166) );
na02f80 g566652 ( .a(x_in_1_8), .b(x_in_0_8), .o(n_3254) );
na02f80 g566653 ( .a(x_in_1_6), .b(x_in_0_6), .o(n_3160) );
in01f80 g566654 ( .a(n_2164), .o(n_2165) );
no02f80 g566655 ( .a(x_in_1_12), .b(x_in_0_12), .o(n_2164) );
na02f80 g566656 ( .a(x_in_1_13), .b(x_in_0_13), .o(n_3154) );
na02f80 g566657 ( .a(x_in_49_15), .b(x_in_48_15), .o(n_1997) );
in01f80 g566658 ( .a(n_2162), .o(n_2163) );
no02f80 g566659 ( .a(x_in_5_13), .b(x_in_4_9), .o(n_2162) );
na02f80 g566660 ( .a(x_in_41_15), .b(x_in_40_15), .o(n_1992) );
in01f80 g566661 ( .a(n_7237), .o(n_2892) );
na02f80 g566662 ( .a(x_in_39_15), .b(FE_OFN35_n_15183), .o(n_7237) );
na02f80 g566663 ( .a(n_2235), .b(n_699), .o(n_2236) );
in01f80 g566664 ( .a(n_2160), .o(n_2161) );
no02f80 g566665 ( .a(x_in_5_9), .b(x_in_4_5), .o(n_2160) );
na02f80 g566666 ( .a(x_in_16_15), .b(x_in_17_15), .o(n_2025) );
na02f80 g566667 ( .a(x_in_25_15), .b(x_in_24_14), .o(n_3341) );
in01f80 g566668 ( .a(n_2158), .o(n_2159) );
na02f80 g566669 ( .a(x_in_57_15), .b(x_in_56_13), .o(n_2158) );
na02f80 g566670 ( .a(x_in_5_7), .b(x_in_4_3), .o(n_3065) );
na02f80 g566671 ( .a(x_in_1_11), .b(x_in_0_11), .o(n_3152) );
in01f80 g566672 ( .a(n_2261), .o(n_2262) );
no02f80 g566673 ( .a(x_in_5_15), .b(x_in_4_11), .o(n_2261) );
na02f80 g566674 ( .a(x_in_47_0), .b(x_in_47_3), .o(n_7989) );
na02f80 g566675 ( .a(x_in_1_9), .b(x_in_0_9), .o(n_3155) );
na02f80 g566676 ( .a(x_in_1_3), .b(x_in_0_3), .o(n_2755) );
na02f80 g566677 ( .a(x_in_5_11), .b(x_in_4_7), .o(n_3272) );
na02f80 g566678 ( .a(x_in_1_7), .b(x_in_0_7), .o(n_3258) );
in01f80 g566679 ( .a(n_2156), .o(n_2157) );
no02f80 g566680 ( .a(x_in_1_6), .b(x_in_0_6), .o(n_2156) );
na02f80 g566681 ( .a(x_in_9_3), .b(x_in_9_6), .o(n_5221) );
no02f80 g566682 ( .a(x_in_1_2), .b(x_in_0_2), .o(n_3256) );
in01f80 g566683 ( .a(n_2154), .o(n_2155) );
no02f80 g566684 ( .a(x_in_1_13), .b(x_in_0_13), .o(n_2154) );
no02f80 g566685 ( .a(x_in_5_6), .b(x_in_4_2), .o(n_2813) );
na02f80 g566686 ( .a(x_in_5_10), .b(x_in_4_6), .o(n_2810) );
in01f80 g566687 ( .a(n_2152), .o(n_2153) );
no02f80 g566688 ( .a(x_in_41_15), .b(x_in_40_14), .o(n_2152) );
na02f80 g566689 ( .a(x_in_1_10), .b(x_in_0_10), .o(n_3268) );
in01f80 g566690 ( .a(n_2265), .o(n_2266) );
na02f80 g566691 ( .a(x_in_1_2), .b(x_in_0_2), .o(n_2265) );
na02f80 g566692 ( .a(n_2230), .b(x_in_9_3), .o(n_5034) );
no02f80 g566693 ( .a(n_2332), .b(x_in_11_0), .o(n_4391) );
in01f80 g566694 ( .a(n_7054), .o(n_4392) );
na02f80 g566695 ( .a(n_2332), .b(x_in_11_0), .o(n_7054) );
na02f80 g566696 ( .a(n_2618), .b(x_in_55_0), .o(n_6504) );
in01f80 g566697 ( .a(n_7076), .o(n_2471) );
na02f80 g566698 ( .a(n_2445), .b(x_in_59_0), .o(n_7076) );
na02f80 g566699 ( .a(n_2646), .b(x_in_23_0), .o(n_7156) );
no02f80 g566700 ( .a(n_2478), .b(x_in_27_0), .o(n_4595) );
no02f80 g566701 ( .a(n_2061), .b(x_in_35_0), .o(n_3864) );
na02f80 g566702 ( .a(n_2616), .b(x_in_47_0), .o(n_7159) );
na02f80 g566703 ( .a(x_in_57_1), .b(x_in_57_0), .o(n_2382) );
no02f80 g566704 ( .a(n_2413), .b(x_in_5_0), .o(n_3354) );
na02f80 g566705 ( .a(n_2707), .b(x_in_13_0), .o(n_7166) );
na02f80 g566706 ( .a(n_2603), .b(x_in_63_0), .o(n_7150) );
in01f80 g566707 ( .a(n_7048), .o(n_4804) );
na02f80 g566708 ( .a(n_2478), .b(x_in_27_0), .o(n_7048) );
na02f80 g566709 ( .a(x_out_38_32), .b(FE_OFN306_n_3069), .o(n_4340) );
in01f80 g566710 ( .a(n_7051), .o(n_4533) );
na02f80 g566711 ( .a(n_2349), .b(x_in_43_0), .o(n_7051) );
in01f80 g566712 ( .a(n_7855), .o(n_4035) );
na02f80 g566713 ( .a(n_2061), .b(x_in_35_0), .o(n_7855) );
na02f80 g566714 ( .a(n_2593), .b(x_in_15_0), .o(n_7162) );
in01f80 g566715 ( .a(n_3292), .o(n_2392) );
na02f80 g566716 ( .a(n_2607), .b(x_in_39_0), .o(n_3292) );
na02f80 g566717 ( .a(n_2660), .b(x_in_31_0), .o(n_7153) );
no02f80 g566718 ( .a(n_2349), .b(x_in_43_0), .o(n_4534) );
na02f80 g566719 ( .a(x_in_9_8), .b(x_in_9_5), .o(n_5219) );
no02f80 g566720 ( .a(x_in_41_1), .b(x_in_41_0), .o(n_2590) );
no02f80 g566721 ( .a(x_in_1_0), .b(x_in_1_1), .o(n_2628) );
na02f80 g566722 ( .a(x_in_36_13), .b(x_in_36_12), .o(n_26962) );
na02f80 g566723 ( .a(x_in_9_9), .b(x_in_9_6), .o(n_5217) );
na02f80 g566724 ( .a(x_in_9_10), .b(x_in_9_7), .o(n_5023) );
na02f80 g566725 ( .a(x_in_9_4), .b(x_in_9_0), .o(n_2003) );
no02f80 g566726 ( .a(x_in_29_12), .b(x_in_29_15), .o(n_5213) );
no02f80 g566727 ( .a(x_in_4_13), .b(x_in_4_12), .o(n_23376) );
na02f80 g566728 ( .a(x_in_49_0), .b(x_in_49_2), .o(n_2030) );
na02f80 g566729 ( .a(x_in_9_4), .b(x_in_9_7), .o(n_5211) );
no02f80 g566730 ( .a(n_2413), .b(n_2539), .o(n_7174) );
na02f80 g566731 ( .a(x_in_57_2), .b(x_in_57_0), .o(n_2029) );
na02f80 g566732 ( .a(x_in_45_0), .b(x_in_45_3), .o(n_7993) );
na02f80 g566733 ( .a(x_in_57_1), .b(x_in_57_2), .o(n_7172) );
na02f80 g566734 ( .a(x_in_11_15), .b(x_in_11_14), .o(n_1979) );
na02f80 g566735 ( .a(x_in_39_3), .b(x_in_39_2), .o(n_9187) );
in01f80 g566736 ( .a(n_3215), .o(n_4076) );
na02f80 g566737 ( .a(n_2537), .b(n_2037), .o(n_3215) );
na02f80 g566738 ( .a(x_in_9_11), .b(x_in_9_8), .o(n_5209) );
in01f80 g566739 ( .a(n_5813), .o(n_6584) );
no02f80 g566740 ( .a(x_in_11_12), .b(x_in_11_15), .o(n_5813) );
no02f80 g566741 ( .a(x_in_39_13), .b(x_in_39_14), .o(n_2625) );
na02f80 g566742 ( .a(x_in_7_2), .b(x_in_7_0), .o(n_7144) );
in01f80 g566743 ( .a(n_2599), .o(n_2247) );
na02f80 g566744 ( .a(x_in_29_11), .b(x_in_29_13), .o(n_2599) );
in01f80 g566745 ( .a(n_4948), .o(n_9295) );
na02f80 g566746 ( .a(x_in_9_14), .b(x_in_9_11), .o(n_4948) );
no02f80 g566747 ( .a(x_in_51_1), .b(x_in_51_0), .o(n_1995) );
in01f80 g566748 ( .a(n_5105), .o(n_2256) );
na02f80 g566749 ( .a(x_in_51_1), .b(x_in_51_0), .o(n_5105) );
in01f80 g566750 ( .a(n_12425), .o(n_2243) );
na02f80 g566751 ( .a(x_in_45_14), .b(x_in_45_11), .o(n_12425) );
na02f80 g566752 ( .a(x_in_45_13), .b(x_in_45_10), .o(n_3100) );
no02f80 g566753 ( .a(x_in_57_3), .b(x_in_57_1), .o(n_1994) );
na02f80 g566754 ( .a(x_in_9_13), .b(x_in_9_10), .o(n_4768) );
no02f80 g566755 ( .a(x_in_29_14), .b(x_in_29_13), .o(n_2002) );
na02f80 g566756 ( .a(x_in_3_0), .b(x_in_3_1), .o(n_4766) );
in01f80 g566757 ( .a(n_3485), .o(n_2151) );
na02f80 g566758 ( .a(x_in_41_13), .b(x_in_41_14), .o(n_3485) );
na02f80 g566759 ( .a(x_in_11_1), .b(x_in_11_2), .o(n_7597) );
in01f80 g566760 ( .a(n_3758), .o(n_5863) );
na02f80 g566761 ( .a(x_in_9_4), .b(x_in_9_1), .o(n_3758) );
na02f80 g566762 ( .a(x_in_43_1), .b(x_in_43_2), .o(n_7594) );
na02f80 g566763 ( .a(x_in_51_2), .b(x_in_51_0), .o(n_6038) );
no02f80 g566764 ( .a(x_in_15_14), .b(x_in_15_13), .o(n_3872) );
no02f80 g566765 ( .a(x_in_47_14), .b(x_in_47_13), .o(n_3870) );
no02f80 g566766 ( .a(x_in_13_13), .b(x_in_13_14), .o(n_2835) );
no02f80 g566767 ( .a(x_in_63_14), .b(x_in_63_13), .o(n_3504) );
in01f80 g566768 ( .a(n_4099), .o(n_4231) );
na02f80 g566769 ( .a(x_in_13_11), .b(x_in_13_13), .o(n_4099) );
na02f80 g566770 ( .a(x_in_9_12), .b(x_in_9_9), .o(n_5207) );
no02f80 g566771 ( .a(x_in_3_12), .b(x_in_3_15), .o(n_5204) );
na02f80 g566772 ( .a(x_in_13_2), .b(x_in_13_1), .o(n_2320) );
in01f80 g566773 ( .a(n_2350), .o(n_2239) );
na02f80 g566774 ( .a(x_in_11_3), .b(x_in_11_1), .o(n_2350) );
in01f80 g566775 ( .a(n_4345), .o(n_3273) );
na02f80 g566776 ( .a(x_in_45_10), .b(x_in_45_7), .o(n_4345) );
in01f80 g566777 ( .a(n_3178), .o(n_2259) );
na02f80 g566778 ( .a(x_in_43_3), .b(x_in_43_1), .o(n_3178) );
in01f80 g566779 ( .a(n_4059), .o(n_4482) );
na02f80 g566780 ( .a(x_in_45_11), .b(x_in_45_8), .o(n_4059) );
no02f80 g566781 ( .a(x_in_49_4), .b(x_in_49_2), .o(n_7924) );
na02f80 g566782 ( .a(n_2452), .b(n_2636), .o(n_2150) );
in01f80 g566783 ( .a(n_5446), .o(n_2238) );
na02f80 g566784 ( .a(x_in_41_3), .b(x_in_41_2), .o(n_5446) );
na02f80 g566785 ( .a(x_in_27_2), .b(x_in_27_1), .o(n_7591) );
in01f80 g566786 ( .a(n_5723), .o(n_5835) );
no02f80 g566787 ( .a(x_in_49_15), .b(x_in_49_12), .o(n_5723) );
in01f80 g566788 ( .a(n_5810), .o(n_6458) );
no02f80 g566789 ( .a(x_in_27_12), .b(x_in_27_15), .o(n_5810) );
in01f80 g566790 ( .a(n_5807), .o(n_6508) );
no02f80 g566791 ( .a(x_in_43_15), .b(x_in_43_12), .o(n_5807) );
in01f80 g566792 ( .a(n_2209), .o(n_2210) );
no02f80 g566793 ( .a(x_in_5_15), .b(x_in_4_13), .o(n_2209) );
na02f80 g566794 ( .a(x_in_25_3), .b(x_in_25_1), .o(n_4144) );
no02f80 g566795 ( .a(x_in_13_4), .b(x_in_13_2), .o(n_4759) );
in01f80 g566796 ( .a(n_2565), .o(n_4065) );
na02f80 g566797 ( .a(x_in_55_5), .b(x_in_55_1), .o(n_2565) );
in01f80 g566798 ( .a(n_3761), .o(n_3762) );
na02f80 g566799 ( .a(x_in_23_5), .b(x_in_23_1), .o(n_3761) );
in01f80 g566800 ( .a(n_2571), .o(n_3764) );
na02f80 g566801 ( .a(x_in_63_5), .b(x_in_63_1), .o(n_2571) );
in01f80 g566802 ( .a(n_2686), .o(n_3749) );
na02f80 g566803 ( .a(x_in_15_5), .b(x_in_15_1), .o(n_2686) );
no02f80 g566804 ( .a(x_in_23_13), .b(x_in_23_14), .o(n_2401) );
in01f80 g566805 ( .a(n_2267), .o(n_2268) );
no02f80 g566806 ( .a(x_in_21_13), .b(x_in_21_15), .o(n_2267) );
no02f80 g566807 ( .a(x_in_55_13), .b(x_in_55_14), .o(n_2532) );
na02f80 g566808 ( .a(x_in_21_1), .b(x_in_21_0), .o(n_4763) );
in01f80 g566809 ( .a(n_7919), .o(n_2148) );
na02f80 g566810 ( .a(x_in_59_2), .b(x_in_59_1), .o(n_7919) );
no02f80 g566811 ( .a(x_in_31_13), .b(x_in_31_14), .o(n_2596) );
in01f80 g566812 ( .a(n_2110), .o(n_2111) );
no02f80 g566813 ( .a(x_in_51_12), .b(x_in_51_15), .o(n_2110) );
no02f80 g566814 ( .a(x_in_29_3), .b(x_in_29_1), .o(n_4250) );
in01f80 g566815 ( .a(n_4800), .o(n_4984) );
no02f80 g566816 ( .a(x_in_33_13), .b(x_in_33_14), .o(n_4800) );
na02f80 g566817 ( .a(x_in_33_14), .b(x_in_33_13), .o(n_3185) );
in01f80 g566818 ( .a(n_4431), .o(n_4433) );
na02f80 g566819 ( .a(x_in_45_6), .b(x_in_45_3), .o(n_4431) );
in01f80 g566820 ( .a(n_4115), .o(n_4596) );
na02f80 g566821 ( .a(x_in_47_11), .b(x_in_47_14), .o(n_4115) );
in01f80 g566822 ( .a(n_3818), .o(n_2147) );
na02f80 g566823 ( .a(x_in_47_5), .b(x_in_47_1), .o(n_3818) );
in01f80 g566824 ( .a(n_4105), .o(n_4415) );
na02f80 g566825 ( .a(x_in_63_11), .b(x_in_63_14), .o(n_4105) );
in01f80 g566826 ( .a(n_4102), .o(n_4405) );
na02f80 g566827 ( .a(x_in_15_11), .b(x_in_15_14), .o(n_4102) );
in01f80 g566828 ( .a(n_3491), .o(n_2205) );
na02f80 g566829 ( .a(x_in_31_5), .b(x_in_31_1), .o(n_3491) );
no02f80 g566830 ( .a(x_in_19_12), .b(x_in_19_15), .o(n_4757) );
na02f80 g566831 ( .a(x_in_19_15), .b(x_in_19_12), .o(n_1988) );
in01f80 g566832 ( .a(n_4317), .o(n_5337) );
no02f80 g566833 ( .a(x_in_33_3), .b(x_in_33_1), .o(n_4317) );
in01f80 g566834 ( .a(n_5319), .o(n_5321) );
na02f80 g566835 ( .a(x_in_33_3), .b(x_in_33_2), .o(n_5319) );
na02f80 g566836 ( .a(x_in_33_2), .b(x_in_33_1), .o(n_2851) );
in01f80 g566837 ( .a(n_2630), .o(n_5416) );
na02f80 g566838 ( .a(x_in_49_3), .b(x_in_49_2), .o(n_2630) );
na02f80 g566839 ( .a(n_23944), .b(n_2112), .o(n_23345) );
in01f80 g566840 ( .a(n_2096), .o(n_2097) );
na02f80 g566841 ( .a(x_in_5_15), .b(x_in_4_12), .o(n_2096) );
in01f80 g566842 ( .a(n_2223), .o(n_2224) );
na02f80 g566843 ( .a(x_in_13_2), .b(x_in_13_3), .o(n_2223) );
in01f80 g566844 ( .a(n_7057), .o(n_2146) );
na02f80 g566845 ( .a(x_in_19_2), .b(x_in_19_1), .o(n_7057) );
no02f80 g566846 ( .a(n_2419), .b(n_3241), .o(n_2817) );
in01f80 g566847 ( .a(n_3752), .o(n_3751) );
na02f80 g566848 ( .a(x_in_41_12), .b(x_in_41_13), .o(n_3752) );
no02f80 g566849 ( .a(x_in_35_12), .b(x_in_35_15), .o(n_5199) );
in01f80 g566850 ( .a(n_3511), .o(n_4475) );
na02f80 g566851 ( .a(x_in_13_4), .b(x_in_13_6), .o(n_3511) );
in01f80 g566852 ( .a(n_9171), .o(n_2290) );
na02f80 g566853 ( .a(x_in_29_3), .b(x_in_29_2), .o(n_9171) );
in01f80 g566854 ( .a(n_2845), .o(n_4453) );
na02f80 g566855 ( .a(x_in_13_9), .b(x_in_13_11), .o(n_2845) );
in01f80 g566856 ( .a(n_4445), .o(n_4447) );
na02f80 g566857 ( .a(x_in_45_9), .b(x_in_45_6), .o(n_4445) );
in01f80 g566858 ( .a(n_3507), .o(n_4416) );
na02f80 g566859 ( .a(x_in_55_11), .b(x_in_55_14), .o(n_3507) );
in01f80 g566860 ( .a(n_3694), .o(n_4518) );
na02f80 g566861 ( .a(x_in_31_11), .b(x_in_31_14), .o(n_3694) );
in01f80 g566862 ( .a(n_3697), .o(n_4424) );
na02f80 g566863 ( .a(x_in_23_11), .b(x_in_23_14), .o(n_3697) );
in01f80 g566864 ( .a(n_3175), .o(n_2068) );
na02f80 g566865 ( .a(x_in_19_3), .b(x_in_19_1), .o(n_3175) );
in01f80 g566866 ( .a(n_3146), .o(n_5342) );
na02f80 g566867 ( .a(n_5252), .b(n_3763), .o(n_3146) );
no02f80 g566868 ( .a(x_in_49_3), .b(x_in_49_1), .o(n_4013) );
in01f80 g566869 ( .a(n_4420), .o(n_4422) );
na02f80 g566870 ( .a(x_in_45_12), .b(x_in_45_9), .o(n_4420) );
in01f80 g566871 ( .a(n_2570), .o(n_5605) );
na02f80 g566872 ( .a(x_in_57_13), .b(x_in_57_14), .o(n_2570) );
na02f80 g566873 ( .a(x_in_25_4), .b(x_in_25_2), .o(n_5700) );
in01f80 g566874 ( .a(n_2144), .o(n_2145) );
no02f80 g566875 ( .a(x_in_25_2), .b(x_in_25_4), .o(n_2144) );
na02f80 g566876 ( .a(x_in_25_3), .b(x_in_25_2), .o(n_7141) );
in01f80 g566877 ( .a(n_4479), .o(n_2040) );
na02f80 g566878 ( .a(x_in_13_5), .b(x_in_13_7), .o(n_4479) );
in01f80 g566879 ( .a(n_3692), .o(n_4480) );
na02f80 g566880 ( .a(x_in_13_7), .b(x_in_13_9), .o(n_3692) );
in01f80 g566881 ( .a(n_4166), .o(n_4165) );
na02f80 g566882 ( .a(x_in_13_6), .b(x_in_13_8), .o(n_4166) );
na02f80 g566883 ( .a(x_in_27_1), .b(x_in_27_3), .o(n_2017) );
na02f80 g566884 ( .a(x_in_49_13), .b(x_in_49_14), .o(n_3170) );
no02f80 g566885 ( .a(x_in_49_13), .b(x_in_49_14), .o(n_4601) );
in01f80 g566886 ( .a(n_5558), .o(n_3917) );
na02f80 g566887 ( .a(x_in_53_1), .b(x_in_53_0), .o(n_5558) );
na02f80 g566888 ( .a(x_in_61_0), .b(x_in_61_1), .o(n_2028) );
in01f80 g566889 ( .a(n_5267), .o(n_2277) );
na02f80 g566890 ( .a(x_in_57_3), .b(x_in_57_2), .o(n_5267) );
in01f80 g566891 ( .a(n_2051), .o(n_2765) );
na02f80 g566892 ( .a(x_in_59_3), .b(x_in_59_1), .o(n_2051) );
na02f80 g566893 ( .a(x_in_33_12), .b(x_in_33_15), .o(n_3143) );
in01f80 g566894 ( .a(n_2042), .o(n_2043) );
no02f80 g566895 ( .a(x_in_33_15), .b(x_in_33_12), .o(n_2042) );
in01f80 g566896 ( .a(n_2044), .o(n_2045) );
no02f80 g566897 ( .a(x_in_17_1), .b(x_in_17_3), .o(n_2044) );
na02f80 g566898 ( .a(x_in_17_3), .b(x_in_17_1), .o(n_2746) );
in01f80 g566899 ( .a(n_9975), .o(n_2046) );
na02f80 g566900 ( .a(x_in_49_4), .b(x_in_49_3), .o(n_9975) );
na02f80 g566901 ( .a(x_in_37_1), .b(x_in_37_0), .o(n_4863) );
no02f80 g566902 ( .a(x_in_37_1), .b(x_in_37_0), .o(n_1981) );
in01f80 g566903 ( .a(n_7138), .o(n_2276) );
no02f80 g566904 ( .a(x_in_13_10), .b(x_in_13_14), .o(n_7138) );
na02f80 g566905 ( .a(x_in_61_2), .b(x_in_61_0), .o(n_6693) );
in01f80 g566906 ( .a(n_5195), .o(n_5747) );
na02f80 g566907 ( .a(x_in_7_3), .b(x_in_7_2), .o(n_5195) );
in01f80 g566908 ( .a(n_2364), .o(n_2260) );
no02f80 g566909 ( .a(x_in_7_3), .b(x_in_7_2), .o(n_2364) );
in01f80 g566910 ( .a(n_4473), .o(n_3686) );
na02f80 g566911 ( .a(x_in_13_5), .b(x_in_13_3), .o(n_4473) );
in01f80 g566912 ( .a(n_4093), .o(n_4520) );
na02f80 g566913 ( .a(x_in_23_6), .b(x_in_23_3), .o(n_4093) );
in01f80 g566914 ( .a(n_4460), .o(n_4462) );
na02f80 g566915 ( .a(x_in_63_6), .b(x_in_63_3), .o(n_4460) );
na02f80 g566916 ( .a(n_5430), .b(n_3075), .o(n_3076) );
na02f80 g566917 ( .a(n_4946), .b(n_2780), .o(n_2781) );
na02f80 g566918 ( .a(x_in_41_4), .b(x_in_41_3), .o(n_4822) );
in01f80 g566919 ( .a(n_4566), .o(n_4583) );
na02f80 g566920 ( .a(x_in_47_6), .b(x_in_47_3), .o(n_4566) );
in01f80 g566921 ( .a(n_4257), .o(n_4259) );
na02f80 g566922 ( .a(x_in_31_6), .b(x_in_31_3), .o(n_4257) );
na02f80 g566923 ( .a(n_5336), .b(n_3079), .o(n_3131) );
na02f80 g566924 ( .a(n_5365), .b(n_2747), .o(n_2753) );
in01f80 g566925 ( .a(n_4457), .o(n_2207) );
na02f80 g566926 ( .a(x_in_15_6), .b(x_in_15_3), .o(n_4457) );
na02f80 g566927 ( .a(n_5351), .b(n_2828), .o(n_3289) );
na02f80 g566928 ( .a(n_5373), .b(n_2721), .o(n_3293) );
in01f80 g566929 ( .a(n_4449), .o(n_4451) );
na02f80 g566930 ( .a(x_in_55_6), .b(x_in_55_3), .o(n_4449) );
in01f80 g566931 ( .a(n_5805), .o(n_7212) );
no02f80 g566932 ( .a(x_in_59_12), .b(x_in_59_15), .o(n_5805) );
no02f80 g566933 ( .a(x_in_11_12), .b(x_in_11_10), .o(n_1978) );
in01f80 g566934 ( .a(n_2705), .o(n_4456) );
na02f80 g566935 ( .a(x_in_13_8), .b(x_in_13_10), .o(n_2705) );
in01f80 g566936 ( .a(n_4185), .o(n_4090) );
na02f80 g566937 ( .a(x_in_45_8), .b(x_in_45_5), .o(n_4185) );
in01f80 g566938 ( .a(n_4435), .o(n_4437) );
na02f80 g566939 ( .a(x_in_45_7), .b(x_in_45_4), .o(n_4435) );
na02f80 g566940 ( .a(n_2060), .b(x_in_9_5), .o(n_4980) );
no02f80 g566941 ( .a(n_5025), .b(x_in_11_15), .o(n_4030) );
in01f80 g566942 ( .a(n_2318), .o(n_2319) );
no02f80 g566943 ( .a(n_1480), .b(x_in_9_0), .o(n_2318) );
in01f80 g566944 ( .a(n_3342), .o(n_2142) );
na02f80 g566945 ( .a(x_in_37_13), .b(x_in_37_14), .o(n_3342) );
in01f80 g566946 ( .a(n_6945), .o(n_2598) );
na02f80 g566947 ( .a(n_2385), .b(x_in_45_0), .o(n_6945) );
no02f80 g566948 ( .a(x_in_3_2), .b(x_in_3_1), .o(n_1980) );
na02f80 g566949 ( .a(x_in_3_2), .b(x_in_3_1), .o(n_7134) );
no02f80 g566950 ( .a(x_in_37_13), .b(x_in_37_14), .o(n_3242) );
na02f80 g566951 ( .a(n_7317), .b(x_in_39_12), .o(n_3208) );
no02f80 g566952 ( .a(n_2222), .b(x_in_57_0), .o(n_3617) );
in01f80 g566953 ( .a(n_2321), .o(n_4972) );
na02f80 g566954 ( .a(n_2036), .b(x_in_39_11), .o(n_2321) );
na02f80 g566955 ( .a(n_2607), .b(x_in_39_2), .o(n_3291) );
in01f80 g566956 ( .a(n_3024), .o(n_7653) );
no02f80 g566957 ( .a(n_5216), .b(x_in_9_5), .o(n_3024) );
in01f80 g566958 ( .a(n_2362), .o(n_3424) );
no02f80 g566959 ( .a(n_2442), .b(x_in_45_0), .o(n_2362) );
na02f80 g566960 ( .a(n_2409), .b(x_in_29_0), .o(n_3516) );
in01f80 g566961 ( .a(n_2594), .o(n_2595) );
na02f80 g566962 ( .a(n_5025), .b(x_in_11_15), .o(n_2594) );
na02f80 g566963 ( .a(n_2699), .b(x_in_7_0), .o(n_2700) );
no02f80 g566964 ( .a(x_in_7_12), .b(x_in_7_15), .o(n_5961) );
in01f80 g566965 ( .a(n_5902), .o(n_3809) );
no02f80 g566966 ( .a(x_in_33_5), .b(x_in_33_3), .o(n_5902) );
in01f80 g566967 ( .a(n_5929), .o(n_2141) );
no02f80 g566968 ( .a(x_in_61_12), .b(x_in_61_15), .o(n_5929) );
in01f80 g566969 ( .a(n_4401), .o(n_3659) );
no02f80 g566970 ( .a(n_2329), .b(n_11297), .o(n_4401) );
in01f80 g566971 ( .a(n_6325), .o(n_2716) );
no02f80 g566972 ( .a(x_in_57_15), .b(x_in_57_14), .o(n_6325) );
in01f80 g566973 ( .a(n_3138), .o(n_5339) );
no02f80 g566974 ( .a(x_in_13_11), .b(x_in_13_12), .o(n_3138) );
na02f80 g566975 ( .a(x_in_51_1), .b(x_in_51_2), .o(n_7907) );
na02f80 g566976 ( .a(x_in_57_15), .b(x_in_57_14), .o(n_2715) );
na02f80 g566977 ( .a(x_in_21_2), .b(x_in_21_0), .o(n_4870) );
na02f80 g566978 ( .a(x_in_53_2), .b(x_in_53_1), .o(n_2672) );
no02f80 g566979 ( .a(x_in_17_2), .b(x_in_17_1), .o(n_1977) );
no02f80 g566980 ( .a(x_in_25_14), .b(x_in_25_15), .o(n_2768) );
in01f80 g566981 ( .a(n_7840), .o(n_7842) );
no02f80 g566982 ( .a(x_in_51_3), .b(x_in_51_1), .o(n_7840) );
no02f80 g566983 ( .a(n_5180), .b(n_4932), .o(n_4742) );
na02f80 g566984 ( .a(x_in_37_2), .b(x_in_37_0), .o(n_3151) );
in01f80 g566985 ( .a(n_2633), .o(n_3757) );
na02f80 g566986 ( .a(x_in_41_5), .b(x_in_41_3), .o(n_2633) );
in01f80 g566987 ( .a(n_9336), .o(n_3723) );
na02f80 g566988 ( .a(x_in_17_1), .b(x_in_17_2), .o(n_9336) );
in01f80 g566989 ( .a(n_4846), .o(n_2103) );
na02f80 g566990 ( .a(x_in_25_14), .b(x_in_25_15), .o(n_4846) );
in01f80 g566991 ( .a(n_5407), .o(n_2423) );
no02f80 g566992 ( .a(n_7915), .b(n_11409), .o(n_5407) );
na02f80 g566993 ( .a(x_in_7_7), .b(x_in_7_6), .o(n_4740) );
in01f80 g566994 ( .a(n_2584), .o(n_5395) );
na02f80 g566995 ( .a(x_in_41_7), .b(x_in_41_6), .o(n_2584) );
na02f80 g566996 ( .a(x_in_41_9), .b(x_in_41_10), .o(n_2617) );
na02f80 g566997 ( .a(n_2540), .b(n_2517), .o(n_2104) );
in01f80 g566998 ( .a(n_2555), .o(n_6724) );
na02f80 g566999 ( .a(x_in_21_10), .b(x_in_21_13), .o(n_2555) );
na02f80 g567000 ( .a(x_in_41_8), .b(x_in_41_7), .o(n_2610) );
in01f80 g567001 ( .a(n_2106), .o(n_2107) );
na02f80 g567002 ( .a(x_in_45_5), .b(x_in_45_1), .o(n_2106) );
no02f80 g567003 ( .a(x_in_11_9), .b(x_in_11_7), .o(n_2008) );
in01f80 g567004 ( .a(n_2641), .o(n_4955) );
na02f80 g567005 ( .a(x_in_41_9), .b(x_in_41_8), .o(n_2641) );
na02f80 g567006 ( .a(n_5352), .b(n_3229), .o(n_2274) );
in01f80 g567007 ( .a(n_3364), .o(n_2769) );
na02f80 g567008 ( .a(x_in_25_13), .b(x_in_25_14), .o(n_3364) );
in01f80 g567009 ( .a(n_6472), .o(n_6473) );
na02f80 g567010 ( .a(x_in_21_11), .b(x_in_21_14), .o(n_6472) );
no02f80 g567011 ( .a(x_in_7_5), .b(x_in_7_3), .o(n_2723) );
in01f80 g567012 ( .a(n_3755), .o(n_3156) );
no02f80 g567013 ( .a(x_in_53_4), .b(x_in_53_2), .o(n_3755) );
na02f80 g567014 ( .a(x_in_7_5), .b(x_in_7_3), .o(n_2724) );
na02f80 g567015 ( .a(x_in_53_4), .b(x_in_53_2), .o(n_3124) );
na02f80 g567016 ( .a(x_in_35_2), .b(x_in_35_1), .o(n_8837) );
no02f80 g567017 ( .a(x_in_61_13), .b(x_in_61_12), .o(n_2010) );
in01f80 g567018 ( .a(n_7554), .o(n_3832) );
na02f80 g567019 ( .a(x_in_61_13), .b(x_in_61_12), .o(n_7554) );
in01f80 g567020 ( .a(n_6769), .o(n_4579) );
na02f80 g567021 ( .a(x_in_61_14), .b(x_in_61_13), .o(n_6769) );
na02f80 g567022 ( .a(x_in_57_13), .b(x_in_57_12), .o(n_5192) );
no02f80 g567023 ( .a(x_in_61_13), .b(x_in_61_14), .o(n_3195) );
in01f80 g567024 ( .a(n_5838), .o(n_8539) );
no02f80 g567025 ( .a(x_in_33_4), .b(x_in_33_2), .o(n_5838) );
in01f80 g567026 ( .a(n_4471), .o(n_2759) );
na02f80 g567027 ( .a(x_in_63_10), .b(x_in_63_13), .o(n_4471) );
in01f80 g567028 ( .a(n_4531), .o(n_3294) );
na02f80 g567029 ( .a(x_in_47_10), .b(x_in_47_13), .o(n_4531) );
na02f80 g567030 ( .a(x_in_33_4), .b(x_in_33_3), .o(n_2573) );
in01f80 g567031 ( .a(n_4369), .o(n_4129) );
na02f80 g567032 ( .a(x_in_15_10), .b(x_in_15_13), .o(n_4369) );
in01f80 g567033 ( .a(n_4732), .o(n_5592) );
na02f80 g567034 ( .a(x_in_7_7), .b(x_in_7_8), .o(n_4732) );
in01f80 g567035 ( .a(n_2113), .o(n_2114) );
no02f80 g567036 ( .a(x_in_5_14), .b(x_in_5_13), .o(n_2113) );
in01f80 g567037 ( .a(n_4570), .o(n_4798) );
na02f80 g567038 ( .a(x_in_23_4), .b(x_in_23_7), .o(n_4570) );
in01f80 g567039 ( .a(n_4506), .o(n_2838) );
na02f80 g567040 ( .a(x_in_15_4), .b(x_in_15_7), .o(n_4506) );
in01f80 g567041 ( .a(n_4441), .o(n_3135) );
na02f80 g567042 ( .a(x_in_31_4), .b(x_in_31_7), .o(n_4441) );
in01f80 g567043 ( .a(n_6784), .o(n_4734) );
na02f80 g567044 ( .a(x_in_7_13), .b(x_in_7_14), .o(n_6784) );
in01f80 g567045 ( .a(n_4464), .o(n_3284) );
na02f80 g567046 ( .a(x_in_63_4), .b(x_in_63_7), .o(n_4464) );
in01f80 g567047 ( .a(n_4487), .o(n_3281) );
na02f80 g567048 ( .a(x_in_47_4), .b(x_in_47_7), .o(n_4487) );
na02f80 g567049 ( .a(n_2430), .b(n_5089), .o(n_2244) );
in01f80 g567050 ( .a(n_4503), .o(n_3140) );
na02f80 g567051 ( .a(x_in_55_7), .b(x_in_55_4), .o(n_4503) );
na02f80 g567052 ( .a(x_in_5_14), .b(x_in_5_13), .o(n_4151) );
in01f80 g567053 ( .a(n_3868), .o(n_2280) );
na02f80 g567054 ( .a(x_in_41_6), .b(x_in_41_5), .o(n_3868) );
in01f80 g567055 ( .a(n_4970), .o(n_6478) );
no02f80 g567056 ( .a(n_4992), .b(n_2635), .o(n_4970) );
in01f80 g567057 ( .a(n_4911), .o(n_6386) );
na02f80 g567058 ( .a(x_in_7_6), .b(x_in_7_5), .o(n_4911) );
na02f80 g567059 ( .a(n_5390), .b(n_5156), .o(n_2795) );
in01f80 g567060 ( .a(n_2794), .o(n_3777) );
na02f80 g567061 ( .a(x_in_35_3), .b(x_in_35_1), .o(n_2794) );
in01f80 g567062 ( .a(n_3853), .o(n_4890) );
na02f80 g567063 ( .a(x_in_13_10), .b(x_in_13_12), .o(n_3853) );
na02f80 g567064 ( .a(x_in_39_14), .b(FE_OFN347_n_4860), .o(n_7424) );
in01f80 g567065 ( .a(n_4511), .o(n_4512) );
na02f80 g567066 ( .a(x_in_55_9), .b(x_in_55_12), .o(n_4511) );
in01f80 g567067 ( .a(n_4466), .o(n_3338) );
na02f80 g567068 ( .a(x_in_63_6), .b(x_in_63_9), .o(n_4466) );
na02f80 g567069 ( .a(n_2139), .b(x_in_3_2), .o(n_4725) );
no02f80 g567070 ( .a(n_2440), .b(x_in_19_0), .o(n_5074) );
in01f80 g567071 ( .a(n_4408), .o(n_2055) );
na02f80 g567072 ( .a(x_in_55_5), .b(x_in_55_8), .o(n_4408) );
in01f80 g567073 ( .a(n_3669), .o(n_4145) );
na02f80 g567074 ( .a(x_in_23_9), .b(x_in_23_12), .o(n_3669) );
na02f80 g567075 ( .a(n_2285), .b(x_in_9_7), .o(n_5130) );
in01f80 g567076 ( .a(n_7757), .o(n_2542) );
na02f80 g567077 ( .a(n_2490), .b(x_in_51_0), .o(n_7757) );
in01f80 g567078 ( .a(n_4413), .o(n_3119) );
na02f80 g567079 ( .a(x_in_23_6), .b(x_in_23_9), .o(n_4413) );
in01f80 g567080 ( .a(n_2245), .o(n_4516) );
na02f80 g567081 ( .a(x_in_15_6), .b(x_in_15_9), .o(n_2245) );
na02f80 g567082 ( .a(n_2589), .b(n_3188), .o(n_2218) );
na02f80 g567083 ( .a(n_2289), .b(x_in_9_4), .o(n_4645) );
in01f80 g567084 ( .a(n_4500), .o(n_3327) );
na02f80 g567085 ( .a(x_in_55_6), .b(x_in_55_9), .o(n_4500) );
in01f80 g567086 ( .a(n_7815), .o(n_2393) );
na02f80 g567087 ( .a(n_2272), .b(x_in_3_0), .o(n_7815) );
na02f80 g567088 ( .a(n_2588), .b(n_5095), .o(n_2216) );
in01f80 g567089 ( .a(n_4522), .o(n_3122) );
na02f80 g567090 ( .a(x_in_63_9), .b(x_in_63_12), .o(n_4522) );
in01f80 g567091 ( .a(n_4883), .o(n_2815) );
na02f80 g567092 ( .a(x_in_31_9), .b(x_in_31_12), .o(n_4883) );
na02f80 g567093 ( .a(n_2488), .b(x_in_9_8), .o(n_4894) );
no02f80 g567094 ( .a(n_5247), .b(x_in_3_15), .o(n_3848) );
in01f80 g567095 ( .a(n_3104), .o(n_7754) );
no02f80 g567096 ( .a(n_2039), .b(x_in_19_2), .o(n_3104) );
in01f80 g567097 ( .a(n_4486), .o(n_2217) );
na02f80 g567098 ( .a(x_in_15_5), .b(x_in_15_8), .o(n_4486) );
in01f80 g567099 ( .a(n_4497), .o(n_2693) );
na02f80 g567100 ( .a(x_in_47_9), .b(x_in_47_12), .o(n_4497) );
na02f80 g567101 ( .a(n_2588), .b(n_2589), .o(n_2225) );
na02f80 g567102 ( .a(n_6726), .b(x_in_9_10), .o(n_3387) );
in01f80 g567103 ( .a(n_4439), .o(n_3420) );
na02f80 g567104 ( .a(x_in_31_6), .b(x_in_31_9), .o(n_4439) );
na02f80 g567105 ( .a(n_2354), .b(x_in_13_12), .o(n_4835) );
in01f80 g567106 ( .a(n_8191), .o(n_2219) );
na02f80 g567107 ( .a(x_in_57_4), .b(x_in_57_3), .o(n_8191) );
na02f80 g567108 ( .a(n_2248), .b(x_in_9_6), .o(n_4608) );
in01f80 g567109 ( .a(n_4426), .o(n_4427) );
na02f80 g567110 ( .a(x_in_15_9), .b(x_in_15_12), .o(n_4426) );
na02f80 g567111 ( .a(n_8957), .b(x_in_9_9), .o(n_5161) );
na02f80 g567112 ( .a(n_610), .b(x_in_51_2), .o(n_2246) );
in01f80 g567113 ( .a(n_3431), .o(n_4217) );
na02f80 g567114 ( .a(x_in_63_5), .b(x_in_63_8), .o(n_3431) );
in01f80 g567115 ( .a(n_4491), .o(n_4493) );
na02f80 g567116 ( .a(x_in_23_5), .b(x_in_23_8), .o(n_4491) );
no02f80 g567117 ( .a(n_4687), .b(x_in_17_0), .o(n_5048) );
in01f80 g567118 ( .a(n_4411), .o(n_3672) );
na02f80 g567119 ( .a(x_in_47_6), .b(x_in_47_9), .o(n_4411) );
in01f80 g567120 ( .a(n_2649), .o(n_2650) );
na02f80 g567121 ( .a(n_5247), .b(x_in_3_15), .o(n_2649) );
no02f80 g567122 ( .a(x_in_57_4), .b(x_in_57_3), .o(n_2007) );
in01f80 g567123 ( .a(n_2330), .o(n_2226) );
na02f80 g567124 ( .a(x_in_59_2), .b(x_in_59_3), .o(n_2330) );
na02f80 g567125 ( .a(n_3186), .b(n_2737), .o(n_2249) );
na02f80 g567126 ( .a(n_5825), .b(n_4419), .o(n_2215) );
in01f80 g567127 ( .a(n_3234), .o(n_3417) );
na02f80 g567128 ( .a(x_in_3_3), .b(x_in_3_1), .o(n_3234) );
in01f80 g567129 ( .a(n_2287), .o(n_2288) );
na02f80 g567130 ( .a(x_in_35_2), .b(x_in_35_5), .o(n_2287) );
na02f80 g567131 ( .a(x_in_51_14), .b(x_in_51_11), .o(n_2696) );
in01f80 g567132 ( .a(n_2220), .o(n_2221) );
no02f80 g567133 ( .a(x_in_51_11), .b(x_in_51_14), .o(n_2220) );
no02f80 g567134 ( .a(x_in_19_5), .b(x_in_19_3), .o(n_4325) );
na02f80 g567135 ( .a(n_5310), .b(n_7818), .o(n_2208) );
in01f80 g567136 ( .a(n_6643), .o(n_2629) );
no02f80 g567137 ( .a(n_3887), .b(n_5977), .o(n_6643) );
no02f80 g567138 ( .a(n_5390), .b(n_5369), .o(n_3987) );
no02f80 g567139 ( .a(x_in_7_7), .b(x_in_7_5), .o(n_2032) );
na02f80 g567140 ( .a(x_in_37_2), .b(x_in_37_1), .o(n_7893) );
in01f80 g567141 ( .a(n_7124), .o(n_2211) );
na02f80 g567142 ( .a(x_in_25_11), .b(x_in_25_14), .o(n_7124) );
in01f80 g567143 ( .a(n_2275), .o(n_4374) );
na02f80 g567144 ( .a(x_in_15_8), .b(x_in_15_11), .o(n_2275) );
in01f80 g567145 ( .a(n_3662), .o(n_4209) );
na02f80 g567146 ( .a(x_in_31_5), .b(x_in_31_8), .o(n_3662) );
na02f80 g567147 ( .a(x_in_37_6), .b(x_in_37_4), .o(n_3202) );
in01f80 g567148 ( .a(n_4198), .o(n_3450) );
na02f80 g567149 ( .a(x_in_63_8), .b(x_in_63_11), .o(n_4198) );
in01f80 g567150 ( .a(n_4495), .o(n_4134) );
na02f80 g567151 ( .a(x_in_47_8), .b(x_in_47_11), .o(n_4495) );
in01f80 g567152 ( .a(n_4443), .o(n_3372) );
na02f80 g567153 ( .a(x_in_23_8), .b(x_in_23_11), .o(n_4443) );
in01f80 g567154 ( .a(n_4429), .o(n_3665) );
na02f80 g567155 ( .a(x_in_55_8), .b(x_in_55_11), .o(n_4429) );
in01f80 g567156 ( .a(n_4458), .o(n_3467) );
na02f80 g567157 ( .a(x_in_31_8), .b(x_in_31_11), .o(n_4458) );
in01f80 g567158 ( .a(n_3459), .o(n_4489) );
na02f80 g567159 ( .a(x_in_47_5), .b(x_in_47_8), .o(n_3459) );
no02f80 g567160 ( .a(x_in_37_4), .b(x_in_37_6), .o(n_3201) );
na02f80 g567161 ( .a(x_in_35_14), .b(x_in_35_11), .o(n_2676) );
in01f80 g567162 ( .a(n_6984), .o(n_4657) );
na02f80 g567163 ( .a(x_in_53_3), .b(x_in_53_2), .o(n_6984) );
no02f80 g567164 ( .a(n_5272), .b(n_8522), .o(n_3351) );
na02f80 g567165 ( .a(x_in_41_12), .b(x_in_41_11), .o(n_2614) );
in01f80 g567166 ( .a(n_4309), .o(n_3300) );
na02f80 g567167 ( .a(x_in_23_10), .b(x_in_23_13), .o(n_4309) );
in01f80 g567168 ( .a(n_4508), .o(n_3306) );
na02f80 g567169 ( .a(x_in_55_10), .b(x_in_55_13), .o(n_4508) );
in01f80 g567170 ( .a(n_4484), .o(n_3114) );
na02f80 g567171 ( .a(x_in_31_10), .b(x_in_31_13), .o(n_4484) );
no02f80 g567172 ( .a(n_3036), .b(n_5869), .o(n_7481) );
in01f80 g567173 ( .a(n_6667), .o(n_7454) );
no02f80 g567174 ( .a(x_in_37_4), .b(x_in_37_2), .o(n_6667) );
no02f80 g567175 ( .a(n_2240), .b(n_3011), .o(n_2241) );
no02f80 g567176 ( .a(x_in_5_4), .b(x_in_5_5), .o(n_2453) );
in01f80 g567177 ( .a(n_6355), .o(n_4843) );
na02f80 g567178 ( .a(x_in_7_8), .b(x_in_7_9), .o(n_6355) );
no02f80 g567179 ( .a(x_in_61_3), .b(x_in_61_1), .o(n_7835) );
na02f80 g567180 ( .a(x_in_57_6), .b(x_in_57_5), .o(n_4722) );
in01f80 g567181 ( .a(n_3753), .o(n_3841) );
no02f80 g567182 ( .a(x_in_19_10), .b(x_in_19_8), .o(n_3753) );
in01f80 g567183 ( .a(n_3849), .o(n_2678) );
na02f80 g567184 ( .a(n_5940), .b(n_5537), .o(n_3849) );
in01f80 g567185 ( .a(n_3263), .o(n_8340) );
na02f80 g567186 ( .a(x_in_59_8), .b(x_in_59_7), .o(n_3263) );
no02f80 g567187 ( .a(n_5691), .b(n_2363), .o(n_6409) );
na02f80 g567188 ( .a(x_in_57_7), .b(x_in_57_8), .o(n_4155) );
na02f80 g567189 ( .a(x_in_57_8), .b(x_in_57_9), .o(n_4720) );
in01f80 g567190 ( .a(n_3780), .o(n_3729) );
no02f80 g567191 ( .a(x_in_19_8), .b(x_in_19_6), .o(n_3780) );
na02f80 g567192 ( .a(x_in_57_7), .b(x_in_57_6), .o(n_4719) );
in01f80 g567193 ( .a(n_2283), .o(n_2855) );
na02f80 g567194 ( .a(x_in_33_13), .b(x_in_33_11), .o(n_2283) );
na02f80 g567195 ( .a(n_9646), .b(n_2520), .o(n_2115) );
in01f80 g567196 ( .a(n_2837), .o(n_4068) );
na02f80 g567197 ( .a(x_in_17_5), .b(x_in_17_3), .o(n_2837) );
in01f80 g567198 ( .a(n_5344), .o(n_5346) );
na02f80 g567199 ( .a(n_5939), .b(n_2440), .o(n_5344) );
no02f80 g567200 ( .a(n_3193), .b(n_2762), .o(n_2763) );
in01f80 g567201 ( .a(n_6307), .o(n_7560) );
na02f80 g567202 ( .a(x_in_7_12), .b(x_in_7_13), .o(n_6307) );
na02f80 g567203 ( .a(x_in_37_12), .b(x_in_37_10), .o(n_2733) );
no02f80 g567204 ( .a(x_in_49_11), .b(x_in_49_10), .o(n_2021) );
no02f80 g567205 ( .a(x_in_37_10), .b(x_in_37_12), .o(n_2732) );
in01f80 g567206 ( .a(n_2656), .o(n_2033) );
no02f80 g567207 ( .a(x_in_53_11), .b(x_in_53_15), .o(n_2656) );
na02f80 g567208 ( .a(x_in_57_9), .b(x_in_57_10), .o(n_4716) );
no02f80 g567209 ( .a(n_5699), .b(n_5275), .o(n_7790) );
na02f80 g567210 ( .a(x_in_37_9), .b(x_in_37_7), .o(n_3204) );
na02f80 g567211 ( .a(x_in_37_7), .b(x_in_37_5), .o(n_3197) );
na02f80 g567212 ( .a(x_in_59_10), .b(x_in_59_9), .o(n_6405) );
in01f80 g567213 ( .a(n_5866), .o(n_5868) );
na02f80 g567214 ( .a(x_in_61_3), .b(x_in_61_2), .o(n_5866) );
in01f80 g567215 ( .a(n_5431), .o(n_4196) );
na02f80 g567216 ( .a(x_in_61_6), .b(x_in_61_5), .o(n_5431) );
na02f80 g567217 ( .a(n_3174), .b(n_5940), .o(n_4664) );
in01f80 g567218 ( .a(n_2088), .o(n_2089) );
na02f80 g567219 ( .a(x_in_35_10), .b(x_in_35_7), .o(n_2088) );
no02f80 g567220 ( .a(x_in_37_7), .b(x_in_37_9), .o(n_3203) );
in01f80 g567221 ( .a(n_4163), .o(n_8564) );
na02f80 g567222 ( .a(x_in_51_3), .b(x_in_51_2), .o(n_4163) );
no02f80 g567223 ( .a(x_in_37_5), .b(x_in_37_7), .o(n_3196) );
no02f80 g567224 ( .a(x_in_7_4), .b(x_in_7_2), .o(n_2000) );
na02f80 g567225 ( .a(x_in_21_1), .b(x_in_21_2), .o(n_7887) );
in01f80 g567226 ( .a(n_3756), .o(n_3157) );
na02f80 g567227 ( .a(x_in_53_5), .b(x_in_53_1), .o(n_3756) );
na02f80 g567228 ( .a(x_in_37_12), .b(x_in_37_11), .o(n_2772) );
no02f80 g567229 ( .a(x_in_37_12), .b(x_in_37_11), .o(n_2771) );
no02f80 g567230 ( .a(x_in_37_3), .b(x_in_37_1), .o(n_2023) );
no02f80 g567231 ( .a(n_4654), .b(n_4376), .o(n_2138) );
na02f80 g567232 ( .a(FE_OFN1110_rst), .b(x_in_43_15), .o(n_8188) );
na02f80 g567233 ( .a(x_in_39_2), .b(n_27194), .o(n_7330) );
in01f80 g567234 ( .a(FE_OFN282_n_7349), .o(n_2773) );
na02f80 g567235 ( .a(x_in_27_15), .b(FE_OFN331_n_4860), .o(n_7349) );
no02f80 g567236 ( .a(x_in_37_8), .b(x_in_37_6), .o(n_2713) );
in01f80 g567237 ( .a(n_6387), .o(n_3447) );
na02f80 g567238 ( .a(x_in_61_7), .b(x_in_61_6), .o(n_6387) );
na02f80 g567239 ( .a(x_in_37_8), .b(x_in_37_6), .o(n_2714) );
na02f80 g567240 ( .a(x_in_35_10), .b(x_in_35_13), .o(n_3978) );
no02f80 g567241 ( .a(x_in_61_7), .b(x_in_61_6), .o(n_1985) );
no02f80 g567242 ( .a(x_in_43_12), .b(x_in_43_10), .o(n_1998) );
no02f80 g567243 ( .a(x_in_27_12), .b(x_in_27_10), .o(n_1986) );
na02f80 g567244 ( .a(n_3736), .b(x_in_29_13), .o(n_3773) );
no02f80 g567245 ( .a(n_5369), .b(n_5098), .o(n_3558) );
no02f80 g567246 ( .a(n_2643), .b(x_in_9_14), .o(n_2991) );
no02f80 g567247 ( .a(x_in_61_3), .b(x_in_61_5), .o(n_3207) );
na02f80 g567248 ( .a(n_6420), .b(x_in_51_15), .o(n_3811) );
no02f80 g567249 ( .a(x_in_3_12), .b(x_in_3_10), .o(n_1991) );
na02f80 g567250 ( .a(x_in_53_8), .b(x_in_53_9), .o(n_3530) );
no02f80 g567251 ( .a(x_in_3_9), .b(x_in_3_7), .o(n_1982) );
in01f80 g567252 ( .a(n_3346), .o(n_2344) );
no02f80 g567253 ( .a(n_2537), .b(x_in_39_2), .o(n_3346) );
na02f80 g567254 ( .a(n_5515), .b(n_5524), .o(n_2048) );
in01f80 g567255 ( .a(n_2390), .o(n_2391) );
na02f80 g567256 ( .a(n_2875), .b(x_in_29_13), .o(n_2390) );
no02f80 g567257 ( .a(n_7263), .b(x_in_43_15), .o(n_3839) );
na02f80 g567258 ( .a(x_in_53_7), .b(x_in_53_8), .o(n_3535) );
na02f80 g567259 ( .a(n_2376), .b(x_in_9_13), .o(n_4205) );
in01f80 g567260 ( .a(n_2338), .o(n_2339) );
na02f80 g567261 ( .a(n_7263), .b(x_in_43_15), .o(n_2338) );
in01f80 g567262 ( .a(n_2057), .o(n_2058) );
na02f80 g567263 ( .a(x_in_61_5), .b(x_in_61_3), .o(n_2057) );
na02f80 g567264 ( .a(x_in_21_6), .b(x_in_21_9), .o(n_6641) );
na02f80 g567265 ( .a(x_in_53_7), .b(x_in_53_6), .o(n_3399) );
in01f80 g567266 ( .a(n_2708), .o(n_2322) );
no02f80 g567267 ( .a(n_3107), .b(x_in_39_3), .o(n_2708) );
na02f80 g567268 ( .a(n_5524), .b(n_5666), .o(n_2047) );
no02f80 g567269 ( .a(n_5244), .b(x_in_19_15), .o(n_3063) );
in01f80 g567270 ( .a(n_3845), .o(n_5046) );
no02f80 g567271 ( .a(n_2875), .b(x_in_29_12), .o(n_3845) );
in01f80 g567272 ( .a(n_7781), .o(n_2090) );
na02f80 g567273 ( .a(x_in_59_6), .b(x_in_59_5), .o(n_7781) );
in01f80 g567274 ( .a(n_3847), .o(n_2342) );
no02f80 g567275 ( .a(n_6420), .b(x_in_51_15), .o(n_3847) );
no02f80 g567276 ( .a(n_7402), .b(x_in_27_15), .o(n_4080) );
in01f80 g567277 ( .a(n_2324), .o(n_2325) );
na02f80 g567278 ( .a(n_7402), .b(x_in_27_15), .o(n_2324) );
in01f80 g567279 ( .a(n_4000), .o(n_2507) );
no02f80 g567280 ( .a(n_8537), .b(x_in_29_12), .o(n_4000) );
na02f80 g567281 ( .a(n_5987), .b(n_2061), .o(n_2062) );
no02f80 g567282 ( .a(n_8206), .b(n_11696), .o(n_2076) );
no02f80 g567283 ( .a(n_7323), .b(n_11041), .o(n_2053) );
no02f80 g567284 ( .a(n_7278), .b(n_11040), .o(n_2252) );
in01f80 g567285 ( .a(n_4239), .o(n_4502) );
na02f80 g567286 ( .a(x_in_15_7), .b(x_in_15_10), .o(n_4239) );
in01f80 g567287 ( .a(n_2562), .o(n_2050) );
no02f80 g567288 ( .a(x_in_27_4), .b(x_in_27_3), .o(n_2562) );
in01f80 g567289 ( .a(n_4110), .o(n_4425) );
na02f80 g567290 ( .a(x_in_31_7), .b(x_in_31_10), .o(n_4110) );
no02f80 g567291 ( .a(n_7247), .b(n_11034), .o(n_2136) );
in01f80 g567292 ( .a(n_4388), .o(n_3110) );
na02f80 g567293 ( .a(x_in_23_7), .b(x_in_23_10), .o(n_4388) );
in01f80 g567294 ( .a(n_4547), .o(n_2866) );
na02f80 g567295 ( .a(x_in_47_7), .b(x_in_47_10), .o(n_4547) );
no02f80 g567296 ( .a(n_7338), .b(n_11037), .o(n_2293) );
no02f80 g567297 ( .a(n_6753), .b(n_11698), .o(n_2291) );
in01f80 g567298 ( .a(n_4223), .o(n_2886) );
na02f80 g567299 ( .a(x_in_55_7), .b(x_in_55_10), .o(n_4223) );
in01f80 g567300 ( .a(n_4468), .o(n_2881) );
na02f80 g567301 ( .a(x_in_63_7), .b(x_in_63_10), .o(n_4468) );
in01f80 g567302 ( .a(n_2099), .o(n_2789) );
na02f80 g567303 ( .a(x_in_21_3), .b(x_in_21_1), .o(n_2099) );
in01f80 g567304 ( .a(n_2254), .o(n_2255) );
no02f80 g567305 ( .a(x_in_21_1), .b(x_in_21_3), .o(n_2254) );
na02f80 g567306 ( .a(x_in_57_12), .b(x_in_57_11), .o(n_5308) );
no02f80 g567307 ( .a(x_in_3_7), .b(x_in_3_5), .o(n_1999) );
no02f80 g567308 ( .a(n_7320), .b(n_8165), .o(n_7551) );
no02f80 g567309 ( .a(x_in_59_5), .b(x_in_59_3), .o(n_3261) );
in01f80 g567310 ( .a(n_2072), .o(n_2073) );
na02f80 g567311 ( .a(x_in_35_12), .b(x_in_35_9), .o(n_2072) );
na02f80 g567312 ( .a(x_in_25_5), .b(x_in_25_4), .o(n_4707) );
in01f80 g567313 ( .a(n_2556), .o(n_2080) );
na02f80 g567314 ( .a(x_in_25_5), .b(x_in_25_3), .o(n_2556) );
na02f80 g567315 ( .a(x_in_35_8), .b(x_in_35_5), .o(n_3971) );
no02f80 g567316 ( .a(x_in_43_9), .b(x_in_43_7), .o(n_2019) );
no02f80 g567317 ( .a(x_in_27_8), .b(x_in_27_6), .o(n_1976) );
in01f80 g567318 ( .a(n_2086), .o(n_2087) );
na02f80 g567319 ( .a(x_in_17_14), .b(x_in_17_11), .o(n_2086) );
no02f80 g567320 ( .a(x_in_37_4), .b(x_in_37_3), .o(n_2026) );
in01f80 g567321 ( .a(n_5716), .o(n_3127) );
na02f80 g567322 ( .a(x_in_37_4), .b(x_in_37_3), .o(n_5716) );
no02f80 g567323 ( .a(x_in_19_12), .b(x_in_19_10), .o(n_5938) );
in01f80 g567324 ( .a(n_4022), .o(n_2064) );
na02f80 g567325 ( .a(x_in_17_6), .b(x_in_17_3), .o(n_4022) );
no02f80 g567326 ( .a(n_23944), .b(n_3169), .o(n_2832) );
in01f80 g567327 ( .a(n_7480), .o(n_5185) );
na02f80 g567328 ( .a(x_in_21_8), .b(x_in_21_5), .o(n_7480) );
in01f80 g567329 ( .a(n_7541), .o(n_4967) );
na02f80 g567330 ( .a(x_in_21_8), .b(x_in_21_11), .o(n_7541) );
no02f80 g567331 ( .a(x_in_37_11), .b(x_in_37_9), .o(n_2031) );
in01f80 g567332 ( .a(n_2372), .o(n_2273) );
na02f80 g567333 ( .a(x_in_53_5), .b(x_in_53_4), .o(n_2372) );
in01f80 g567334 ( .a(n_2098), .o(n_6363) );
na02f80 g567335 ( .a(x_in_21_7), .b(x_in_21_4), .o(n_2098) );
na02f80 g567336 ( .a(x_in_57_10), .b(x_in_57_11), .o(n_4352) );
na02f80 g567337 ( .a(x_in_53_5), .b(x_in_53_6), .o(n_3968) );
na02f80 g567338 ( .a(x_in_37_10), .b(x_in_37_8), .o(n_2720) );
no02f80 g567339 ( .a(x_in_3_5), .b(x_in_3_3), .o(n_1987) );
no02f80 g567340 ( .a(x_in_37_8), .b(x_in_37_10), .o(n_2719) );
no02f80 g567341 ( .a(x_in_27_10), .b(x_in_27_8), .o(n_2018) );
no02f80 g567342 ( .a(x_in_43_10), .b(x_in_43_8), .o(n_1990) );
no02f80 g567343 ( .a(x_in_43_8), .b(x_in_43_6), .o(n_1989) );
no02f80 g567344 ( .a(x_in_27_9), .b(x_in_27_7), .o(n_2024) );
in01f80 g567345 ( .a(n_3415), .o(n_3838) );
no02f80 g567346 ( .a(x_in_19_6), .b(x_in_19_4), .o(n_3415) );
in01f80 g567347 ( .a(n_6767), .o(n_4651) );
na02f80 g567348 ( .a(x_in_61_12), .b(x_in_61_11), .o(n_6767) );
in01f80 g567349 ( .a(n_5820), .o(n_2135) );
no02f80 g567350 ( .a(x_in_33_7), .b(x_in_33_5), .o(n_5820) );
no02f80 g567351 ( .a(x_in_61_12), .b(x_in_61_11), .o(n_2027) );
na02f80 g567352 ( .a(x_in_33_7), .b(x_in_33_5), .o(n_2798) );
in01f80 g567353 ( .a(n_3177), .o(n_2092) );
no02f80 g567354 ( .a(x_in_43_4), .b(x_in_43_5), .o(n_3177) );
na02f80 g567355 ( .a(x_in_53_9), .b(x_in_53_10), .o(n_3545) );
na02f80 g567356 ( .a(x_in_53_12), .b(x_in_53_11), .o(n_4138) );
na02f80 g567357 ( .a(x_in_7_11), .b(x_in_7_12), .o(n_6653) );
in01f80 g567358 ( .a(n_6748), .o(n_4355) );
na02f80 g567359 ( .a(x_in_7_10), .b(x_in_7_11), .o(n_6748) );
no02f80 g567360 ( .a(x_in_27_7), .b(x_in_27_5), .o(n_1996) );
in01f80 g567361 ( .a(n_2741), .o(n_2547) );
na02f80 g567362 ( .a(n_4654), .b(n_5742), .o(n_2741) );
na02f80 g567363 ( .a(n_5931), .b(n_5515), .o(n_2094) );
na02f80 g567364 ( .a(x_in_37_5), .b(x_in_37_3), .o(n_4573) );
no02f80 g567365 ( .a(x_in_19_5), .b(x_in_19_4), .o(n_2009) );
in01f80 g567366 ( .a(n_5730), .o(n_4976) );
na02f80 g567367 ( .a(x_in_37_3), .b(x_in_37_2), .o(n_5730) );
na02f80 g567368 ( .a(x_in_63_15), .b(n_27012), .o(n_8198) );
na02f80 g567369 ( .a(x_in_15_15), .b(n_27012), .o(n_8056) );
na02f80 g567370 ( .a(x_in_47_15), .b(n_27012), .o(n_7406) );
na02f80 g567371 ( .a(x_in_31_15), .b(n_27012), .o(n_7575) );
na02f80 g567372 ( .a(x_in_55_15), .b(FE_OFN146_n_2667), .o(n_7361) );
na02f80 g567373 ( .a(x_in_23_15), .b(FE_OFN146_n_2667), .o(n_8204) );
in01f80 g567374 ( .a(n_5596), .o(n_6731) );
na02f80 g567375 ( .a(x_in_61_8), .b(x_in_61_7), .o(n_5596) );
na02f80 g567376 ( .a(x_in_53_10), .b(x_in_53_11), .o(n_3963) );
no02f80 g567377 ( .a(x_in_61_8), .b(x_in_61_7), .o(n_2012) );
in01f80 g567378 ( .a(n_8756), .o(n_2119) );
no02f80 g567379 ( .a(x_in_53_10), .b(x_in_53_14), .o(n_8756) );
na02f80 g567380 ( .a(n_8206), .b(x_in_63_15), .o(n_2212) );
na02f80 g567381 ( .a(n_8032), .b(x_in_41_13), .o(n_3796) );
na02f80 g567382 ( .a(n_7247), .b(x_in_47_15), .o(n_2133) );
in01f80 g567383 ( .a(n_4461), .o(n_4463) );
no02f80 g567384 ( .a(n_5351), .b(x_in_63_1), .o(n_4461) );
no02f80 g567385 ( .a(n_2528), .b(x_in_45_10), .o(n_4659) );
na02f80 g567386 ( .a(n_5032), .b(x_in_35_15), .o(n_3902) );
no02f80 g567387 ( .a(n_2134), .b(x_in_45_13), .o(n_4604) );
in01f80 g567388 ( .a(n_2504), .o(n_10829) );
na02f80 g567389 ( .a(n_2214), .b(x_in_41_12), .o(n_2504) );
no02f80 g567390 ( .a(n_7216), .b(x_in_45_10), .o(n_2065) );
in01f80 g567391 ( .a(n_3903), .o(n_2612) );
no02f80 g567392 ( .a(n_5032), .b(x_in_35_15), .o(n_3903) );
in01f80 g567393 ( .a(n_6952), .o(n_2587) );
no02f80 g567394 ( .a(n_2517), .b(x_in_5_2), .o(n_6952) );
na02f80 g567395 ( .a(n_7338), .b(x_in_15_15), .o(n_2100) );
in01f80 g567396 ( .a(n_2373), .o(n_4574) );
na02f80 g567397 ( .a(n_2538), .b(x_in_33_12), .o(n_2373) );
na02f80 g567398 ( .a(n_7323), .b(x_in_23_15), .o(n_2059) );
no02f80 g567399 ( .a(n_2527), .b(x_in_45_11), .o(n_4958) );
na02f80 g567400 ( .a(n_3077), .b(x_in_13_13), .o(n_3827) );
in01f80 g567401 ( .a(n_4258), .o(n_4260) );
no02f80 g567402 ( .a(n_5373), .b(x_in_31_1), .o(n_4258) );
in01f80 g567403 ( .a(n_4582), .o(n_4567) );
no02f80 g567404 ( .a(n_5365), .b(x_in_47_1), .o(n_4582) );
na02f80 g567405 ( .a(n_7278), .b(x_in_55_15), .o(n_2281) );
in01f80 g567406 ( .a(n_3287), .o(n_2444) );
no02f80 g567407 ( .a(n_4946), .b(x_in_15_1), .o(n_3287) );
in01f80 g567408 ( .a(n_3859), .o(n_2389) );
no02f80 g567409 ( .a(n_7216), .b(x_in_45_14), .o(n_3859) );
na02f80 g567410 ( .a(n_2049), .b(x_in_45_12), .o(n_3324) );
in01f80 g567411 ( .a(n_2658), .o(n_2659) );
na02f80 g567412 ( .a(n_10486), .b(x_in_45_11), .o(n_2658) );
in01f80 g567413 ( .a(n_4450), .o(n_4452) );
no02f80 g567414 ( .a(n_5336), .b(x_in_55_1), .o(n_4450) );
na02f80 g567415 ( .a(n_6753), .b(x_in_31_15), .o(n_2063) );
in01f80 g567416 ( .a(n_2503), .o(n_5401) );
na02f80 g567417 ( .a(n_2214), .b(x_in_41_14), .o(n_2503) );
na02f80 g567418 ( .a(n_2214), .b(x_in_41_15), .o(n_2213) );
in01f80 g567419 ( .a(n_4521), .o(n_4094) );
no02f80 g567420 ( .a(n_5430), .b(x_in_23_1), .o(n_4521) );
na02f80 g567421 ( .a(x_in_19_11), .b(x_in_19_13), .o(n_4698) );
in01f80 g567422 ( .a(n_2198), .o(n_2949) );
na02f80 g567423 ( .a(x_in_53_4), .b(x_in_53_3), .o(n_2198) );
in01f80 g567424 ( .a(n_3323), .o(n_6955) );
no02f80 g567425 ( .a(n_2668), .b(n_8482), .o(n_3323) );
na02f80 g567426 ( .a(x_in_59_12), .b(x_in_59_11), .o(n_8336) );
in01f80 g567427 ( .a(n_2263), .o(n_2264) );
na02f80 g567428 ( .a(x_in_35_11), .b(x_in_35_8), .o(n_2263) );
in01f80 g567429 ( .a(n_7088), .o(n_2132) );
na02f80 g567430 ( .a(x_in_25_7), .b(x_in_25_4), .o(n_7088) );
na02f80 g567431 ( .a(x_in_51_4), .b(x_in_51_2), .o(n_2939) );
no02f80 g567432 ( .a(x_in_51_4), .b(x_in_51_2), .o(n_2938) );
na02f80 g567433 ( .a(x_in_25_6), .b(x_in_25_5), .o(n_4004) );
no02f80 g567434 ( .a(x_in_27_11), .b(x_in_27_9), .o(n_2006) );
no02f80 g567435 ( .a(x_in_43_11), .b(x_in_43_9), .o(n_1993) );
na02f80 g567436 ( .a(n_5931), .b(n_5963), .o(n_2233) );
no02f80 g567437 ( .a(x_in_27_5), .b(x_in_27_4), .o(n_2004) );
no02f80 g567438 ( .a(x_in_3_11), .b(x_in_3_9), .o(n_2015) );
no02f80 g567439 ( .a(x_in_61_2), .b(x_in_61_4), .o(n_3209) );
na02f80 g567440 ( .a(x_in_61_4), .b(x_in_61_2), .o(n_3210) );
in01f80 g567441 ( .a(n_7082), .o(n_2054) );
na02f80 g567442 ( .a(x_in_25_8), .b(x_in_25_5), .o(n_7082) );
no02f80 g567443 ( .a(x_in_51_10), .b(x_in_51_12), .o(n_3262) );
in01f80 g567444 ( .a(n_3781), .o(n_2511) );
na02f80 g567445 ( .a(n_5537), .b(n_7765), .o(n_3781) );
no02f80 g567446 ( .a(x_in_59_6), .b(x_in_59_4), .o(n_2016) );
na02f80 g567447 ( .a(x_in_59_6), .b(x_in_59_4), .o(n_2878) );
in01f80 g567448 ( .a(n_4386), .o(n_7776) );
na02f80 g567449 ( .a(x_in_59_5), .b(x_in_59_4), .o(n_4386) );
in01f80 g567450 ( .a(n_2130), .o(n_2131) );
na02f80 g567451 ( .a(x_in_35_7), .b(x_in_35_4), .o(n_2130) );
in01f80 g567452 ( .a(n_7443), .o(n_4923) );
na02f80 g567453 ( .a(x_in_61_9), .b(x_in_61_8), .o(n_7443) );
no02f80 g567454 ( .a(x_in_61_9), .b(x_in_61_8), .o(n_2011) );
na02f80 g567455 ( .a(x_in_53_14), .b(x_in_53_13), .o(n_3052) );
in01f80 g567456 ( .a(n_5153), .o(n_5137) );
no02f80 g567457 ( .a(x_in_53_14), .b(x_in_53_13), .o(n_5153) );
in01f80 g567458 ( .a(n_2122), .o(n_3309) );
na02f80 g567459 ( .a(x_in_61_4), .b(x_in_61_3), .o(n_2122) );
in01f80 g567460 ( .a(n_5571), .o(n_6716) );
na02f80 g567461 ( .a(x_in_21_6), .b(x_in_21_3), .o(n_5571) );
in01f80 g567462 ( .a(n_7079), .o(n_2129) );
na02f80 g567463 ( .a(x_in_25_13), .b(x_in_25_10), .o(n_7079) );
no02f80 g567464 ( .a(n_7434), .b(n_8557), .o(n_2206) );
in01f80 g567465 ( .a(n_7445), .o(n_3576) );
no02f80 g567466 ( .a(n_4914), .b(n_3833), .o(n_7445) );
in01f80 g567467 ( .a(n_4203), .o(n_3015) );
no02f80 g567468 ( .a(x_in_33_6), .b(x_in_33_4), .o(n_4203) );
no02f80 g567469 ( .a(x_in_61_10), .b(x_in_61_9), .o(n_2020) );
na02f80 g567470 ( .a(x_in_33_6), .b(x_in_33_4), .o(n_2877) );
na02f80 g567471 ( .a(x_in_53_13), .b(x_in_53_12), .o(n_3954) );
in01f80 g567472 ( .a(n_4887), .o(n_4888) );
na02f80 g567473 ( .a(x_in_31_14), .b(FE_OFN1171_n_4860), .o(n_4887) );
in01f80 g567474 ( .a(n_2986), .o(n_2987) );
na02f80 g567475 ( .a(x_in_55_14), .b(n_15183), .o(n_2986) );
in01f80 g567476 ( .a(n_4319), .o(n_4320) );
na02f80 g567477 ( .a(x_in_23_14), .b(FE_OFN1155_n_14586), .o(n_4319) );
no02f80 g567478 ( .a(n_3043), .b(x_in_21_15), .o(n_4063) );
no02f80 g567479 ( .a(n_3746), .b(x_in_21_0), .o(n_2140) );
no02f80 g567480 ( .a(n_5435), .b(x_in_41_3), .o(n_2128) );
in01f80 g567481 ( .a(n_4474), .o(n_3687) );
na02f80 g567482 ( .a(n_2707), .b(x_in_13_2), .o(n_4474) );
in01f80 g567483 ( .a(n_4011), .o(n_2663) );
no02f80 g567484 ( .a(n_2451), .b(x_in_33_0), .o(n_4011) );
in01f80 g567485 ( .a(n_2857), .o(n_2662) );
no02f80 g567486 ( .a(n_2424), .b(x_in_41_2), .o(n_2857) );
na02f80 g567487 ( .a(n_2234), .b(x_in_49_2), .o(n_5126) );
na02f80 g567488 ( .a(n_2535), .b(x_in_25_3), .o(n_2948) );
na02f80 g567489 ( .a(n_3043), .b(x_in_21_15), .o(n_4062) );
no02f80 g567490 ( .a(n_7434), .b(x_in_21_0), .o(n_4148) );
in01f80 g567491 ( .a(n_4027), .o(n_4228) );
no02f80 g567492 ( .a(n_2597), .b(x_in_29_11), .o(n_4027) );
no02f80 g567493 ( .a(n_2066), .b(x_in_21_1), .o(n_2067) );
no02f80 g567494 ( .a(x_in_51_10), .b(x_in_51_8), .o(n_3199) );
in01f80 g567495 ( .a(n_5228), .o(n_3106) );
no02f80 g567496 ( .a(x_in_33_8), .b(x_in_33_10), .o(n_5228) );
na02f80 g567497 ( .a(x_in_51_10), .b(x_in_51_8), .o(n_2682) );
na02f80 g567498 ( .a(x_in_51_8), .b(x_in_51_6), .o(n_2669) );
in01f80 g567499 ( .a(n_3776), .o(n_2084) );
na02f80 g567500 ( .a(x_in_17_7), .b(x_in_17_10), .o(n_3776) );
in01f80 g567501 ( .a(n_6723), .o(n_4397) );
na02f80 g567502 ( .a(x_in_61_11), .b(x_in_61_10), .o(n_6723) );
na02f80 g567503 ( .a(x_in_33_8), .b(x_in_33_6), .o(n_3072) );
na02f80 g567504 ( .a(x_in_33_9), .b(x_in_33_7), .o(n_3070) );
no02f80 g567505 ( .a(x_in_51_8), .b(x_in_51_6), .o(n_2695) );
in01f80 g567506 ( .a(n_5231), .o(n_3073) );
no02f80 g567507 ( .a(x_in_33_9), .b(x_in_33_7), .o(n_5231) );
no02f80 g567508 ( .a(x_in_61_11), .b(x_in_61_10), .o(n_2005) );
na02f80 g567509 ( .a(x_in_33_10), .b(x_in_33_8), .o(n_2879) );
in01f80 g567510 ( .a(n_4692), .o(n_5230) );
no02f80 g567511 ( .a(x_in_33_6), .b(x_in_33_8), .o(n_4692) );
in01f80 g567512 ( .a(n_3393), .o(n_2035) );
na02f80 g567513 ( .a(x_in_17_5), .b(x_in_17_8), .o(n_3393) );
na02f80 g567514 ( .a(x_in_25_13), .b(x_in_25_12), .o(n_3949) );
na02f80 g567515 ( .a(x_in_17_12), .b(x_in_17_9), .o(n_3734) );
in01f80 g567516 ( .a(n_5226), .o(n_3173) );
no02f80 g567517 ( .a(x_in_33_10), .b(x_in_33_12), .o(n_5226) );
na02f80 g567518 ( .a(x_in_25_7), .b(x_in_25_6), .o(n_3946) );
in01f80 g567519 ( .a(n_2077), .o(n_2078) );
na02f80 g567520 ( .a(x_in_33_12), .b(x_in_33_10), .o(n_2077) );
in01f80 g567521 ( .a(n_7073), .o(n_2074) );
na02f80 g567522 ( .a(x_in_25_9), .b(x_in_25_6), .o(n_7073) );
no02f80 g567523 ( .a(x_in_21_4), .b(x_in_21_3), .o(n_1984) );
na02f80 g567524 ( .a(x_in_21_5), .b(x_in_21_3), .o(n_2001) );
na02f80 g567525 ( .a(x_in_33_11), .b(x_in_33_9), .o(n_2805) );
in01f80 g567526 ( .a(n_3760), .o(n_2038) );
na02f80 g567527 ( .a(x_in_17_7), .b(x_in_17_4), .o(n_3760) );
in01f80 g567528 ( .a(n_5224), .o(n_3311) );
no02f80 g567529 ( .a(x_in_33_9), .b(x_in_33_11), .o(n_5224) );
no02f80 g567530 ( .a(x_in_51_9), .b(x_in_51_7), .o(n_3314) );
na02f80 g567531 ( .a(x_in_25_10), .b(x_in_25_9), .o(n_3472) );
na02f80 g567532 ( .a(x_in_51_9), .b(x_in_51_7), .o(n_3315) );
na02f80 g567533 ( .a(x_in_25_8), .b(x_in_25_7), .o(n_3464) );
na02f80 g567534 ( .a(x_in_25_9), .b(x_in_25_8), .o(n_3943) );
na02f80 g567535 ( .a(x_in_25_10), .b(x_in_25_7), .o(n_7070) );
no02f80 g567536 ( .a(x_in_51_6), .b(x_in_51_4), .o(n_3212) );
na02f80 g567537 ( .a(x_in_51_6), .b(x_in_51_4), .o(n_2647) );
no02f80 g567538 ( .a(x_in_19_11), .b(x_in_19_12), .o(n_2352) );
na02f80 g567539 ( .a(x_in_59_15), .b(n_4270), .o(n_7239) );
na02f80 g567540 ( .a(x_in_7_15), .b(FE_OFN146_n_2667), .o(n_7261) );
na02f80 g567541 ( .a(x_in_17_9), .b(x_in_17_6), .o(n_3732) );
in01f80 g567542 ( .a(n_7064), .o(n_2127) );
na02f80 g567543 ( .a(x_in_25_9), .b(x_in_25_12), .o(n_7064) );
na02f80 g567544 ( .a(x_in_25_10), .b(x_in_25_11), .o(n_3563) );
in01f80 g567545 ( .a(n_7067), .o(n_2126) );
na02f80 g567546 ( .a(x_in_25_11), .b(x_in_25_8), .o(n_7067) );
in01f80 g567547 ( .a(n_5383), .o(n_2500) );
no02f80 g567548 ( .a(n_7213), .b(x_in_39_11), .o(n_5383) );
no02f80 g567549 ( .a(n_2533), .b(x_in_33_14), .o(n_2856) );
no02f80 g567550 ( .a(n_5689), .b(x_in_51_14), .o(n_3385) );
in01f80 g567551 ( .a(n_3398), .o(n_2600) );
no02f80 g567552 ( .a(n_7340), .b(x_in_7_15), .o(n_3398) );
na02f80 g567553 ( .a(n_2419), .b(x_in_37_15), .o(n_2056) );
no02f80 g567554 ( .a(n_8957), .b(x_in_9_15), .o(n_9207) );
in01f80 g567555 ( .a(n_2499), .o(n_6904) );
no02f80 g567556 ( .a(n_2052), .b(x_in_33_13), .o(n_2499) );
in01f80 g567557 ( .a(n_4213), .o(n_2498) );
na02f80 g567558 ( .a(n_2513), .b(x_in_45_3), .o(n_4213) );
in01f80 g567559 ( .a(n_2496), .o(n_2497) );
na02f80 g567560 ( .a(n_5689), .b(x_in_51_14), .o(n_2496) );
in01f80 g567561 ( .a(n_2998), .o(n_2315) );
na02f80 g567562 ( .a(n_2605), .b(x_in_61_4), .o(n_2998) );
na02f80 g567563 ( .a(n_9118), .b(x_in_49_13), .o(n_4903) );
no02f80 g567564 ( .a(n_2124), .b(x_in_11_13), .o(n_3388) );
in01f80 g567565 ( .a(n_5265), .o(n_4476) );
no02f80 g567566 ( .a(n_2516), .b(x_in_13_2), .o(n_5265) );
na02f80 g567567 ( .a(n_4143), .b(x_in_61_0), .o(n_3310) );
na02f80 g567568 ( .a(n_2691), .b(x_in_49_14), .o(n_2125) );
na02f80 g567569 ( .a(n_2605), .b(x_in_61_2), .o(n_3325) );
in01f80 g567570 ( .a(n_4186), .o(n_4091) );
na02f80 g567571 ( .a(n_2439), .b(x_in_45_4), .o(n_4186) );
in01f80 g567572 ( .a(n_4436), .o(n_4438) );
no02f80 g567573 ( .a(n_2439), .b(x_in_45_2), .o(n_4436) );
in01f80 g567574 ( .a(n_12616), .o(n_2366) );
no02f80 g567575 ( .a(n_2124), .b(x_in_11_11), .o(n_12616) );
na02f80 g567576 ( .a(n_7340), .b(x_in_7_15), .o(n_3397) );
in01f80 g567577 ( .a(n_8517), .o(n_2410) );
na02f80 g567578 ( .a(n_2624), .b(x_in_7_11), .o(n_8517) );
in01f80 g567579 ( .a(n_2368), .o(n_2369) );
na02f80 g567580 ( .a(n_4992), .b(x_in_59_15), .o(n_2368) );
na02f80 g567581 ( .a(n_5252), .b(x_in_19_1), .o(n_2123) );
na02f80 g567582 ( .a(n_4825), .b(x_in_53_0), .o(n_2950) );
in01f80 g567583 ( .a(n_3806), .o(n_3389) );
na02f80 g567584 ( .a(n_2124), .b(x_in_11_13), .o(n_3806) );
no02f80 g567585 ( .a(n_2601), .b(x_in_57_2), .o(n_6938) );
no02f80 g567586 ( .a(n_4992), .b(x_in_59_15), .o(n_3834) );
na02f80 g567587 ( .a(n_2439), .b(x_in_45_6), .o(n_2075) );
in01f80 g567588 ( .a(n_3096), .o(n_2495) );
na02f80 g567589 ( .a(n_2409), .b(x_in_29_2), .o(n_3096) );
in01f80 g567590 ( .a(n_2494), .o(n_12646) );
no02f80 g567591 ( .a(n_2269), .b(x_in_51_11), .o(n_2494) );
na02f80 g567592 ( .a(x_in_17_11), .b(x_in_17_8), .o(n_3731) );
na02f80 g567593 ( .a(x_in_25_11), .b(x_in_25_12), .o(n_3927) );
in01f80 g567594 ( .a(n_3770), .o(n_2091) );
na02f80 g567595 ( .a(x_in_17_10), .b(x_in_17_13), .o(n_3770) );
na02f80 g567596 ( .a(x_in_51_11), .b(x_in_51_9), .o(n_2357) );
no02f80 g567597 ( .a(x_in_51_9), .b(x_in_51_11), .o(n_3198) );
in01f80 g567598 ( .a(n_4194), .o(n_4195) );
na02f80 g567599 ( .a(x_in_47_13), .b(FE_OFN357_n_4860), .o(n_4194) );
in01f80 g567600 ( .a(n_4192), .o(n_4193) );
na02f80 g567601 ( .a(x_in_15_13), .b(FE_OFN355_n_4860), .o(n_4192) );
in01f80 g567602 ( .a(n_4315), .o(n_4316) );
na02f80 g567603 ( .a(x_in_63_13), .b(FE_OFN357_n_4860), .o(n_4315) );
in01f80 g567604 ( .a(n_2808), .o(n_2411) );
na02f80 g567605 ( .a(n_2673), .b(x_in_13_11), .o(n_2808) );
na02f80 g567606 ( .a(n_3126), .b(x_in_37_1), .o(n_2093) );
in01f80 g567607 ( .a(n_4218), .o(n_3432) );
no02f80 g567608 ( .a(n_3737), .b(x_in_63_3), .o(n_4218) );
na02f80 g567609 ( .a(n_2234), .b(x_in_49_3), .o(n_2270) );
na02f80 g567610 ( .a(n_5313), .b(x_in_57_14), .o(n_8701) );
in01f80 g567611 ( .a(n_2493), .o(n_3980) );
no02f80 g567612 ( .a(n_2492), .b(x_in_25_15), .o(n_2493) );
in01f80 g567613 ( .a(n_7760), .o(n_8527) );
na02f80 g567614 ( .a(n_2655), .b(x_in_61_11), .o(n_7760) );
in01f80 g567615 ( .a(n_4951), .o(n_4774) );
no02f80 g567616 ( .a(n_2575), .b(x_in_15_11), .o(n_4951) );
na02f80 g567617 ( .a(n_4376), .b(x_in_37_0), .o(n_2101) );
na02f80 g567618 ( .a(n_3238), .b(x_in_49_4), .o(n_2271) );
in01f80 g567619 ( .a(n_8693), .o(n_2417) );
na02f80 g567620 ( .a(n_5872), .b(x_in_21_14), .o(n_8693) );
in01f80 g567621 ( .a(n_3285), .o(n_4465) );
no02f80 g567622 ( .a(n_2828), .b(x_in_63_2), .o(n_3285) );
in01f80 g567623 ( .a(n_3282), .o(n_4488) );
no02f80 g567624 ( .a(n_2747), .b(x_in_47_2), .o(n_3282) );
in01f80 g567625 ( .a(n_4964), .o(n_4393) );
no02f80 g567626 ( .a(n_2448), .b(x_in_47_11), .o(n_4964) );
in01f80 g567627 ( .a(n_3741), .o(n_2425) );
no02f80 g567628 ( .a(n_3742), .b(x_in_55_3), .o(n_3741) );
na02f80 g567629 ( .a(n_10486), .b(x_in_45_9), .o(n_4997) );
na02f80 g567630 ( .a(n_5180), .b(x_in_51_1), .o(n_2105) );
na02f80 g567631 ( .a(n_3724), .b(x_in_29_2), .o(n_5790) );
in01f80 g567632 ( .a(n_3822), .o(n_2429) );
no02f80 g567633 ( .a(n_2353), .b(x_in_61_15), .o(n_3822) );
in01f80 g567634 ( .a(n_4797), .o(n_4571) );
no02f80 g567635 ( .a(n_3075), .b(x_in_23_2), .o(n_4797) );
na02f80 g567636 ( .a(n_2520), .b(x_in_17_1), .o(n_2121) );
in01f80 g567637 ( .a(n_6032), .o(n_4170) );
na02f80 g567638 ( .a(n_2433), .b(x_in_13_5), .o(n_6032) );
in01f80 g567639 ( .a(n_3044), .o(n_6773) );
na02f80 g567640 ( .a(n_3043), .b(x_in_21_13), .o(n_3044) );
in01f80 g567641 ( .a(n_4490), .o(n_3460) );
no02f80 g567642 ( .a(n_3445), .b(x_in_47_3), .o(n_4490) );
in01f80 g567643 ( .a(n_4636), .o(n_2508) );
na02f80 g567644 ( .a(n_2588), .b(x_in_49_4), .o(n_4636) );
na02f80 g567645 ( .a(n_4794), .b(x_in_17_15), .o(n_5396) );
na02f80 g567646 ( .a(n_3641), .b(x_in_57_14), .o(n_3821) );
no02f80 g567647 ( .a(n_3011), .b(x_in_37_0), .o(n_4639) );
na02f80 g567648 ( .a(n_2353), .b(x_in_61_15), .o(n_3716) );
no02f80 g567649 ( .a(n_2424), .b(x_in_41_4), .o(n_2168) );
in01f80 g567650 ( .a(n_4210), .o(n_3663) );
no02f80 g567651 ( .a(n_3739), .b(x_in_31_3), .o(n_4210) );
in01f80 g567652 ( .a(n_3144), .o(n_3878) );
no02f80 g567653 ( .a(n_2433), .b(x_in_13_3), .o(n_3144) );
in01f80 g567654 ( .a(n_3481), .o(n_2524) );
no02f80 g567655 ( .a(n_3482), .b(x_in_15_3), .o(n_3481) );
na02f80 g567656 ( .a(n_5926), .b(x_in_13_11), .o(n_3025) );
in01f80 g567657 ( .a(n_2839), .o(n_4507) );
no02f80 g567658 ( .a(n_2780), .b(x_in_15_2), .o(n_2839) );
in01f80 g567659 ( .a(n_2751), .o(n_2620) );
na02f80 g567660 ( .a(n_2549), .b(x_in_17_12), .o(n_2751) );
in01f80 g567661 ( .a(n_10793), .o(n_2398) );
no02f80 g567662 ( .a(n_3560), .b(x_in_57_14), .o(n_10793) );
no02f80 g567663 ( .a(n_2428), .b(x_in_45_8), .o(n_3101) );
in01f80 g567664 ( .a(n_5348), .o(n_4779) );
no02f80 g567665 ( .a(n_2523), .b(x_in_63_11), .o(n_5348) );
no02f80 g567666 ( .a(n_2513), .b(x_in_45_9), .o(n_4146) );
in01f80 g567667 ( .a(n_4492), .o(n_4494) );
no02f80 g567668 ( .a(n_3744), .b(x_in_23_3), .o(n_4492) );
in01f80 g567669 ( .a(n_3136), .o(n_4442) );
no02f80 g567670 ( .a(n_2721), .b(x_in_31_2), .o(n_3136) );
in01f80 g567671 ( .a(n_3141), .o(n_4504) );
no02f80 g567672 ( .a(n_3079), .b(x_in_55_2), .o(n_3141) );
in01f80 g567673 ( .a(n_2611), .o(n_21777) );
na02f80 g567674 ( .a(n_2492), .b(x_in_25_15), .o(n_2611) );
no02f80 g567675 ( .a(n_5381), .b(x_in_41_3), .o(n_9095) );
no02f80 g567676 ( .a(n_3641), .b(x_in_57_14), .o(n_3820) );
no02f80 g567677 ( .a(n_3591), .b(x_in_29_2), .o(n_3172) );
in01f80 g567678 ( .a(n_4349), .o(n_4350) );
na02f80 g567679 ( .a(x_in_39_9), .b(FE_OFN1171_n_4860), .o(n_4349) );
in01f80 g567680 ( .a(n_4311), .o(n_4312) );
na02f80 g567681 ( .a(x_in_39_5), .b(FE_OFN336_n_4860), .o(n_4311) );
in01f80 g567682 ( .a(n_2578), .o(n_2579) );
na02f80 g567683 ( .a(n_5272), .b(x_in_7_4), .o(n_2578) );
in01f80 g567684 ( .a(n_3379), .o(n_2415) );
no02f80 g567685 ( .a(n_2752), .b(x_in_35_13), .o(n_3379) );
in01f80 g567686 ( .a(n_2809), .o(n_2685) );
no02f80 g567687 ( .a(n_4514), .b(x_in_39_8), .o(n_2809) );
in01f80 g567688 ( .a(n_4168), .o(n_2491) );
no02f80 g567689 ( .a(n_6500), .b(x_in_39_5), .o(n_4168) );
no02f80 g567690 ( .a(n_5247), .b(x_in_3_14), .o(n_6932) );
in01f80 g567691 ( .a(n_5115), .o(n_3592) );
na02f80 g567692 ( .a(n_3470), .b(x_in_29_3), .o(n_5115) );
in01f80 g567693 ( .a(n_2767), .o(n_2582) );
no02f80 g567694 ( .a(n_7325), .b(x_in_39_6), .o(n_2767) );
in01f80 g567695 ( .a(n_5127), .o(n_2378) );
na02f80 g567696 ( .a(n_2597), .b(x_in_29_10), .o(n_5127) );
in01f80 g567697 ( .a(n_4226), .o(n_2316) );
no02f80 g567698 ( .a(n_3035), .b(x_in_29_9), .o(n_4226) );
in01f80 g567699 ( .a(n_2613), .o(n_4121) );
na02f80 g567700 ( .a(n_2422), .b(x_in_59_13), .o(n_2613) );
in01f80 g567701 ( .a(n_6921), .o(n_6919) );
na02f80 g567702 ( .a(n_2752), .b(x_in_35_12), .o(n_6921) );
in01f80 g567703 ( .a(n_4122), .o(n_4410) );
no02f80 g567704 ( .a(n_2422), .b(x_in_59_13), .o(n_4122) );
in01f80 g567705 ( .a(n_12696), .o(n_12057) );
no02f80 g567706 ( .a(n_2422), .b(x_in_59_11), .o(n_12696) );
na02f80 g567707 ( .a(n_2864), .b(x_in_29_9), .o(n_3056) );
in01f80 g567708 ( .a(n_4929), .o(n_4928) );
na02f80 g567709 ( .a(n_2522), .b(x_in_13_9), .o(n_4929) );
in01f80 g567710 ( .a(n_4421), .o(n_4423) );
no02f80 g567711 ( .a(n_2527), .b(x_in_45_7), .o(n_4421) );
na02f80 g567712 ( .a(n_8522), .b(x_in_7_3), .o(n_3322) );
in01f80 g567713 ( .a(n_3384), .o(n_2602) );
na02f80 g567714 ( .a(n_6746), .b(x_in_3_14), .o(n_3384) );
in01f80 g567715 ( .a(n_5264), .o(n_5263) );
na02f80 g567716 ( .a(n_2506), .b(x_in_13_7), .o(n_5264) );
in01f80 g567717 ( .a(n_4454), .o(n_4455) );
na02f80 g567718 ( .a(n_2657), .b(x_in_13_8), .o(n_4454) );
no02f80 g567719 ( .a(n_2231), .b(x_in_53_3), .o(n_2232) );
in01f80 g567720 ( .a(n_6372), .o(n_4481) );
no02f80 g567721 ( .a(n_2506), .b(x_in_13_5), .o(n_6372) );
in01f80 g567722 ( .a(n_4483), .o(n_4060) );
no02f80 g567723 ( .a(n_2528), .b(x_in_45_6), .o(n_4483) );
in01f80 g567724 ( .a(n_3098), .o(n_2515) );
no02f80 g567725 ( .a(n_4338), .b(x_in_39_4), .o(n_3098) );
in01f80 g567726 ( .a(n_4957), .o(n_4232) );
no02f80 g567727 ( .a(n_2673), .b(x_in_13_9), .o(n_4957) );
in01f80 g567728 ( .a(n_2661), .o(n_3498) );
na02f80 g567729 ( .a(n_2752), .b(x_in_35_13), .o(n_2661) );
in01f80 g567730 ( .a(n_3274), .o(n_4346) );
no02f80 g567731 ( .a(n_2513), .b(x_in_45_5), .o(n_3274) );
in01f80 g567732 ( .a(n_3045), .o(n_4618) );
no02f80 g567733 ( .a(n_2438), .b(x_in_45_8), .o(n_3045) );
no02f80 g567734 ( .a(n_2442), .b(x_in_45_7), .o(n_4220) );
no02f80 g567735 ( .a(n_6746), .b(x_in_3_14), .o(n_4034) );
in01f80 g567736 ( .a(n_7734), .o(n_5695) );
no02f80 g567737 ( .a(n_5827), .b(x_in_53_2), .o(n_7734) );
no02f80 g567738 ( .a(n_3724), .b(x_in_29_3), .o(n_3206) );
in01f80 g567739 ( .a(n_12670), .o(n_2580) );
na02f80 g567740 ( .a(n_8524), .b(x_in_35_14), .o(n_12670) );
in01f80 g567741 ( .a(n_11217), .o(n_12643) );
no02f80 g567742 ( .a(n_2317), .b(x_in_3_11), .o(n_11217) );
in01f80 g567743 ( .a(n_8598), .o(n_4853) );
na02f80 g567744 ( .a(n_4825), .b(x_in_53_2), .o(n_8598) );
in01f80 g567745 ( .a(n_5904), .o(n_2472) );
no02f80 g567746 ( .a(n_8851), .b(x_in_39_9), .o(n_5904) );
na02f80 g567747 ( .a(x_in_7_2), .b(n_27194), .o(n_6737) );
in01f80 g567748 ( .a(n_4881), .o(n_4882) );
na02f80 g567749 ( .a(x_in_27_14), .b(FE_OFN352_n_4860), .o(n_4881) );
in01f80 g567750 ( .a(n_4089), .o(n_4291) );
no02f80 g567751 ( .a(n_3390), .b(x_in_29_8), .o(n_4089) );
in01f80 g567752 ( .a(n_2543), .o(n_2544) );
na02f80 g567753 ( .a(n_3390), .b(x_in_29_7), .o(n_2543) );
no02f80 g567754 ( .a(n_4847), .b(x_in_61_13), .o(n_3298) );
na02f80 g567755 ( .a(n_3724), .b(x_in_29_5), .o(n_2876) );
in01f80 g567756 ( .a(n_2644), .o(n_5789) );
na02f80 g567757 ( .a(n_3390), .b(x_in_29_4), .o(n_2644) );
na02f80 g567758 ( .a(n_9329), .b(x_in_41_10), .o(n_3326) );
na02f80 g567759 ( .a(n_4343), .b(x_in_37_14), .o(n_2143) );
in01f80 g567760 ( .a(n_2486), .o(n_8441) );
no02f80 g567761 ( .a(n_4343), .b(x_in_37_14), .o(n_2486) );
na02f80 g567762 ( .a(n_5900), .b(x_in_21_1), .o(n_2120) );
no02f80 g567763 ( .a(n_5968), .b(x_in_7_5), .o(n_3220) );
no02f80 g567764 ( .a(n_14997), .b(x_in_27_13), .o(n_3501) );
in01f80 g567765 ( .a(n_3233), .o(n_2671) );
na02f80 g567766 ( .a(n_2377), .b(x_in_35_2), .o(n_3233) );
in01f80 g567767 ( .a(n_2563), .o(n_2564) );
na02f80 g567768 ( .a(n_2583), .b(x_in_41_6), .o(n_2563) );
in01f80 g567769 ( .a(n_2559), .o(n_2560) );
na02f80 g567770 ( .a(n_2272), .b(x_in_3_1), .o(n_2559) );
in01f80 g567771 ( .a(n_3725), .o(n_4336) );
no02f80 g567772 ( .a(n_3470), .b(x_in_29_7), .o(n_3725) );
na02f80 g567773 ( .a(n_6781), .b(x_in_21_1), .o(n_2149) );
in01f80 g567774 ( .a(n_2336), .o(n_2337) );
no02f80 g567775 ( .a(n_5256), .b(x_in_7_6), .o(n_2336) );
na02f80 g567776 ( .a(n_3470), .b(x_in_29_6), .o(n_2865) );
no02f80 g567777 ( .a(n_5869), .b(x_in_21_13), .o(n_4616) );
in01f80 g567778 ( .a(n_3879), .o(n_2609) );
no02f80 g567779 ( .a(n_3187), .b(x_in_49_12), .o(n_3879) );
in01f80 g567780 ( .a(n_3027), .o(n_4602) );
na02f80 g567781 ( .a(n_2737), .b(x_in_49_11), .o(n_3027) );
in01f80 g567782 ( .a(n_3885), .o(n_3655) );
no02f80 g567783 ( .a(n_2518), .b(x_in_61_14), .o(n_3885) );
in01f80 g567784 ( .a(n_4920), .o(n_4623) );
no02f80 g567785 ( .a(n_7231), .b(x_in_55_11), .o(n_4920) );
na02f80 g567786 ( .a(n_6494), .b(x_in_7_6), .o(n_3333) );
no02f80 g567787 ( .a(n_5931), .b(x_in_3_2), .o(n_7748) );
na02f80 g567788 ( .a(n_3746), .b(x_in_21_5), .o(n_2041) );
no02f80 g567789 ( .a(n_2377), .b(x_in_35_2), .o(n_3526) );
in01f80 g567790 ( .a(n_3788), .o(n_3500) );
na02f80 g567791 ( .a(n_14997), .b(x_in_27_13), .o(n_3788) );
in01f80 g567792 ( .a(n_5378), .o(n_4626) );
no02f80 g567793 ( .a(n_6488), .b(x_in_23_11), .o(n_5378) );
in01f80 g567794 ( .a(n_3039), .o(n_4323) );
na02f80 g567795 ( .a(n_9610), .b(x_in_41_7), .o(n_3039) );
in01f80 g567796 ( .a(n_4172), .o(n_2443) );
na02f80 g567797 ( .a(n_8537), .b(x_in_29_8), .o(n_4172) );
in01f80 g567798 ( .a(n_12582), .o(n_2400) );
no02f80 g567799 ( .a(n_14997), .b(x_in_27_11), .o(n_12582) );
no02f80 g567800 ( .a(n_5296), .b(x_in_5_3), .o(n_6926) );
in01f80 g567801 ( .a(n_8696), .o(n_2374) );
na02f80 g567802 ( .a(n_4180), .b(x_in_37_14), .o(n_8696) );
in01f80 g567803 ( .a(n_2750), .o(n_2677) );
no02f80 g567804 ( .a(n_8133), .b(x_in_39_7), .o(n_2750) );
no02f80 g567805 ( .a(n_2272), .b(x_in_3_1), .o(n_3629) );
in01f80 g567806 ( .a(n_2484), .o(n_2485) );
na02f80 g567807 ( .a(n_5968), .b(x_in_7_7), .o(n_2484) );
in01f80 g567808 ( .a(n_5354), .o(n_4247) );
no02f80 g567809 ( .a(n_7291), .b(x_in_31_11), .o(n_5354) );
in01f80 g567810 ( .a(n_2387), .o(n_3643) );
na02f80 g567811 ( .a(n_7915), .b(x_in_41_11), .o(n_2387) );
no02f80 g567812 ( .a(n_2864), .b(x_in_29_7), .o(n_3225) );
in01f80 g567813 ( .a(n_4307), .o(n_4308) );
na02f80 g567814 ( .a(x_in_7_14), .b(FE_OFN86_n_14586), .o(n_4307) );
in01f80 g567815 ( .a(n_4515), .o(n_2679) );
no02f80 g567816 ( .a(n_4746), .b(x_in_15_4), .o(n_4515) );
in01f80 g567817 ( .a(n_6895), .o(n_2323) );
no02f80 g567818 ( .a(n_5291), .b(x_in_5_6), .o(n_6895) );
in01f80 g567819 ( .a(n_6875), .o(n_2483) );
na02f80 g567820 ( .a(n_2517), .b(x_in_5_6), .o(n_6875) );
in01f80 g567821 ( .a(n_3082), .o(n_2680) );
no02f80 g567822 ( .a(n_4057), .b(x_in_19_13), .o(n_3082) );
no02f80 g567823 ( .a(n_15590), .b(x_in_7_13), .o(n_2868) );
in01f80 g567824 ( .a(n_3120), .o(n_4414) );
no02f80 g567825 ( .a(n_4744), .b(x_in_23_4), .o(n_3120) );
in01f80 g567826 ( .a(n_2880), .o(n_4672) );
na02f80 g567827 ( .a(n_9608), .b(x_in_41_11), .o(n_2880) );
no02f80 g567828 ( .a(n_7311), .b(x_in_43_13), .o(n_3438) );
no02f80 g567829 ( .a(n_5369), .b(x_in_35_3), .o(n_3782) );
in01f80 g567830 ( .a(n_3650), .o(n_3437) );
na02f80 g567831 ( .a(n_7311), .b(x_in_43_13), .o(n_3650) );
in01f80 g567832 ( .a(n_2481), .o(n_2482) );
no02f80 g567833 ( .a(n_6494), .b(x_in_7_8), .o(n_2481) );
in01f80 g567834 ( .a(n_12599), .o(n_2480) );
no02f80 g567835 ( .a(n_7311), .b(x_in_43_11), .o(n_12599) );
in01f80 g567836 ( .a(n_3222), .o(n_2479) );
na02f80 g567837 ( .a(n_5369), .b(x_in_35_3), .o(n_3222) );
in01f80 g567838 ( .a(n_3328), .o(n_4501) );
no02f80 g567839 ( .a(n_4329), .b(x_in_55_4), .o(n_3328) );
in01f80 g567840 ( .a(n_10790), .o(n_2361) );
na02f80 g567841 ( .a(n_3169), .b(x_in_5_13), .o(n_10790) );
no02f80 g567842 ( .a(n_5156), .b(x_in_35_3), .o(n_2034) );
in01f80 g567843 ( .a(n_3339), .o(n_4467) );
no02f80 g567844 ( .a(n_4745), .b(x_in_63_4), .o(n_3339) );
in01f80 g567845 ( .a(n_5772), .o(n_5856) );
no02f80 g567846 ( .a(n_5986), .b(x_in_45_5), .o(n_5772) );
no02f80 g567847 ( .a(n_2438), .b(x_in_45_2), .o(n_3803) );
no02f80 g567848 ( .a(n_5418), .b(x_in_17_14), .o(n_2842) );
in01f80 g567849 ( .a(n_4446), .o(n_4448) );
no02f80 g567850 ( .a(n_2438), .b(x_in_45_4), .o(n_4446) );
no02f80 g567851 ( .a(n_3887), .b(x_in_21_12), .o(n_3313) );
in01f80 g567852 ( .a(n_2406), .o(n_2407) );
no02f80 g567853 ( .a(n_5977), .b(x_in_21_9), .o(n_2406) );
in01f80 g567854 ( .a(n_2334), .o(n_6935) );
na02f80 g567855 ( .a(n_4794), .b(x_in_17_12), .o(n_2334) );
in01f80 g567856 ( .a(n_4412), .o(n_3673) );
na02f80 g567857 ( .a(n_3445), .b(x_in_47_5), .o(n_4412) );
in01f80 g567858 ( .a(n_12596), .o(n_2379) );
na02f80 g567859 ( .a(n_7336), .b(x_in_7_14), .o(n_12596) );
in01f80 g567860 ( .a(n_12817), .o(n_12815) );
na02f80 g567861 ( .a(n_7765), .b(x_in_19_14), .o(n_12817) );
na02f80 g567862 ( .a(n_9612), .b(x_in_41_9), .o(n_3019) );
in01f80 g567863 ( .a(n_7683), .o(n_2477) );
na02f80 g567864 ( .a(n_5869), .b(x_in_21_12), .o(n_7683) );
in01f80 g567865 ( .a(n_4432), .o(n_4434) );
no02f80 g567866 ( .a(n_5986), .b(x_in_45_1), .o(n_4432) );
in01f80 g567867 ( .a(n_4159), .o(n_2476) );
no02f80 g567868 ( .a(n_3238), .b(x_in_49_5), .o(n_4159) );
no02f80 g567869 ( .a(n_9646), .b(x_in_17_3), .o(n_6929) );
na02f80 g567870 ( .a(n_9327), .b(x_in_41_8), .o(n_3252) );
in01f80 g567871 ( .a(n_4440), .o(n_3421) );
na02f80 g567872 ( .a(n_3739), .b(x_in_31_5), .o(n_4440) );
na02f80 g567873 ( .a(n_4654), .b(x_in_37_1), .o(n_2278) );
in01f80 g567874 ( .a(n_2474), .o(n_2475) );
no02f80 g567875 ( .a(n_5556), .b(x_in_19_14), .o(n_2474) );
no02f80 g567876 ( .a(n_7304), .b(x_in_7_7), .o(n_2848) );
in01f80 g567877 ( .a(n_2869), .o(n_3789) );
no02f80 g567878 ( .a(n_7285), .b(x_in_7_14), .o(n_2869) );
in01f80 g567879 ( .a(n_2776), .o(n_2777) );
na02f80 g567880 ( .a(x_in_23_9), .b(n_15183), .o(n_2776) );
na02f80 g567881 ( .a(x_in_23_2), .b(FE_OFN290_n_27194), .o(n_7283) );
na02f80 g567882 ( .a(x_in_55_2), .b(n_4276), .o(n_7364) );
na02f80 g567883 ( .a(x_in_15_2), .b(FE_OFN290_n_27194), .o(n_7359) );
in01f80 g567884 ( .a(n_4201), .o(n_4202) );
na02f80 g567885 ( .a(x_in_15_7), .b(FE_OFN355_n_4860), .o(n_4201) );
in01f80 g567886 ( .a(n_4211), .o(n_4212) );
na02f80 g567887 ( .a(x_in_31_7), .b(FE_OFN1171_n_4860), .o(n_4211) );
in01f80 g567888 ( .a(n_2796), .o(n_2797) );
na02f80 g567889 ( .a(x_in_63_7), .b(FE_OFN1115_rst), .o(n_2796) );
in01f80 g567890 ( .a(n_2799), .o(n_2800) );
na02f80 g567891 ( .a(x_in_63_5), .b(FE_OFN1106_rst), .o(n_2799) );
na02f80 g567892 ( .a(x_in_63_2), .b(n_4276), .o(n_7347) );
in01f80 g567893 ( .a(n_4301), .o(n_4302) );
na02f80 g567894 ( .a(x_in_31_9), .b(FE_OFN1171_n_4860), .o(n_4301) );
in01f80 g567895 ( .a(n_4299), .o(n_4300) );
na02f80 g567896 ( .a(x_in_55_9), .b(FE_OFN86_n_14586), .o(n_4299) );
in01f80 g567897 ( .a(n_4297), .o(n_4298) );
na02f80 g567898 ( .a(x_in_63_9), .b(n_4860), .o(n_4297) );
na02f80 g567899 ( .a(x_in_31_2), .b(n_27194), .o(n_7446) );
in01f80 g567900 ( .a(n_4221), .o(n_4222) );
na02f80 g567901 ( .a(x_in_15_5), .b(n_4860), .o(n_4221) );
na02f80 g567902 ( .a(x_in_47_2), .b(FE_OFN290_n_27194), .o(n_7254) );
in01f80 g567903 ( .a(n_4233), .o(n_4234) );
na02f80 g567904 ( .a(x_in_23_5), .b(FE_OFN1155_n_14586), .o(n_4233) );
in01f80 g567905 ( .a(n_2859), .o(n_2860) );
na02f80 g567906 ( .a(x_in_23_7), .b(n_15183), .o(n_2859) );
in01f80 g567907 ( .a(n_2821), .o(n_2822) );
na02f80 g567908 ( .a(x_in_15_9), .b(FE_OFN1112_rst), .o(n_2821) );
na02f80 g567909 ( .a(x_in_27_3), .b(n_4276), .o(n_7250) );
in01f80 g567910 ( .a(n_2823), .o(n_2824) );
na02f80 g567911 ( .a(x_in_47_9), .b(FE_OFN34_n_15183), .o(n_2823) );
in01f80 g567912 ( .a(n_3348), .o(n_3349) );
na02f80 g567913 ( .a(x_in_55_7), .b(n_15183), .o(n_3348) );
in01f80 g567914 ( .a(n_4295), .o(n_4296) );
na02f80 g567915 ( .a(x_in_47_7), .b(n_4860), .o(n_4295) );
in01f80 g567916 ( .a(n_4293), .o(n_4294) );
na02f80 g567917 ( .a(x_in_55_5), .b(FE_OFN86_n_14586), .o(n_4293) );
in01f80 g567918 ( .a(n_4523), .o(n_4524) );
no02f80 g567919 ( .a(n_7272), .b(x_in_63_7), .o(n_4523) );
no02f80 g567920 ( .a(n_2421), .b(x_in_27_4), .o(n_3634) );
in01f80 g567921 ( .a(n_4469), .o(n_4470) );
no02f80 g567922 ( .a(n_6711), .b(x_in_63_5), .o(n_4469) );
in01f80 g567923 ( .a(n_4459), .o(n_3468) );
na02f80 g567924 ( .a(n_6483), .b(x_in_31_7), .o(n_4459) );
in01f80 g567925 ( .a(n_4642), .o(n_2447) );
na02f80 g567926 ( .a(n_3186), .b(x_in_49_9), .o(n_4642) );
in01f80 g567927 ( .a(n_4224), .o(n_4225) );
no02f80 g567928 ( .a(n_6685), .b(x_in_55_5), .o(n_4224) );
in01f80 g567929 ( .a(n_4884), .o(n_4885) );
no02f80 g567930 ( .a(n_8200), .b(x_in_31_7), .o(n_4884) );
in01f80 g567931 ( .a(n_7613), .o(n_2367) );
no02f80 g567932 ( .a(n_5888), .b(x_in_5_10), .o(n_7613) );
in01f80 g567933 ( .a(n_4430), .o(n_3666) );
na02f80 g567934 ( .a(n_6685), .b(x_in_55_7), .o(n_4430) );
in01f80 g567935 ( .a(n_6907), .o(n_2487) );
na02f80 g567936 ( .a(n_5296), .b(x_in_5_7), .o(n_6907) );
in01f80 g567937 ( .a(n_6802), .o(n_2296) );
no02f80 g567938 ( .a(n_5388), .b(x_in_5_8), .o(n_6802) );
no02f80 g567939 ( .a(n_23944), .b(x_in_5_14), .o(n_15752) );
in01f80 g567940 ( .a(n_6015), .o(n_4111) );
no02f80 g567941 ( .a(n_6483), .b(x_in_31_5), .o(n_6015) );
in01f80 g567942 ( .a(n_8071), .o(n_4103) );
no02f80 g567943 ( .a(n_11037), .b(x_in_15_9), .o(n_8071) );
in01f80 g567944 ( .a(n_8063), .o(n_3508) );
no02f80 g567945 ( .a(n_11040), .b(x_in_55_9), .o(n_8063) );
in01f80 g567946 ( .a(n_8067), .o(n_4106) );
no02f80 g567947 ( .a(n_11696), .b(x_in_63_9), .o(n_8067) );
in01f80 g567948 ( .a(n_3054), .o(n_2519) );
na02f80 g567949 ( .a(n_2421), .b(x_in_27_4), .o(n_3054) );
in01f80 g567950 ( .a(n_2760), .o(n_4472) );
no02f80 g567951 ( .a(n_10916), .b(x_in_63_8), .o(n_2760) );
in01f80 g567952 ( .a(n_3301), .o(n_4310) );
no02f80 g567953 ( .a(n_10918), .b(x_in_23_8), .o(n_3301) );
no02f80 g567954 ( .a(n_2512), .b(x_in_57_4), .o(n_6892) );
in01f80 g567955 ( .a(n_6766), .o(n_2632) );
no02f80 g567956 ( .a(n_5849), .b(x_in_37_10), .o(n_6766) );
in01f80 g567957 ( .a(n_2529), .o(n_2530) );
na02f80 g567958 ( .a(n_3193), .b(x_in_53_11), .o(n_2529) );
in01f80 g567959 ( .a(n_6805), .o(n_2300) );
no02f80 g567960 ( .a(n_6000), .b(x_in_5_7), .o(n_6805) );
no02f80 g567961 ( .a(n_4654), .b(x_in_37_4), .o(n_2286) );
in01f80 g567962 ( .a(n_3295), .o(n_4532) );
no02f80 g567963 ( .a(n_10913), .b(x_in_47_8), .o(n_3295) );
in01f80 g567964 ( .a(n_2301), .o(n_5108) );
na02f80 g567965 ( .a(n_3191), .b(x_in_49_7), .o(n_2301) );
in01f80 g567966 ( .a(n_7710), .o(n_2473) );
na02f80 g567967 ( .a(n_5860), .b(x_in_21_10), .o(n_7710) );
na02f80 g567968 ( .a(n_3193), .b(x_in_53_14), .o(n_3235) );
no02f80 g567969 ( .a(n_2240), .b(x_in_37_3), .o(n_2242) );
in01f80 g567970 ( .a(n_4403), .o(n_4402) );
na02f80 g567971 ( .a(n_3193), .b(x_in_53_12), .o(n_4403) );
no02f80 g567972 ( .a(n_2240), .b(x_in_37_6), .o(n_2109) );
in01f80 g567973 ( .a(n_4373), .o(n_2302) );
no02f80 g567974 ( .a(n_7904), .b(x_in_15_6), .o(n_4373) );
no02f80 g567975 ( .a(n_5095), .b(x_in_49_7), .o(n_5107) );
in01f80 g567976 ( .a(n_6023), .o(n_4428) );
no02f80 g567977 ( .a(n_6492), .b(x_in_15_7), .o(n_6023) );
in01f80 g567978 ( .a(n_8058), .o(n_3695) );
no02f80 g567979 ( .a(n_11698), .b(x_in_31_9), .o(n_8058) );
no02f80 g567980 ( .a(n_7320), .b(x_in_7_8), .o(n_2844) );
in01f80 g567981 ( .a(n_7681), .o(n_2303) );
no02f80 g567982 ( .a(n_5884), .b(x_in_37_4), .o(n_7681) );
in01f80 g567983 ( .a(n_6923), .o(n_2414) );
no02f80 g567984 ( .a(n_5754), .b(x_in_5_9), .o(n_6923) );
na02f80 g567985 ( .a(n_2240), .b(x_in_37_2), .o(n_2082) );
in01f80 g567986 ( .a(n_4498), .o(n_4499) );
no02f80 g567987 ( .a(n_7241), .b(x_in_47_7), .o(n_4498) );
in01f80 g567988 ( .a(n_6889), .o(n_2304) );
no02f80 g567989 ( .a(n_4668), .b(x_in_57_3), .o(n_6889) );
no02f80 g567990 ( .a(n_7765), .b(x_in_19_13), .o(n_3022) );
in01f80 g567991 ( .a(n_6021), .o(n_3670) );
no02f80 g567992 ( .a(n_7270), .b(x_in_23_7), .o(n_6021) );
in01f80 g567993 ( .a(n_6013), .o(n_4240) );
no02f80 g567994 ( .a(n_6687), .b(x_in_15_5), .o(n_6013) );
in01f80 g567995 ( .a(n_4199), .o(n_3451) );
na02f80 g567996 ( .a(n_6711), .b(x_in_63_7), .o(n_4199) );
no02f80 g567997 ( .a(n_3188), .b(x_in_49_10), .o(n_5125) );
in01f80 g567998 ( .a(n_4444), .o(n_3373) );
na02f80 g567999 ( .a(n_6689), .b(x_in_23_7), .o(n_4444) );
na02f80 g568000 ( .a(n_5869), .b(x_in_21_7), .o(n_3084) );
in01f80 g568001 ( .a(n_4389), .o(n_4390) );
no02f80 g568002 ( .a(n_6689), .b(x_in_23_5), .o(n_4389) );
no02f80 g568003 ( .a(n_3193), .b(x_in_53_14), .o(n_3362) );
in01f80 g568004 ( .a(n_2306), .o(n_2307) );
no02f80 g568005 ( .a(n_7304), .b(x_in_7_9), .o(n_2306) );
in01f80 g568006 ( .a(n_2576), .o(n_2577) );
na02f80 g568007 ( .a(n_3036), .b(x_in_21_10), .o(n_2576) );
in01f80 g568008 ( .a(n_8069), .o(n_4116) );
no02f80 g568009 ( .a(n_11034), .b(x_in_47_9), .o(n_8069) );
in01f80 g568010 ( .a(n_2898), .o(n_8299) );
na02f80 g568011 ( .a(n_3011), .b(x_in_37_4), .o(n_2898) );
in01f80 g568012 ( .a(n_3307), .o(n_4509) );
no02f80 g568013 ( .a(n_10915), .b(x_in_55_8), .o(n_3307) );
in01f80 g568014 ( .a(n_4370), .o(n_4130) );
na02f80 g568015 ( .a(n_6492), .b(x_in_15_9), .o(n_4370) );
in01f80 g568016 ( .a(n_4548), .o(n_4549) );
no02f80 g568017 ( .a(n_6683), .b(x_in_47_5), .o(n_4548) );
in01f80 g568018 ( .a(n_8061), .o(n_3698) );
no02f80 g568019 ( .a(n_11041), .b(x_in_23_9), .o(n_8061) );
na02f80 g568020 ( .a(n_5754), .b(x_in_5_14), .o(n_8690) );
in01f80 g568021 ( .a(n_3115), .o(n_4485) );
no02f80 g568022 ( .a(n_10914), .b(x_in_31_8), .o(n_3115) );
in01f80 g568023 ( .a(n_4496), .o(n_4135) );
na02f80 g568024 ( .a(n_6683), .b(x_in_47_7), .o(n_4496) );
in01f80 g568025 ( .a(n_2883), .o(n_4605) );
na02f80 g568026 ( .a(n_3188), .b(x_in_49_6), .o(n_2883) );
in01f80 g568027 ( .a(n_6022), .o(n_4513) );
no02f80 g568028 ( .a(n_7315), .b(x_in_55_7), .o(n_6022) );
in01f80 g568029 ( .a(n_2436), .o(n_2437) );
no02f80 g568030 ( .a(n_2583), .b(x_in_41_4), .o(n_2436) );
in01f80 g568031 ( .a(n_4141), .o(n_4142) );
na02f80 g568032 ( .a(x_in_31_5), .b(FE_OFN1171_n_4860), .o(n_4141) );
in01f80 g568033 ( .a(n_4305), .o(n_4306) );
na02f80 g568034 ( .a(x_in_47_5), .b(n_4860), .o(n_4305) );
in01f80 g568035 ( .a(n_2591), .o(n_2592) );
na02f80 g568036 ( .a(n_2363), .b(x_in_59_8), .o(n_2591) );
in01f80 g568037 ( .a(n_6912), .o(n_2416) );
no02f80 g568038 ( .a(n_5313), .b(x_in_57_9), .o(n_6912) );
in01f80 g568039 ( .a(n_3095), .o(n_5408) );
no02f80 g568040 ( .a(n_5962), .b(x_in_37_7), .o(n_3095) );
no02f80 g568041 ( .a(n_5699), .b(x_in_59_6), .o(n_3632) );
in01f80 g568042 ( .a(n_3040), .o(n_7700) );
no02f80 g568043 ( .a(n_5881), .b(x_in_37_6), .o(n_3040) );
no02f80 g568044 ( .a(n_5940), .b(x_in_19_9), .o(n_3033) );
no02f80 g568045 ( .a(n_2363), .b(x_in_59_8), .o(n_3358) );
no02f80 g568046 ( .a(n_5939), .b(x_in_19_6), .o(n_3239) );
na02f80 g568047 ( .a(n_5839), .b(x_in_61_6), .o(n_3083) );
in01f80 g568048 ( .a(n_6881), .o(n_2470) );
no02f80 g568049 ( .a(n_3409), .b(x_in_57_8), .o(n_6881) );
no02f80 g568050 ( .a(n_2652), .b(x_in_35_7), .o(n_3449) );
na02f80 g568051 ( .a(n_5691), .b(x_in_59_7), .o(n_3368) );
no02f80 g568052 ( .a(n_5293), .b(x_in_43_5), .o(n_3448) );
in01f80 g568053 ( .a(n_6814), .o(n_2514) );
no02f80 g568054 ( .a(n_2627), .b(x_in_57_6), .o(n_6814) );
in01f80 g568055 ( .a(n_7679), .o(n_2689) );
na02f80 g568056 ( .a(n_5742), .b(x_in_37_7), .o(n_7679) );
in01f80 g568057 ( .a(n_2468), .o(n_2469) );
na02f80 g568058 ( .a(n_5180), .b(x_in_51_2), .o(n_2468) );
in01f80 g568059 ( .a(n_2638), .o(n_2639) );
no02f80 g568060 ( .a(n_5242), .b(x_in_61_6), .o(n_2638) );
na02f80 g568061 ( .a(n_5244), .b(x_in_19_10), .o(n_3047) );
in01f80 g568062 ( .a(n_3255), .o(n_2311) );
na02f80 g568063 ( .a(n_2652), .b(x_in_35_7), .o(n_3255) );
na02f80 g568064 ( .a(n_5554), .b(x_in_19_6), .o(n_3026) );
no02f80 g568065 ( .a(n_5537), .b(x_in_19_11), .o(n_3108) );
in01f80 g568066 ( .a(n_2466), .o(n_2467) );
na02f80 g568067 ( .a(n_5699), .b(x_in_59_6), .o(n_2466) );
no02f80 g568068 ( .a(n_5761), .b(x_in_61_5), .o(n_2804) );
in01f80 g568069 ( .a(n_2665), .o(n_2666) );
no02f80 g568070 ( .a(n_5691), .b(x_in_59_7), .o(n_2665) );
in01f80 g568071 ( .a(n_2347), .o(n_2348) );
no02f80 g568072 ( .a(n_2668), .b(x_in_59_9), .o(n_2347) );
in01f80 g568073 ( .a(n_11195), .o(n_12688) );
no02f80 g568074 ( .a(n_4847), .b(x_in_61_11), .o(n_11195) );
no02f80 g568075 ( .a(n_5180), .b(x_in_51_2), .o(n_3453) );
in01f80 g568076 ( .a(n_6817), .o(n_2501) );
na02f80 g568077 ( .a(n_4668), .b(x_in_57_7), .o(n_6817) );
no02f80 g568078 ( .a(n_3174), .b(x_in_19_7), .o(n_3034) );
na02f80 g568079 ( .a(n_2668), .b(x_in_59_9), .o(n_3875) );
in01f80 g568080 ( .a(n_2345), .o(n_2346) );
na02f80 g568081 ( .a(n_5293), .b(x_in_43_5), .o(n_2345) );
in01f80 g568082 ( .a(n_7702), .o(n_2465) );
na02f80 g568083 ( .a(n_3409), .b(x_in_57_12), .o(n_7702) );
in01f80 g568084 ( .a(n_6811), .o(n_2335) );
no02f80 g568085 ( .a(n_3245), .b(x_in_57_7), .o(n_6811) );
in01f80 g568086 ( .a(n_2674), .o(n_2675) );
na02f80 g568087 ( .a(n_5761), .b(x_in_61_7), .o(n_2674) );
na02f80 g568088 ( .a(n_3020), .b(x_in_19_8), .o(n_3021) );
na02f80 g568089 ( .a(n_4942), .b(x_in_35_4), .o(n_3784) );
in01f80 g568090 ( .a(n_3305), .o(n_7731) );
na02f80 g568091 ( .a(n_5905), .b(x_in_3_11), .o(n_3305) );
no02f80 g568092 ( .a(n_2550), .b(x_in_53_10), .o(n_2095) );
in01f80 g568093 ( .a(n_7693), .o(n_2464) );
no02f80 g568094 ( .a(n_5872), .b(x_in_21_9), .o(n_7693) );
in01f80 g568095 ( .a(n_7687), .o(n_2463) );
na02f80 g568096 ( .a(n_8557), .b(x_in_21_6), .o(n_7687) );
in01f80 g568097 ( .a(n_7650), .o(n_2462) );
no02f80 g568098 ( .a(n_5860), .b(x_in_21_6), .o(n_7650) );
no02f80 g568099 ( .a(n_4180), .b(x_in_37_9), .o(n_8305) );
na02f80 g568100 ( .a(n_5515), .b(x_in_3_8), .o(n_7655) );
in01f80 g568101 ( .a(n_2297), .o(n_2298) );
no02f80 g568102 ( .a(n_5900), .b(x_in_21_8), .o(n_2297) );
in01f80 g568103 ( .a(n_6374), .o(n_6376) );
na02f80 g568104 ( .a(n_2626), .b(x_in_53_6), .o(n_6374) );
na02f80 g568105 ( .a(n_8929), .b(x_in_61_5), .o(n_2901) );
in01f80 g568106 ( .a(n_2370), .o(n_2371) );
no02f80 g568107 ( .a(n_5914), .b(x_in_21_9), .o(n_2370) );
na02f80 g568108 ( .a(n_5275), .b(x_in_59_5), .o(n_3691) );
no02f80 g568109 ( .a(n_5860), .b(x_in_21_5), .o(n_3248) );
in01f80 g568110 ( .a(n_3042), .o(n_5567) );
no02f80 g568111 ( .a(n_2653), .b(x_in_53_9), .o(n_3042) );
no02f80 g568112 ( .a(n_4021), .b(x_in_17_2), .o(n_7728) );
in01f80 g568113 ( .a(n_6382), .o(n_6383) );
no02f80 g568114 ( .a(n_2550), .b(x_in_53_8), .o(n_6382) );
in01f80 g568115 ( .a(n_2997), .o(n_7669) );
na02f80 g568116 ( .a(n_5757), .b(x_in_3_9), .o(n_2997) );
in01f80 g568117 ( .a(n_2404), .o(n_2405) );
na02f80 g568118 ( .a(n_5860), .b(x_in_21_11), .o(n_2404) );
na02f80 g568119 ( .a(n_5524), .b(x_in_3_10), .o(n_7645) );
in01f80 g568120 ( .a(n_2340), .o(n_2341) );
na02f80 g568121 ( .a(n_5369), .b(x_in_35_9), .o(n_2340) );
in01f80 g568122 ( .a(n_2312), .o(n_2313) );
na02f80 g568123 ( .a(n_3036), .b(x_in_21_4), .o(n_2312) );
no02f80 g568124 ( .a(n_4939), .b(x_in_35_5), .o(n_3353) );
no02f80 g568125 ( .a(n_5271), .b(x_in_59_5), .o(n_3477) );
no02f80 g568126 ( .a(n_8524), .b(x_in_35_8), .o(n_3543) );
in01f80 g568127 ( .a(n_2801), .o(n_6797) );
no02f80 g568128 ( .a(n_5247), .b(x_in_3_10), .o(n_2801) );
in01f80 g568129 ( .a(n_4857), .o(n_6378) );
no02f80 g568130 ( .a(n_3038), .b(x_in_53_3), .o(n_4857) );
in01f80 g568131 ( .a(n_3257), .o(n_2375) );
na02f80 g568132 ( .a(n_4939), .b(x_in_35_5), .o(n_3257) );
in01f80 g568133 ( .a(n_3037), .o(n_7690) );
no02f80 g568134 ( .a(n_3036), .b(x_in_21_5), .o(n_3037) );
in01f80 g568135 ( .a(n_2380), .o(n_2381) );
no02f80 g568136 ( .a(n_7320), .b(x_in_7_10), .o(n_2380) );
in01f80 g568137 ( .a(n_6362), .o(n_6360) );
no02f80 g568138 ( .a(n_2654), .b(x_in_53_7), .o(n_6362) );
in01f80 g568139 ( .a(n_2383), .o(n_2384) );
na02f80 g568140 ( .a(n_3608), .b(x_in_61_4), .o(n_2383) );
no02f80 g568141 ( .a(n_3887), .b(x_in_21_6), .o(n_3334) );
in01f80 g568142 ( .a(n_5633), .o(n_2388) );
na02f80 g568143 ( .a(n_3038), .b(x_in_53_5), .o(n_5633) );
no02f80 g568144 ( .a(n_8165), .b(x_in_7_9), .o(n_2728) );
na02f80 g568145 ( .a(n_5963), .b(x_in_3_7), .o(n_7697) );
no02f80 g568146 ( .a(n_2525), .b(x_in_53_8), .o(n_2085) );
in01f80 g568147 ( .a(n_2355), .o(n_2356) );
na02f80 g568148 ( .a(n_5242), .b(x_in_61_4), .o(n_2355) );
in01f80 g568149 ( .a(n_2396), .o(n_2397) );
no02f80 g568150 ( .a(n_5275), .b(x_in_59_5), .o(n_2396) );
na02f80 g568151 ( .a(n_5931), .b(x_in_3_6), .o(n_7380) );
in01f80 g568152 ( .a(n_3090), .o(n_2399) );
na02f80 g568153 ( .a(n_5032), .b(x_in_35_9), .o(n_3090) );
in01f80 g568154 ( .a(n_3211), .o(n_8010) );
no02f80 g568155 ( .a(n_3887), .b(x_in_21_7), .o(n_3211) );
na02f80 g568156 ( .a(n_2651), .b(x_in_53_5), .o(n_2108) );
na02f80 g568157 ( .a(n_5872), .b(x_in_21_8), .o(n_3330) );
no02f80 g568158 ( .a(n_5032), .b(x_in_35_9), .o(n_3386) );
in01f80 g568159 ( .a(n_2359), .o(n_2360) );
no02f80 g568160 ( .a(n_4942), .b(x_in_35_4), .o(n_2359) );
in01f80 g568161 ( .a(n_6369), .o(n_6367) );
no02f80 g568162 ( .a(n_2525), .b(x_in_53_6), .o(n_6369) );
in01f80 g568163 ( .a(n_3321), .o(n_2690) );
na02f80 g568164 ( .a(n_5247), .b(x_in_3_11), .o(n_3321) );
na02f80 g568165 ( .a(n_6781), .b(x_in_21_6), .o(n_2888) );
no02f80 g568166 ( .a(n_2654), .b(x_in_53_9), .o(n_2279) );
no02f80 g568167 ( .a(n_2651), .b(x_in_53_7), .o(n_2070) );
na02f80 g568168 ( .a(n_8557), .b(x_in_21_7), .o(n_3223) );
na02f80 g568169 ( .a(n_8929), .b(x_in_61_3), .o(n_2906) );
in01f80 g568170 ( .a(n_2460), .o(n_2461) );
na02f80 g568171 ( .a(n_5914), .b(x_in_21_3), .o(n_2460) );
no02f80 g568172 ( .a(n_5369), .b(x_in_35_9), .o(n_3366) );
in01f80 g568173 ( .a(n_2827), .o(n_2459) );
na02f80 g568174 ( .a(n_8524), .b(x_in_35_8), .o(n_2827) );
na02f80 g568175 ( .a(n_5742), .b(x_in_37_3), .o(n_2253) );
no02f80 g568176 ( .a(n_5827), .b(x_in_53_4), .o(n_2071) );
in01f80 g568177 ( .a(n_8303), .o(n_2426) );
na02f80 g568178 ( .a(n_4654), .b(x_in_37_5), .o(n_8303) );
in01f80 g568179 ( .a(n_2457), .o(n_2458) );
no02f80 g568180 ( .a(n_5839), .b(x_in_61_8), .o(n_2457) );
in01f80 g568181 ( .a(n_2806), .o(n_7658) );
na02f80 g568182 ( .a(n_5881), .b(x_in_37_10), .o(n_2806) );
no02f80 g568183 ( .a(n_4937), .b(x_in_61_7), .o(n_3332) );
in01f80 g568184 ( .a(n_3031), .o(n_7665) );
na02f80 g568185 ( .a(n_5825), .b(x_in_3_5), .o(n_3031) );
in01f80 g568186 ( .a(n_7675), .o(n_7677) );
no02f80 g568187 ( .a(n_2548), .b(x_in_53_14), .o(n_7675) );
no02f80 g568188 ( .a(n_7434), .b(x_in_21_4), .o(n_2118) );
no02f80 g568189 ( .a(n_9651), .b(x_in_17_5), .o(n_6898) );
in01f80 g568190 ( .a(n_3041), .o(n_7707) );
no02f80 g568191 ( .a(n_8557), .b(x_in_21_2), .o(n_3041) );
in01f80 g568192 ( .a(n_2791), .o(n_7715) );
no02f80 g568193 ( .a(n_5900), .b(x_in_21_3), .o(n_2791) );
na02f80 g568194 ( .a(n_5360), .b(x_in_17_5), .o(n_3046) );
no02f80 g568195 ( .a(n_6781), .b(x_in_21_5), .o(n_2282) );
in01f80 g568196 ( .a(n_2621), .o(n_2622) );
no02f80 g568197 ( .a(n_4914), .b(x_in_61_10), .o(n_2621) );
no02f80 g568198 ( .a(n_3833), .b(x_in_61_9), .o(n_3081) );
in01f80 g568199 ( .a(n_2449), .o(n_2450) );
na02f80 g568200 ( .a(n_4914), .b(x_in_61_8), .o(n_2449) );
in01f80 g568201 ( .a(n_4621), .o(n_2623) );
na02f80 g568202 ( .a(n_5244), .b(x_in_19_11), .o(n_4621) );
na02f80 g568203 ( .a(n_4937), .b(x_in_61_9), .o(n_3078) );
na02f80 g568204 ( .a(x_in_43_4), .b(n_4276), .o(n_6481) );
no02f80 g568205 ( .a(n_3792), .b(x_in_51_4), .o(n_3331) );
na02f80 g568206 ( .a(n_5415), .b(x_in_17_9), .o(n_3200) );
no02f80 g568207 ( .a(n_9654), .b(x_in_17_7), .o(n_6878) );
in01f80 g568208 ( .a(n_2455), .o(n_2456) );
no02f80 g568209 ( .a(n_5979), .b(x_in_51_5), .o(n_2455) );
in01f80 g568210 ( .a(n_4540), .o(n_3638) );
no02f80 g568211 ( .a(n_5418), .b(x_in_17_12), .o(n_4540) );
in01f80 g568212 ( .a(n_6843), .o(n_2454) );
no02f80 g568213 ( .a(n_5415), .b(x_in_17_10), .o(n_6843) );
na02f80 g568214 ( .a(n_5360), .b(x_in_17_10), .o(n_6901) );
na02f80 g568215 ( .a(n_5359), .b(x_in_17_7), .o(n_3345) );
na02f80 g568216 ( .a(n_9651), .b(x_in_17_4), .o(n_2841) );
na02f80 g568217 ( .a(n_10477), .b(x_in_17_10), .o(n_3050) );
in01f80 g568218 ( .a(n_2734), .o(n_4801) );
na02f80 g568219 ( .a(n_12635), .b(x_in_33_11), .o(n_2734) );
na02f80 g568220 ( .a(n_9654), .b(x_in_17_6), .o(n_3336) );
na02f80 g568221 ( .a(n_12178), .b(x_in_33_12), .o(n_2735) );
no02f80 g568222 ( .a(n_5418), .b(x_in_17_9), .o(n_6872) );
na02f80 g568223 ( .a(n_5418), .b(x_in_17_8), .o(n_2830) );
no02f80 g568224 ( .a(n_5362), .b(x_in_17_4), .o(n_6869) );
no02f80 g568225 ( .a(n_5360), .b(x_in_17_6), .o(n_6846) );
in01f80 g568226 ( .a(x_out_29_6), .o(n_1122) );
in01f80 g568227 ( .a(x_out_27_27), .o(n_1744) );
in01f80 g568228 ( .a(x_out_38_0), .o(n_1519) );
in01f80 g568229 ( .a(x_out_55_9), .o(n_771) );
in01f80 g568230 ( .a(x_out_35_21), .o(n_1251) );
in01f80 g568231 ( .a(x_out_42_31), .o(n_1158) );
in01f80 g568232 ( .a(x_out_42_4), .o(n_690) );
in01f80 g568233 ( .a(x_out_3_9), .o(n_1118) );
in01f80 g568234 ( .a(x_out_6_25), .o(n_1787) );
in01f80 g568235 ( .a(x_out_7_0), .o(n_125) );
in01f80 g568236 ( .a(x_out_40_6), .o(n_1544) );
in01f80 g568237 ( .a(x_out_55_3), .o(n_118) );
in01f80 g568238 ( .a(x_out_3_20), .o(n_1062) );
in01f80 g568239 ( .a(x_out_22_20), .o(n_541) );
in01f80 g568240 ( .a(x_out_14_27), .o(n_1432) );
in01f80 g568241 ( .a(x_out_60_26), .o(n_576) );
in01f80 g568242 ( .a(x_out_10_21), .o(n_1305) );
in01f80 g568243 ( .a(x_out_16_29), .o(n_499) );
in01f80 g568244 ( .a(x_out_59_10), .o(n_1891) );
in01f80 g568245 ( .a(x_out_38_21), .o(n_1411) );
in01f80 g568246 ( .a(x_out_26_33), .o(n_809) );
in01f80 g568247 ( .a(x_out_6_1), .o(n_829) );
in01f80 g568248 ( .a(x_out_52_13), .o(n_1093) );
in01f80 g568249 ( .a(x_out_49_27), .o(n_87) );
in01f80 g568250 ( .a(x_out_10_0), .o(n_107) );
in01f80 g568251 ( .a(x_out_27_31), .o(n_1393) );
in01f80 g568252 ( .a(x_out_21_12), .o(n_163) );
in01f80 g568253 ( .a(x_out_43_11), .o(n_506) );
in01f80 g568254 ( .a(x_out_29_26), .o(n_807) );
in01f80 g568255 ( .a(x_out_62_12), .o(n_1240) );
in01f80 g568256 ( .a(x_out_55_23), .o(n_573) );
in01f80 g568257 ( .a(x_out_59_7), .o(n_1739) );
in01f80 g568258 ( .a(x_out_5_28), .o(n_436) );
in01f80 g568259 ( .a(x_out_25_9), .o(n_481) );
in01f80 g568260 ( .a(x_out_41_20), .o(n_969) );
in01f80 g568261 ( .a(x_out_29_24), .o(n_1468) );
in01f80 g568262 ( .a(x_out_5_29), .o(n_1778) );
in01f80 g568263 ( .a(x_out_18_30), .o(n_1589) );
in01f80 g568264 ( .a(x_out_62_11), .o(n_1687) );
in01f80 g568265 ( .a(x_out_63_32), .o(n_82) );
in01f80 g568266 ( .a(x_out_23_22), .o(n_1577) );
in01f80 g568267 ( .a(x_out_23_5), .o(n_1079) );
in01f80 g568268 ( .a(x_out_13_7), .o(n_170) );
in01f80 g568269 ( .a(x_out_16_11), .o(n_842) );
in01f80 g568270 ( .a(x_out_16_32), .o(n_1695) );
in01f80 g568271 ( .a(x_out_26_10), .o(n_1727) );
in01f80 g568272 ( .a(x_out_26_28), .o(n_320) );
in01f80 g568273 ( .a(x_out_31_3), .o(n_801) );
in01f80 g568274 ( .a(x_out_15_14), .o(n_828) );
in01f80 g568275 ( .a(x_out_23_29), .o(n_351) );
in01f80 g568276 ( .a(x_out_21_20), .o(n_1591) );
in01f80 g568277 ( .a(x_out_34_4), .o(n_1507) );
in01f80 g568278 ( .a(x_out_56_1), .o(n_833) );
in01f80 g568279 ( .a(x_out_50_27), .o(n_188) );
in01f80 g568280 ( .a(x_out_55_27), .o(n_291) );
in01f80 g568281 ( .a(x_out_63_18), .o(n_1665) );
in01f80 g568282 ( .a(x_out_18_18), .o(n_452) );
in01f80 g568283 ( .a(x_out_21_32), .o(n_702) );
in01f80 g568284 ( .a(x_out_7_24), .o(n_1465) );
in01f80 g568285 ( .a(x_out_21_10), .o(n_1963) );
in01f80 g568286 ( .a(x_out_56_6), .o(n_257) );
in01f80 g568287 ( .a(x_out_36_27), .o(n_1649) );
in01f80 g568288 ( .a(x_out_10_15), .o(n_1138) );
in01f80 g568289 ( .a(x_out_5_3), .o(n_1919) );
in01f80 g568290 ( .a(x_out_56_2), .o(n_1362) );
in01f80 g568291 ( .a(x_out_55_0), .o(n_1281) );
in01f80 g568292 ( .a(x_out_25_29), .o(n_931) );
in01f80 g568293 ( .a(x_out_41_12), .o(n_115) );
in01f80 g568294 ( .a(x_out_55_4), .o(n_963) );
in01f80 g568295 ( .a(x_out_35_32), .o(n_937) );
in01f80 g568296 ( .a(x_out_30_21), .o(n_737) );
in01f80 g568297 ( .a(x_out_44_33), .o(n_751) );
in01f80 g568298 ( .a(x_out_19_6), .o(n_1873) );
in01f80 g568299 ( .a(x_out_61_15), .o(n_238) );
in01f80 g568300 ( .a(x_out_25_1), .o(n_274) );
in01f80 g568301 ( .a(x_out_57_29), .o(n_1059) );
in01f80 g568302 ( .a(x_out_46_2), .o(n_1167) );
in01f80 g568303 ( .a(x_out_35_4), .o(n_354) );
in01f80 g568304 ( .a(x_out_51_30), .o(n_1288) );
in01f80 g568305 ( .a(x_out_31_26), .o(n_1087) );
in01f80 g568306 ( .a(x_out_0_12), .o(n_1182) );
in01f80 g568307 ( .a(x_out_50_32), .o(n_216) );
in01f80 g568308 ( .a(x_out_31_27), .o(n_525) );
in01f80 g568309 ( .a(x_out_46_4), .o(n_168) );
in01f80 g568310 ( .a(x_out_21_28), .o(n_75) );
in01f80 g568311 ( .a(x_out_46_1), .o(n_834) );
in01f80 g568312 ( .a(x_out_51_4), .o(n_1340) );
in01f80 g568313 ( .a(x_out_23_2), .o(n_1336) );
in01f80 g568314 ( .a(x_out_62_10), .o(n_1851) );
in01f80 g568315 ( .a(x_out_42_15), .o(n_1922) );
in01f80 g568316 ( .a(x_out_11_4), .o(n_384) );
in01f80 g568317 ( .a(x_out_24_21), .o(n_1799) );
in01f80 g568318 ( .a(x_out_55_21), .o(n_1398) );
in01f80 g568319 ( .a(x_out_50_1), .o(n_1437) );
in01f80 g568320 ( .a(x_out_35_0), .o(n_72) );
in01f80 g568321 ( .a(x_out_38_10), .o(n_344) );
in01f80 g568322 ( .a(x_out_57_14), .o(n_735) );
in01f80 g568323 ( .a(x_out_44_15), .o(n_502) );
in01f80 g568324 ( .a(x_out_62_28), .o(n_173) );
in01f80 g568325 ( .a(x_out_49_26), .o(n_358) );
in01f80 g568326 ( .a(x_out_0_2), .o(n_1433) );
in01f80 g568327 ( .a(x_out_12_0), .o(n_1543) );
in01f80 g568328 ( .a(x_out_60_6), .o(n_1225) );
in01f80 g568329 ( .a(x_out_11_26), .o(n_1381) );
in01f80 g568330 ( .a(x_out_46_3), .o(n_1934) );
in01f80 g568331 ( .a(x_out_36_14), .o(n_450) );
in01f80 g568332 ( .a(x_out_6_24), .o(n_1953) );
in01f80 g568333 ( .a(x_out_39_15), .o(n_1326) );
in01f80 g568334 ( .a(x_out_39_7), .o(n_1631) );
in01f80 g568335 ( .a(x_out_4_31), .o(n_756) );
in01f80 g568336 ( .a(x_out_27_8), .o(n_29) );
in01f80 g568337 ( .a(x_out_2_22), .o(n_1961) );
in01f80 g568338 ( .a(x_out_60_22), .o(n_713) );
in01f80 g568339 ( .a(x_out_17_27), .o(n_762) );
in01f80 g568340 ( .a(x_out_49_13), .o(n_1137) );
in01f80 g568341 ( .a(x_out_36_8), .o(n_345) );
in01f80 g568342 ( .a(x_out_21_26), .o(n_237) );
in01f80 g568343 ( .a(x_out_5_14), .o(n_1648) );
in01f80 g568344 ( .a(x_out_24_22), .o(n_1216) );
in01f80 g568345 ( .a(x_out_44_12), .o(n_1908) );
in01f80 g568346 ( .a(x_out_25_25), .o(n_1229) );
in01f80 g568347 ( .a(x_out_51_8), .o(n_1268) );
in01f80 g568348 ( .a(x_out_58_8), .o(n_1482) );
in01f80 g568349 ( .a(x_out_25_27), .o(n_42) );
in01f80 g568350 ( .a(x_out_37_22), .o(n_703) );
in01f80 g568351 ( .a(x_out_56_8), .o(n_307) );
in01f80 g568352 ( .a(x_out_1_11), .o(n_1455) );
in01f80 g568353 ( .a(x_out_19_25), .o(n_37) );
in01f80 g568354 ( .a(x_out_34_12), .o(n_1841) );
in01f80 g568355 ( .a(x_out_4_11), .o(n_924) );
in01f80 g568356 ( .a(x_out_27_26), .o(n_1662) );
in01f80 g568357 ( .a(x_out_60_3), .o(n_719) );
in01f80 g568358 ( .a(x_out_37_0), .o(n_1253) );
in01f80 g568359 ( .a(x_out_22_29), .o(n_1698) );
in01f80 g568360 ( .a(x_out_53_21), .o(n_293) );
in01f80 g568361 ( .a(x_out_54_21), .o(n_1064) );
in01f80 g568362 ( .a(x_out_41_14), .o(n_1256) );
in01f80 g568363 ( .a(x_out_18_27), .o(n_633) );
in01f80 g568364 ( .a(x_out_54_2), .o(n_1218) );
in01f80 g568365 ( .a(x_out_7_30), .o(n_960) );
in01f80 g568366 ( .a(x_out_3_28), .o(n_1569) );
in01f80 g568367 ( .a(x_out_4_23), .o(n_1751) );
in01f80 g568368 ( .a(x_out_44_20), .o(n_1025) );
in01f80 g568369 ( .a(x_out_60_15), .o(n_1923) );
in01f80 g568370 ( .a(x_out_56_25), .o(n_1592) );
in01f80 g568371 ( .a(x_out_59_20), .o(n_694) );
in01f80 g568372 ( .a(x_out_46_9), .o(n_609) );
in01f80 g568373 ( .a(x_out_18_7), .o(n_720) );
in01f80 g568374 ( .a(x_out_12_13), .o(n_1299) );
in01f80 g568375 ( .a(x_out_43_30), .o(n_995) );
in01f80 g568376 ( .a(x_out_3_0), .o(n_194) );
in01f80 g568377 ( .a(x_out_6_5), .o(n_613) );
in01f80 g568378 ( .a(x_out_32_7), .o(n_1888) );
in01f80 g568379 ( .a(x_out_47_18), .o(n_1539) );
in01f80 g568380 ( .a(x_out_8_33), .o(n_18) );
in01f80 g568381 ( .a(x_out_28_8), .o(n_511) );
in01f80 g568382 ( .a(x_out_53_2), .o(n_1474) );
in01f80 g568383 ( .a(x_out_54_13), .o(n_1178) );
in01f80 g568384 ( .a(x_out_63_14), .o(n_8) );
in01f80 g568385 ( .a(x_out_1_18), .o(n_1066) );
in01f80 g568386 ( .a(x_out_14_12), .o(n_1707) );
in01f80 g568387 ( .a(x_out_47_33), .o(n_726) );
in01f80 g568388 ( .a(x_out_49_12), .o(n_602) );
in01f80 g568389 ( .a(x_out_46_20), .o(n_1016) );
in01f80 g568390 ( .a(x_out_48_27), .o(n_455) );
in01f80 g568391 ( .a(x_out_33_33), .o(n_1389) );
in01f80 g568392 ( .a(x_out_22_3), .o(n_184) );
in01f80 g568393 ( .a(x_out_23_12), .o(n_1518) );
in01f80 g568394 ( .a(x_out_15_5), .o(n_240) );
in01f80 g568395 ( .a(x_out_15_13), .o(n_739) );
in01f80 g568396 ( .a(x_out_57_32), .o(n_1024) );
in01f80 g568397 ( .a(x_out_11_32), .o(n_80) );
in01f80 g568398 ( .a(x_out_29_18), .o(n_1499) );
in01f80 g568399 ( .a(x_out_6_29), .o(n_1061) );
in01f80 g568400 ( .a(x_out_4_28), .o(n_1156) );
in01f80 g568401 ( .a(x_out_33_0), .o(n_472) );
in01f80 g568402 ( .a(x_out_47_14), .o(n_1132) );
in01f80 g568403 ( .a(x_out_55_20), .o(n_653) );
in01f80 g568404 ( .a(x_out_41_24), .o(n_1274) );
in01f80 g568405 ( .a(x_out_49_18), .o(n_1410) );
in01f80 g568406 ( .a(x_out_62_6), .o(n_1193) );
in01f80 g568407 ( .a(x_out_35_11), .o(n_516) );
in01f80 g568408 ( .a(x_out_34_22), .o(n_839) );
in01f80 g568409 ( .a(x_out_51_33), .o(n_1536) );
in01f80 g568410 ( .a(x_out_39_8), .o(n_41) );
in01f80 g568411 ( .a(x_out_37_33), .o(n_1295) );
in01f80 g568412 ( .a(x_out_42_9), .o(n_263) );
in01f80 g568413 ( .a(x_out_61_8), .o(n_1918) );
in01f80 g568414 ( .a(x_out_41_15), .o(n_1420) );
in01f80 g568415 ( .a(x_out_45_3), .o(n_1870) );
in01f80 g568416 ( .a(x_out_51_15), .o(n_808) );
in01f80 g568417 ( .a(x_out_57_23), .o(n_1005) );
in01f80 g568418 ( .a(x_out_56_9), .o(n_889) );
in01f80 g568419 ( .a(x_out_46_8), .o(n_1525) );
in01f80 g568420 ( .a(x_out_41_6), .o(n_389) );
in01f80 g568421 ( .a(x_out_53_30), .o(n_421) );
in01f80 g568422 ( .a(x_out_27_6), .o(n_677) );
in01f80 g568423 ( .a(x_out_30_13), .o(n_1653) );
in01f80 g568424 ( .a(x_out_47_10), .o(n_483) );
in01f80 g568425 ( .a(x_out_22_27), .o(n_841) );
in01f80 g568426 ( .a(x_out_24_30), .o(n_226) );
in01f80 g568427 ( .a(x_out_33_4), .o(n_89) );
in01f80 g568428 ( .a(x_out_23_9), .o(n_1259) );
in01f80 g568429 ( .a(x_out_10_27), .o(n_915) );
in01f80 g568430 ( .a(x_out_52_8), .o(n_826) );
in01f80 g568431 ( .a(x_out_49_22), .o(n_350) );
in01f80 g568432 ( .a(x_out_25_4), .o(n_743) );
in01f80 g568433 ( .a(x_out_15_20), .o(n_1335) );
in01f80 g568434 ( .a(x_out_27_30), .o(n_1522) );
in01f80 g568435 ( .a(x_out_7_13), .o(n_1226) );
in01f80 g568436 ( .a(x_out_3_13), .o(n_914) );
in01f80 g568437 ( .a(x_out_47_25), .o(n_646) );
in01f80 g568438 ( .a(x_out_22_5), .o(n_1658) );
in01f80 g568439 ( .a(x_out_27_28), .o(n_457) );
in01f80 g568440 ( .a(x_out_40_23), .o(n_142) );
in01f80 g568441 ( .a(x_out_18_20), .o(n_1619) );
in01f80 g568442 ( .a(x_out_0_0), .o(n_1535) );
in01f80 g568443 ( .a(x_out_40_25), .o(n_977) );
in01f80 g568444 ( .a(x_out_28_22), .o(n_1365) );
in01f80 g568445 ( .a(x_out_51_32), .o(n_1719) );
in01f80 g568446 ( .a(x_out_51_24), .o(n_1332) );
in01f80 g568447 ( .a(x_out_3_2), .o(n_275) );
in01f80 g568448 ( .a(x_out_47_11), .o(n_877) );
in01f80 g568449 ( .a(x_out_36_13), .o(n_1273) );
in01f80 g568450 ( .a(x_out_16_33), .o(n_172) );
in01f80 g568451 ( .a(x_out_57_11), .o(n_412) );
in01f80 g568452 ( .a(x_out_30_0), .o(n_1363) );
in01f80 g568453 ( .a(x_out_36_5), .o(n_1545) );
in01f80 g568454 ( .a(x_out_25_23), .o(n_857) );
in01f80 g568455 ( .a(x_out_62_5), .o(n_867) );
in01f80 g568456 ( .a(x_out_59_28), .o(n_1505) );
in01f80 g568457 ( .a(x_out_1_5), .o(n_177) );
in01f80 g568458 ( .a(x_out_61_18), .o(n_1026) );
in01f80 g568459 ( .a(x_out_4_22), .o(n_760) );
in01f80 g568460 ( .a(x_out_4_25), .o(n_1467) );
in01f80 g568461 ( .a(x_out_49_6), .o(n_504) );
in01f80 g568462 ( .a(x_out_51_10), .o(n_1319) );
in01f80 g568463 ( .a(x_out_14_20), .o(n_127) );
in01f80 g568464 ( .a(x_out_35_1), .o(n_1472) );
in01f80 g568465 ( .a(x_out_58_22), .o(n_104) );
in01f80 g568466 ( .a(x_out_11_10), .o(n_1058) );
in01f80 g568467 ( .a(x_out_25_24), .o(n_1974) );
in01f80 g568468 ( .a(x_out_13_25), .o(n_231) );
in01f80 g568469 ( .a(x_out_6_7), .o(n_1609) );
in01f80 g568470 ( .a(x_out_48_18), .o(n_1260) );
in01f80 g568471 ( .a(x_out_26_2), .o(n_151) );
in01f80 g568472 ( .a(x_out_23_1), .o(n_330) );
in01f80 g568473 ( .a(x_out_53_23), .o(n_721) );
in01f80 g568474 ( .a(x_out_7_14), .o(n_805) );
in01f80 g568475 ( .a(x_out_58_33), .o(n_547) );
in01f80 g568476 ( .a(x_out_24_15), .o(n_855) );
in01f80 g568477 ( .a(x_out_22_2), .o(n_813) );
in01f80 g568478 ( .a(x_out_15_7), .o(n_1669) );
in01f80 g568479 ( .a(x_out_35_29), .o(n_1723) );
in01f80 g568480 ( .a(x_out_38_33), .o(n_306) );
in01f80 g568481 ( .a(x_out_8_3), .o(n_1202) );
in01f80 g568482 ( .a(x_out_41_2), .o(n_564) );
in01f80 g568483 ( .a(x_out_4_7), .o(n_423) );
in01f80 g568484 ( .a(x_out_62_2), .o(n_1354) );
in01f80 g568485 ( .a(x_out_25_15), .o(n_1487) );
in01f80 g568486 ( .a(x_out_22_7), .o(n_1386) );
in01f80 g568487 ( .a(x_out_5_19), .o(n_1485) );
in01f80 g568488 ( .a(x_out_41_27), .o(n_786) );
in01f80 g568489 ( .a(x_out_38_22), .o(n_492) );
in01f80 g568490 ( .a(x_out_30_27), .o(n_891) );
in01f80 g568491 ( .a(x_out_12_32), .o(n_1213) );
in01f80 g568492 ( .a(x_out_50_18), .o(n_1188) );
in01f80 g568493 ( .a(x_out_8_0), .o(n_858) );
in01f80 g568494 ( .a(x_out_11_2), .o(n_1252) );
in01f80 g568495 ( .a(x_out_7_7), .o(n_1282) );
in01f80 g568496 ( .a(x_out_42_24), .o(n_1390) );
in01f80 g568497 ( .a(x_out_44_29), .o(n_812) );
in01f80 g568498 ( .a(x_out_4_18), .o(n_103) );
in01f80 g568499 ( .a(x_out_54_7), .o(n_1532) );
in01f80 g568500 ( .a(x_out_35_13), .o(n_340) );
in01f80 g568501 ( .a(x_out_20_10), .o(n_540) );
in01f80 g568502 ( .a(x_out_62_4), .o(n_77) );
in01f80 g568503 ( .a(x_out_18_28), .o(n_1752) );
in01f80 g568504 ( .a(x_out_49_7), .o(n_1861) );
in01f80 g568505 ( .a(x_out_44_8), .o(n_1017) );
in01f80 g568506 ( .a(x_out_55_14), .o(n_335) );
in01f80 g568507 ( .a(x_out_62_9), .o(n_370) );
in01f80 g568508 ( .a(x_out_26_31), .o(n_1887) );
in01f80 g568509 ( .a(x_out_2_10), .o(n_88) );
in01f80 g568510 ( .a(x_out_31_21), .o(n_1074) );
in01f80 g568511 ( .a(x_out_17_18), .o(n_259) );
in01f80 g568512 ( .a(x_out_36_22), .o(n_58) );
in01f80 g568513 ( .a(x_out_38_11), .o(n_159) );
in01f80 g568514 ( .a(x_out_33_10), .o(n_999) );
in01f80 g568515 ( .a(x_out_17_32), .o(n_959) );
in01f80 g568516 ( .a(x_out_46_25), .o(n_1674) );
in01f80 g568517 ( .a(x_out_59_18), .o(n_128) );
in01f80 g568518 ( .a(x_out_39_28), .o(n_734) );
in01f80 g568519 ( .a(x_out_35_12), .o(n_478) );
in01f80 g568520 ( .a(x_out_12_3), .o(n_92) );
in01f80 g568521 ( .a(x_out_15_11), .o(n_220) );
in01f80 g568522 ( .a(x_out_42_22), .o(n_973) );
in01f80 g568523 ( .a(x_out_59_33), .o(n_21) );
in01f80 g568524 ( .a(x_out_48_33), .o(n_1387) );
in01f80 g568525 ( .a(x_out_22_8), .o(n_1822) );
in01f80 g568526 ( .a(x_out_54_25), .o(n_1359) );
in01f80 g568527 ( .a(x_out_28_15), .o(n_1133) );
in01f80 g568528 ( .a(x_out_11_24), .o(n_904) );
in01f80 g568529 ( .a(x_out_4_4), .o(n_1725) );
in01f80 g568530 ( .a(x_out_57_8), .o(n_1714) );
in01f80 g568531 ( .a(x_out_1_14), .o(n_1165) );
in01f80 g568532 ( .a(x_out_43_29), .o(n_598) );
in01f80 g568533 ( .a(x_out_12_2), .o(n_1426) );
in01f80 g568534 ( .a(x_out_46_13), .o(n_1912) );
in01f80 g568535 ( .a(x_out_47_1), .o(n_532) );
in01f80 g568536 ( .a(x_out_60_5), .o(n_748) );
in01f80 g568537 ( .a(x_out_28_9), .o(n_1832) );
in01f80 g568538 ( .a(x_out_21_4), .o(n_363) );
in01f80 g568539 ( .a(x_out_3_27), .o(n_470) );
in01f80 g568540 ( .a(x_out_26_18), .o(n_1938) );
in01f80 g568541 ( .a(x_out_21_13), .o(n_894) );
in01f80 g568542 ( .a(x_out_35_33), .o(n_317) );
in01f80 g568543 ( .a(x_out_53_20), .o(n_411) );
in01f80 g568544 ( .a(x_out_60_11), .o(n_770) );
in01f80 g568545 ( .a(x_out_26_24), .o(n_1852) );
in01f80 g568546 ( .a(x_out_44_13), .o(n_790) );
in01f80 g568547 ( .a(x_out_49_4), .o(n_1657) );
in01f80 g568548 ( .a(x_out_45_21), .o(n_1680) );
in01f80 g568549 ( .a(x_out_50_8), .o(n_267) );
in01f80 g568550 ( .a(x_out_20_7), .o(n_322) );
in01f80 g568551 ( .a(x_out_39_24), .o(n_1080) );
in01f80 g568552 ( .a(x_out_25_13), .o(n_268) );
in01f80 g568553 ( .a(x_out_56_4), .o(n_443) );
in01f80 g568554 ( .a(x_out_28_0), .o(n_1902) );
in01f80 g568555 ( .a(x_out_28_19), .o(n_1402) );
in01f80 g568556 ( .a(x_out_8_9), .o(n_365) );
in01f80 g568557 ( .a(x_out_1_3), .o(n_233) );
in01f80 g568558 ( .a(x_out_57_0), .o(n_1654) );
in01f80 g568559 ( .a(x_out_31_19), .o(n_1191) );
in01f80 g568560 ( .a(x_out_28_27), .o(n_922) );
in01f80 g568561 ( .a(x_out_47_12), .o(n_933) );
in01f80 g568562 ( .a(x_out_44_11), .o(n_155) );
in01f80 g568563 ( .a(x_out_45_7), .o(n_1899) );
in01f80 g568564 ( .a(x_out_13_26), .o(n_1423) );
in01f80 g568565 ( .a(x_out_29_28), .o(n_7) );
in01f80 g568566 ( .a(x_out_55_5), .o(n_1171) );
in01f80 g568567 ( .a(x_out_8_5), .o(n_116) );
in01f80 g568568 ( .a(x_out_53_24), .o(n_1661) );
in01f80 g568569 ( .a(x_out_59_24), .o(n_1773) );
in01f80 g568570 ( .a(x_out_45_23), .o(n_635) );
in01f80 g568571 ( .a(x_out_22_13), .o(n_53) );
in01f80 g568572 ( .a(x_out_58_5), .o(n_1733) );
in01f80 g568573 ( .a(x_out_18_5), .o(n_766) );
in01f80 g568574 ( .a(x_out_42_3), .o(n_850) );
in01f80 g568575 ( .a(x_out_13_4), .o(n_898) );
in01f80 g568576 ( .a(x_out_34_24), .o(n_1640) );
in01f80 g568577 ( .a(x_out_9_26), .o(n_1430) );
in01f80 g568578 ( .a(x_out_42_25), .o(n_1818) );
in01f80 g568579 ( .a(x_out_25_30), .o(n_1049) );
in01f80 g568580 ( .a(x_out_12_1), .o(n_1811) );
in01f80 g568581 ( .a(x_out_32_9), .o(n_1484) );
in01f80 g568582 ( .a(x_out_37_21), .o(n_414) );
in01f80 g568583 ( .a(x_out_42_2), .o(n_1924) );
in01f80 g568584 ( .a(x_out_40_24), .o(n_1228) );
in01f80 g568585 ( .a(x_out_54_22), .o(n_1515) );
in01f80 g568586 ( .a(x_out_8_23), .o(n_462) );
in01f80 g568587 ( .a(x_out_39_18), .o(n_591) );
in01f80 g568588 ( .a(x_out_15_27), .o(n_161) );
in01f80 g568589 ( .a(x_out_4_1), .o(n_1766) );
in01f80 g568590 ( .a(x_out_55_24), .o(n_1767) );
in01f80 g568591 ( .a(x_out_48_23), .o(n_907) );
in01f80 g568592 ( .a(x_out_1_8), .o(n_36) );
in01f80 g568593 ( .a(x_out_2_26), .o(n_1703) );
in01f80 g568594 ( .a(x_out_5_26), .o(n_617) );
in01f80 g568595 ( .a(x_out_51_2), .o(n_817) );
in01f80 g568596 ( .a(x_out_48_12), .o(n_791) );
in01f80 g568597 ( .a(x_out_23_27), .o(n_245) );
in01f80 g568598 ( .a(x_out_59_12), .o(n_885) );
in01f80 g568599 ( .a(x_out_22_14), .o(n_1618) );
in01f80 g568600 ( .a(x_out_56_22), .o(n_1173) );
in01f80 g568601 ( .a(x_out_33_11), .o(n_1845) );
in01f80 g568602 ( .a(x_out_31_30), .o(n_656) );
in01f80 g568603 ( .a(x_out_23_3), .o(n_1699) );
in01f80 g568604 ( .a(x_out_20_15), .o(n_24) );
in01f80 g568605 ( .a(x_out_18_15), .o(n_749) );
in01f80 g568606 ( .a(x_out_51_18), .o(n_1623) );
in01f80 g568607 ( .a(x_out_15_6), .o(n_1360) );
in01f80 g568608 ( .a(x_out_15_10), .o(n_197) );
in01f80 g568609 ( .a(x_out_33_5), .o(n_1614) );
in01f80 g568610 ( .a(x_out_19_26), .o(n_1014) );
in01f80 g568611 ( .a(x_out_42_0), .o(n_1905) );
in01f80 g568612 ( .a(x_out_60_18), .o(n_1837) );
in01f80 g568613 ( .a(x_out_19_13), .o(n_1749) );
in01f80 g568614 ( .a(x_out_14_23), .o(n_1551) );
in01f80 g568615 ( .a(x_out_2_28), .o(n_792) );
in01f80 g568616 ( .a(x_out_22_21), .o(n_60) );
in01f80 g568617 ( .a(x_out_14_18), .o(n_137) );
in01f80 g568618 ( .a(x_out_57_20), .o(n_555) );
in01f80 g568619 ( .a(x_out_11_18), .o(n_331) );
in01f80 g568620 ( .a(x_out_53_14), .o(n_1019) );
in01f80 g568621 ( .a(x_out_47_2), .o(n_1896) );
in01f80 g568622 ( .a(x_out_37_4), .o(n_1479) );
in01f80 g568623 ( .a(x_out_27_12), .o(n_1043) );
in01f80 g568624 ( .a(x_out_4_32), .o(n_1448) );
in01f80 g568625 ( .a(x_out_7_22), .o(n_375) );
in01f80 g568626 ( .a(x_out_27_14), .o(n_1081) );
in01f80 g568627 ( .a(x_out_8_13), .o(n_1827) );
in01f80 g568628 ( .a(x_out_26_14), .o(n_942) );
in01f80 g568629 ( .a(x_out_55_32), .o(n_552) );
in01f80 g568630 ( .a(x_out_13_13), .o(n_961) );
in01f80 g568631 ( .a(x_out_30_30), .o(n_1394) );
in01f80 g568632 ( .a(x_out_16_19), .o(n_1761) );
in01f80 g568633 ( .a(x_out_22_24), .o(n_1796) );
in01f80 g568634 ( .a(x_out_62_13), .o(n_1279) );
in01f80 g568635 ( .a(x_out_2_12), .o(n_1289) );
in01f80 g568636 ( .a(x_out_23_21), .o(n_1972) );
in01f80 g568637 ( .a(x_out_26_13), .o(n_182) );
in01f80 g568638 ( .a(x_out_18_12), .o(n_1792) );
in01f80 g568639 ( .a(x_out_30_18), .o(n_1671) );
in01f80 g568640 ( .a(x_out_61_7), .o(n_1051) );
in01f80 g568641 ( .a(x_out_37_1), .o(n_954) );
in01f80 g568642 ( .a(x_out_36_7), .o(n_1890) );
in01f80 g568643 ( .a(x_out_5_20), .o(n_34) );
in01f80 g568644 ( .a(x_out_61_1), .o(n_279) );
in01f80 g568645 ( .a(x_out_38_12), .o(n_767) );
in01f80 g568646 ( .a(x_out_54_28), .o(n_1450) );
in01f80 g568647 ( .a(x_out_3_6), .o(n_687) );
in01f80 g568648 ( .a(x_out_7_23), .o(n_469) );
in01f80 g568649 ( .a(x_out_7_1), .o(n_1162) );
in01f80 g568650 ( .a(x_out_21_6), .o(n_1070) );
in01f80 g568651 ( .a(x_out_61_2), .o(n_367) );
in01f80 g568652 ( .a(x_out_53_6), .o(n_324) );
in01f80 g568653 ( .a(x_out_16_14), .o(n_489) );
in01f80 g568654 ( .a(x_out_3_5), .o(n_1159) );
in01f80 g568655 ( .a(x_out_28_31), .o(n_952) );
in01f80 g568656 ( .a(x_out_43_6), .o(n_733) );
in01f80 g568657 ( .a(x_out_17_21), .o(n_1768) );
in01f80 g568658 ( .a(x_out_17_7), .o(n_562) );
in01f80 g568659 ( .a(x_out_45_24), .o(n_1872) );
in01f80 g568660 ( .a(x_out_54_23), .o(n_1730) );
in01f80 g568661 ( .a(x_out_6_26), .o(n_1724) );
in01f80 g568662 ( .a(x_out_32_1), .o(n_905) );
in01f80 g568663 ( .a(x_out_1_2), .o(n_1611) );
in01f80 g568664 ( .a(x_out_9_4), .o(n_1688) );
in01f80 g568665 ( .a(x_out_35_20), .o(n_1220) );
in01f80 g568666 ( .a(x_out_44_14), .o(n_1350) );
in01f80 g568667 ( .a(x_out_53_5), .o(n_916) );
in01f80 g568668 ( .a(x_out_35_31), .o(n_997) );
in01f80 g568669 ( .a(x_out_18_26), .o(n_1862) );
in01f80 g568670 ( .a(x_out_40_9), .o(n_1004) );
in01f80 g568671 ( .a(x_out_26_3), .o(n_856) );
in01f80 g568672 ( .a(x_out_36_11), .o(n_409) );
in01f80 g568673 ( .a(x_out_9_14), .o(n_711) );
in01f80 g568674 ( .a(x_out_11_20), .o(n_438) );
in01f80 g568675 ( .a(x_out_31_8), .o(n_755) );
in01f80 g568676 ( .a(x_out_57_1), .o(n_209) );
in01f80 g568677 ( .a(x_out_10_19), .o(n_759) );
in01f80 g568678 ( .a(x_out_41_13), .o(n_1348) );
in01f80 g568679 ( .a(x_out_61_20), .o(n_1063) );
in01f80 g568680 ( .a(x_out_44_4), .o(n_1670) );
in01f80 g568681 ( .a(x_out_5_10), .o(n_584) );
in01f80 g568682 ( .a(x_out_9_0), .o(n_1900) );
in01f80 g568683 ( .a(x_out_30_32), .o(n_648) );
in01f80 g568684 ( .a(x_out_27_10), .o(n_1055) );
in01f80 g568685 ( .a(x_out_29_0), .o(n_1756) );
in01f80 g568686 ( .a(x_out_43_12), .o(n_804) );
in01f80 g568687 ( .a(x_out_27_1), .o(n_1349) );
in01f80 g568688 ( .a(x_out_25_22), .o(n_252) );
in01f80 g568689 ( .a(x_out_34_3), .o(n_927) );
in01f80 g568690 ( .a(x_out_3_32), .o(n_1099) );
in01f80 g568691 ( .a(x_out_32_10), .o(n_1937) );
in01f80 g568692 ( .a(x_out_27_24), .o(n_285) );
in01f80 g568693 ( .a(x_out_18_21), .o(n_1759) );
in01f80 g568694 ( .a(x_out_8_11), .o(n_1304) );
in01f80 g568695 ( .a(x_out_43_22), .o(n_854) );
in01f80 g568696 ( .a(x_out_6_9), .o(n_1696) );
in01f80 g568697 ( .a(x_out_19_0), .o(n_604) );
in01f80 g568698 ( .a(x_out_48_15), .o(n_1844) );
in01f80 g568699 ( .a(x_out_44_21), .o(n_157) );
in01f80 g568700 ( .a(x_out_5_24), .o(n_271) );
in01f80 g568701 ( .a(x_out_10_8), .o(n_134) );
in01f80 g568702 ( .a(x_out_27_23), .o(n_132) );
in01f80 g568703 ( .a(x_out_62_32), .o(n_595) );
in01f80 g568704 ( .a(x_out_14_26), .o(n_1339) );
in01f80 g568705 ( .a(x_out_39_21), .o(n_1933) );
in01f80 g568706 ( .a(x_out_40_3), .o(n_601) );
in01f80 g568707 ( .a(x_out_46_26), .o(n_248) );
in01f80 g568708 ( .a(x_out_30_25), .o(n_769) );
in01f80 g568709 ( .a(x_out_17_25), .o(n_1581) );
in01f80 g568710 ( .a(x_out_48_9), .o(n_413) );
in01f80 g568711 ( .a(x_out_40_29), .o(n_1602) );
in01f80 g568712 ( .a(x_out_4_2), .o(n_140) );
in01f80 g568713 ( .a(x_out_29_9), .o(n_589) );
in01f80 g568714 ( .a(x_out_24_27), .o(n_435) );
in01f80 g568715 ( .a(x_out_54_1), .o(n_623) );
in01f80 g568716 ( .a(x_out_2_4), .o(n_232) );
in01f80 g568717 ( .a(x_out_49_9), .o(n_1367) );
in01f80 g568718 ( .a(x_out_5_11), .o(n_235) );
in01f80 g568719 ( .a(x_out_13_2), .o(n_1456) );
in01f80 g568720 ( .a(x_out_48_5), .o(n_597) );
in01f80 g568721 ( .a(x_out_47_7), .o(n_189) );
in01f80 g568722 ( .a(x_out_44_24), .o(n_1804) );
in01f80 g568723 ( .a(x_out_33_18), .o(n_50) );
in01f80 g568724 ( .a(x_out_21_1), .o(n_524) );
in01f80 g568725 ( .a(x_out_8_10), .o(n_579) );
in01f80 g568726 ( .a(x_out_49_32), .o(n_428) );
in01f80 g568727 ( .a(x_out_2_2), .o(n_401) );
in01f80 g568728 ( .a(x_out_23_26), .o(n_1830) );
in01f80 g568729 ( .a(x_out_22_22), .o(n_1865) );
in01f80 g568730 ( .a(x_out_42_27), .o(n_1760) );
in01f80 g568731 ( .a(x_out_12_4), .o(n_652) );
in01f80 g568732 ( .a(x_out_30_2), .o(n_356) );
in01f80 g568733 ( .a(x_out_14_25), .o(n_852) );
in01f80 g568734 ( .a(x_out_13_9), .o(n_456) );
in01f80 g568735 ( .a(x_out_18_4), .o(n_1276) );
in01f80 g568736 ( .a(x_out_16_9), .o(n_113) );
in01f80 g568737 ( .a(x_out_30_5), .o(n_1294) );
in01f80 g568738 ( .a(x_out_57_26), .o(n_1561) );
in01f80 g568739 ( .a(x_out_60_32), .o(n_1575) );
in01f80 g568740 ( .a(x_out_10_4), .o(n_288) );
in01f80 g568741 ( .a(x_out_63_7), .o(n_1529) );
in01f80 g568742 ( .a(x_out_35_23), .o(n_1626) );
in01f80 g568743 ( .a(x_out_11_8), .o(n_395) );
in01f80 g568744 ( .a(x_out_47_15), .o(n_1103) );
in01f80 g568745 ( .a(x_out_49_29), .o(n_680) );
in01f80 g568746 ( .a(x_out_7_3), .o(n_1396) );
in01f80 g568747 ( .a(x_out_11_21), .o(n_28) );
in01f80 g568748 ( .a(x_out_6_22), .o(n_490) );
in01f80 g568749 ( .a(x_out_27_11), .o(n_1868) );
in01f80 g568750 ( .a(x_out_58_24), .o(n_740) );
in01f80 g568751 ( .a(x_out_39_29), .o(n_859) );
in01f80 g568752 ( .a(x_out_16_21), .o(n_64) );
in01f80 g568753 ( .a(x_out_24_23), .o(n_346) );
in01f80 g568754 ( .a(x_out_38_8), .o(n_1136) );
in01f80 g568755 ( .a(x_out_28_14), .o(n_129) );
in01f80 g568756 ( .a(x_out_12_8), .o(n_1112) );
in01f80 g568757 ( .a(x_out_59_22), .o(n_514) );
in01f80 g568758 ( .a(x_out_14_8), .o(n_398) );
in01f80 g568759 ( .a(x_out_31_22), .o(n_1460) );
in01f80 g568760 ( .a(x_out_33_25), .o(n_823) );
in01f80 g568761 ( .a(x_out_50_28), .o(n_1957) );
in01f80 g568762 ( .a(x_out_24_10), .o(n_625) );
in01f80 g568763 ( .a(x_out_24_26), .o(n_1034) );
in01f80 g568764 ( .a(x_out_17_2), .o(n_956) );
in01f80 g568765 ( .a(x_out_33_31), .o(n_1238) );
in01f80 g568766 ( .a(x_out_15_28), .o(n_1130) );
in01f80 g568767 ( .a(x_out_2_6), .o(n_292) );
in01f80 g568768 ( .a(x_out_13_19), .o(n_253) );
in01f80 g568769 ( .a(x_out_38_2), .o(n_1721) );
in01f80 g568770 ( .a(x_out_20_8), .o(n_166) );
in01f80 g568771 ( .a(x_out_27_18), .o(n_1812) );
in01f80 g568772 ( .a(x_out_11_12), .o(n_1552) );
in01f80 g568773 ( .a(x_out_57_22), .o(n_1380) );
in01f80 g568774 ( .a(x_out_9_11), .o(n_187) );
in01f80 g568775 ( .a(x_out_14_11), .o(n_530) );
in01f80 g568776 ( .a(x_out_62_24), .o(n_1681) );
in01f80 g568777 ( .a(x_out_16_5), .o(n_1190) );
in01f80 g568778 ( .a(x_out_34_23), .o(n_1110) );
in01f80 g568779 ( .a(x_out_38_7), .o(n_54) );
in01f80 g568780 ( .a(x_out_51_1), .o(n_1195) );
in01f80 g568781 ( .a(x_out_28_2), .o(n_863) );
in01f80 g568782 ( .a(x_out_19_11), .o(n_385) );
in01f80 g568783 ( .a(x_out_18_29), .o(n_1425) );
in01f80 g568784 ( .a(x_out_16_30), .o(n_1819) );
in01f80 g568785 ( .a(x_out_56_28), .o(n_1601) );
in01f80 g568786 ( .a(x_out_5_9), .o(n_5) );
in01f80 g568787 ( .a(x_out_10_10), .o(n_213) );
in01f80 g568788 ( .a(x_out_31_29), .o(n_35) );
in01f80 g568789 ( .a(x_out_4_3), .o(n_122) );
in01f80 g568790 ( .a(x_out_27_7), .o(n_1419) );
in01f80 g568791 ( .a(x_out_24_5), .o(n_862) );
in01f80 g568792 ( .a(x_out_53_12), .o(n_1906) );
in01f80 g568793 ( .a(x_out_14_6), .o(n_1434) );
in01f80 g568794 ( .a(x_out_37_23), .o(n_1615) );
in01f80 g568795 ( .a(x_out_41_4), .o(n_90) );
in01f80 g568796 ( .a(x_out_11_9), .o(n_1644) );
in01f80 g568797 ( .a(x_out_62_20), .o(n_1076) );
in01f80 g568798 ( .a(x_out_18_2), .o(n_673) );
in01f80 g568799 ( .a(x_out_3_21), .o(n_386) );
in01f80 g568800 ( .a(x_out_6_13), .o(n_1956) );
in01f80 g568801 ( .a(x_out_22_25), .o(n_768) );
in01f80 g568802 ( .a(x_out_34_30), .o(n_1084) );
in01f80 g568803 ( .a(x_out_42_12), .o(n_1312) );
in01f80 g568804 ( .a(x_out_58_0), .o(n_382) );
in01f80 g568805 ( .a(x_out_54_9), .o(n_1139) );
in01f80 g568806 ( .a(x_out_24_1), .o(n_211) );
in01f80 g568807 ( .a(x_out_53_8), .o(n_1142) );
in01f80 g568808 ( .a(x_out_61_0), .o(n_1572) );
in01f80 g568809 ( .a(x_out_10_5), .o(n_1743) );
in01f80 g568810 ( .a(x_out_2_21), .o(n_1639) );
in01f80 g568811 ( .a(x_out_32_12), .o(n_518) );
in01f80 g568812 ( .a(x_out_10_9), .o(n_570) );
in01f80 g568813 ( .a(x_out_13_29), .o(n_1166) );
in01f80 g568814 ( .a(x_out_19_29), .o(n_935) );
in01f80 g568815 ( .a(x_out_22_26), .o(n_1711) );
in01f80 g568816 ( .a(x_out_16_2), .o(n_1414) );
in01f80 g568817 ( .a(x_out_45_4), .o(n_1442) );
in01f80 g568818 ( .a(x_out_27_25), .o(n_1101) );
in01f80 g568819 ( .a(x_out_3_14), .o(n_277) );
in01f80 g568820 ( .a(x_out_29_31), .o(n_1344) );
in01f80 g568821 ( .a(x_out_43_3), .o(n_1001) );
in01f80 g568822 ( .a(x_out_40_15), .o(n_746) );
in01f80 g568823 ( .a(x_out_52_1), .o(n_1715) );
in01f80 g568824 ( .a(x_out_51_20), .o(n_1643) );
in01f80 g568825 ( .a(x_out_51_26), .o(n_1054) );
in01f80 g568826 ( .a(x_out_61_12), .o(n_1239) );
in01f80 g568827 ( .a(x_out_63_33), .o(n_1065) );
in01f80 g568828 ( .a(x_out_37_10), .o(n_1429) );
in01f80 g568829 ( .a(x_out_6_31), .o(n_611) );
in01f80 g568830 ( .a(x_out_13_24), .o(n_359) );
in01f80 g568831 ( .a(x_out_61_5), .o(n_326) );
in01f80 g568832 ( .a(x_out_42_8), .o(n_1763) );
in01f80 g568833 ( .a(x_out_4_15), .o(n_553) );
in01f80 g568834 ( .a(x_out_25_5), .o(n_1373) );
in01f80 g568835 ( .a(x_out_7_31), .o(n_476) );
in01f80 g568836 ( .a(x_out_25_33), .o(n_1418) );
in01f80 g568837 ( .a(x_out_14_14), .o(n_93) );
in01f80 g568838 ( .a(x_out_44_31), .o(n_453) );
in01f80 g568839 ( .a(x_out_37_9), .o(n_311) );
in01f80 g568840 ( .a(x_out_1_23), .o(n_590) );
in01f80 g568841 ( .a(x_out_20_1), .o(n_688) );
in01f80 g568842 ( .a(x_out_11_14), .o(n_47) );
in01f80 g568843 ( .a(x_out_16_6), .o(n_522) );
in01f80 g568844 ( .a(x_out_26_4), .o(n_334) );
in01f80 g568845 ( .a(x_out_36_2), .o(n_848) );
in01f80 g568846 ( .a(x_out_36_15), .o(n_1391) );
in01f80 g568847 ( .a(x_out_51_25), .o(n_1198) );
in01f80 g568848 ( .a(x_out_58_13), .o(n_1320) );
in01f80 g568849 ( .a(x_out_50_25), .o(n_774) );
in01f80 g568850 ( .a(x_out_17_4), .o(n_156) );
in01f80 g568851 ( .a(x_out_38_29), .o(n_1975) );
in01f80 g568852 ( .a(x_out_3_19), .o(n_13) );
in01f80 g568853 ( .a(x_out_9_10), .o(n_445) );
in01f80 g568854 ( .a(x_out_35_18), .o(n_780) );
in01f80 g568855 ( .a(x_out_22_6), .o(n_1007) );
in01f80 g568856 ( .a(x_out_40_0), .o(n_868) );
in01f80 g568857 ( .a(x_out_5_21), .o(n_337) );
in01f80 g568858 ( .a(x_out_12_7), .o(n_1710) );
in01f80 g568859 ( .a(x_out_59_4), .o(n_94) );
in01f80 g568860 ( .a(x_out_59_11), .o(n_186) );
in01f80 g568861 ( .a(x_out_37_31), .o(n_1050) );
in01f80 g568862 ( .a(x_out_21_22), .o(n_1196) );
in01f80 g568863 ( .a(x_out_40_20), .o(n_943) );
in01f80 g568864 ( .a(x_out_60_10), .o(n_154) );
in01f80 g568865 ( .a(x_out_30_28), .o(n_178) );
in01f80 g568866 ( .a(x_out_1_19), .o(n_1969) );
in01f80 g568867 ( .a(x_out_39_11), .o(n_434) );
in01f80 g568868 ( .a(x_out_45_29), .o(n_607) );
in01f80 g568869 ( .a(x_out_59_27), .o(n_1807) );
in01f80 g568870 ( .a(x_out_3_30), .o(n_684) );
in01f80 g568871 ( .a(x_out_8_1), .o(n_181) );
in01f80 g568872 ( .a(x_out_29_14), .o(n_701) );
in01f80 g568873 ( .a(x_out_28_33), .o(n_360) );
in01f80 g568874 ( .a(x_out_29_30), .o(n_1233) );
in01f80 g568875 ( .a(x_out_58_28), .o(n_1355) );
in01f80 g568876 ( .a(x_out_8_27), .o(n_1405) );
in01f80 g568877 ( .a(x_out_1_22), .o(n_1141) );
in01f80 g568878 ( .a(x_out_17_23), .o(n_886) );
in01f80 g568879 ( .a(x_out_2_15), .o(n_1746) );
in01f80 g568880 ( .a(x_out_34_20), .o(n_254) );
in01f80 g568881 ( .a(x_out_18_9), .o(n_1664) );
in01f80 g568882 ( .a(x_out_36_10), .o(n_1131) );
in01f80 g568883 ( .a(x_out_41_9), .o(n_84) );
in01f80 g568884 ( .a(x_out_39_5), .o(n_1635) );
in01f80 g568885 ( .a(x_out_34_8), .o(n_1453) );
in01f80 g568886 ( .a(x_out_36_29), .o(n_1098) );
in01f80 g568887 ( .a(x_out_41_22), .o(n_940) );
in01f80 g568888 ( .a(x_out_39_10), .o(n_328) );
in01f80 g568889 ( .a(x_out_6_28), .o(n_473) );
in01f80 g568890 ( .a(x_out_14_15), .o(n_1598) );
in01f80 g568891 ( .a(x_out_54_27), .o(n_1346) );
in01f80 g568892 ( .a(x_out_3_12), .o(n_531) );
in01f80 g568893 ( .a(x_out_31_7), .o(n_1573) );
in01f80 g568894 ( .a(x_out_56_26), .o(n_1128) );
in01f80 g568895 ( .a(x_out_46_6), .o(n_1686) );
in01f80 g568896 ( .a(x_out_13_20), .o(n_299) );
in01f80 g568897 ( .a(x_out_15_1), .o(n_1958) );
in01f80 g568898 ( .a(x_out_41_28), .o(n_549) );
in01f80 g568899 ( .a(x_out_10_3), .o(n_1245) );
in01f80 g568900 ( .a(x_out_44_0), .o(n_678) );
in01f80 g568901 ( .a(x_out_7_21), .o(n_1737) );
in01f80 g568902 ( .a(x_out_9_3), .o(n_212) );
in01f80 g568903 ( .a(x_out_25_21), .o(n_1234) );
in01f80 g568904 ( .a(x_out_50_3), .o(n_1765) );
in01f80 g568905 ( .a(x_out_36_30), .o(n_795) );
in01f80 g568906 ( .a(x_out_18_23), .o(n_1904) );
in01f80 g568907 ( .a(x_out_27_9), .o(n_782) );
in01f80 g568908 ( .a(x_out_36_24), .o(n_1802) );
in01f80 g568909 ( .a(x_out_10_6), .o(n_1403) );
in01f80 g568910 ( .a(x_out_54_26), .o(n_1774) );
in01f80 g568911 ( .a(x_out_16_24), .o(n_183) );
in01f80 g568912 ( .a(x_out_42_30), .o(n_81) );
in01f80 g568913 ( .a(x_out_26_20), .o(n_980) );
in01f80 g568914 ( .a(x_out_8_31), .o(n_1347) );
in01f80 g568915 ( .a(x_out_44_28), .o(n_1096) );
in01f80 g568916 ( .a(x_out_42_10), .o(n_1313) );
in01f80 g568917 ( .a(x_out_33_1), .o(n_294) );
in01f80 g568918 ( .a(x_out_2_18), .o(n_778) );
in01f80 g568919 ( .a(x_out_2_1), .o(n_919) );
in01f80 g568920 ( .a(x_out_15_24), .o(n_1452) );
in01f80 g568921 ( .a(x_out_42_20), .o(n_1027) );
in01f80 g568922 ( .a(x_out_39_12), .o(n_1540) );
in01f80 g568923 ( .a(x_out_3_29), .o(n_1221) );
in01f80 g568924 ( .a(x_out_42_1), .o(n_1123) );
in01f80 g568925 ( .a(x_out_21_30), .o(n_1169) );
in01f80 g568926 ( .a(x_out_1_0), .o(n_988) );
in01f80 g568927 ( .a(x_out_33_27), .o(n_1882) );
in01f80 g568928 ( .a(x_out_46_23), .o(n_1784) );
in01f80 g568929 ( .a(x_out_51_12), .o(n_662) );
in01f80 g568930 ( .a(x_out_55_11), .o(n_1864) );
in01f80 g568931 ( .a(x_out_3_8), .o(n_1824) );
in01f80 g568932 ( .a(x_out_62_14), .o(n_1230) );
in01f80 g568933 ( .a(x_out_11_5), .o(n_515) );
in01f80 g568934 ( .a(x_out_40_14), .o(n_1095) );
in01f80 g568935 ( .a(x_out_2_23), .o(n_6) );
in01f80 g568936 ( .a(x_out_4_14), .o(n_1667) );
in01f80 g568937 ( .a(x_out_22_11), .o(n_121) );
in01f80 g568938 ( .a(x_out_2_3), .o(n_1473) );
in01f80 g568939 ( .a(x_out_5_33), .o(n_1836) );
in01f80 g568940 ( .a(x_out_39_2), .o(n_377) );
in01f80 g568941 ( .a(x_out_15_0), .o(n_1520) );
in01f80 g568942 ( .a(x_out_53_10), .o(n_284) );
in01f80 g568943 ( .a(x_out_11_19), .o(n_996) );
in01f80 g568944 ( .a(x_out_28_11), .o(n_1672) );
in01f80 g568945 ( .a(x_out_16_31), .o(n_402) );
in01f80 g568946 ( .a(x_out_26_19), .o(n_1921) );
in01f80 g568947 ( .a(x_out_24_18), .o(n_494) );
in01f80 g568948 ( .a(x_out_6_0), .o(n_1753) );
in01f80 g568949 ( .a(x_out_54_15), .o(n_14) );
in01f80 g568950 ( .a(x_out_6_3), .o(n_840) );
in01f80 g568951 ( .a(x_out_13_22), .o(n_1032) );
in01f80 g568952 ( .a(x_out_59_0), .o(n_349) );
in01f80 g568953 ( .a(x_out_22_33), .o(n_222) );
in01f80 g568954 ( .a(x_out_24_33), .o(n_918) );
in01f80 g568955 ( .a(x_out_35_5), .o(n_25) );
in01f80 g568956 ( .a(x_out_27_0), .o(n_1124) );
in01f80 g568957 ( .a(x_out_7_20), .o(n_550) );
in01f80 g568958 ( .a(x_out_16_23), .o(n_890) );
in01f80 g568959 ( .a(x_out_19_5), .o(n_896) );
in01f80 g568960 ( .a(x_out_56_13), .o(n_1444) );
in01f80 g568961 ( .a(x_out_44_18), .o(n_180) );
in01f80 g568962 ( .a(x_out_58_29), .o(n_592) );
in01f80 g568963 ( .a(x_out_54_24), .o(n_1135) );
in01f80 g568964 ( .a(x_out_23_28), .o(n_816) );
in01f80 g568965 ( .a(x_out_31_13), .o(n_1588) );
in01f80 g568966 ( .a(x_out_6_21), .o(n_1323) );
in01f80 g568967 ( .a(x_out_0_7), .o(n_1060) );
in01f80 g568968 ( .a(x_out_53_22), .o(n_315) );
in01f80 g568969 ( .a(x_out_17_20), .o(n_865) );
in01f80 g568970 ( .a(x_out_35_26), .o(n_725) );
in01f80 g568971 ( .a(x_out_62_3), .o(n_1878) );
in01f80 g568972 ( .a(x_out_18_31), .o(n_1343) );
in01f80 g568973 ( .a(x_out_1_28), .o(n_1324) );
in01f80 g568974 ( .a(x_out_34_7), .o(n_1493) );
in01f80 g568975 ( .a(x_out_55_8), .o(n_665) );
in01f80 g568976 ( .a(x_out_27_19), .o(n_1809) );
in01f80 g568977 ( .a(x_out_59_2), .o(n_1407) );
in01f80 g568978 ( .a(x_out_47_20), .o(n_1789) );
in01f80 g568979 ( .a(x_out_57_2), .o(n_821) );
in01f80 g568980 ( .a(x_out_48_24), .o(n_1881) );
in01f80 g568981 ( .a(x_out_60_20), .o(n_1057) );
in01f80 g568982 ( .a(x_out_45_14), .o(n_449) );
in01f80 g568983 ( .a(x_out_43_14), .o(n_1950) );
in01f80 g568984 ( .a(x_out_10_13), .o(n_426) );
in01f80 g568985 ( .a(x_out_55_31), .o(n_1261) );
in01f80 g568986 ( .a(x_out_11_30), .o(n_1399) );
in01f80 g568987 ( .a(x_out_39_22), .o(n_1314) );
in01f80 g568988 ( .a(x_out_59_3), .o(n_794) );
in01f80 g568989 ( .a(x_out_1_20), .o(n_1146) );
in01f80 g568990 ( .a(x_out_47_26), .o(n_1464) );
in01f80 g568991 ( .a(x_out_34_6), .o(n_1184) );
in01f80 g568992 ( .a(x_out_6_19), .o(n_971) );
in01f80 g568993 ( .a(x_out_44_10), .o(n_998) );
in01f80 g568994 ( .a(x_out_56_19), .o(n_1570) );
in01f80 g568995 ( .a(x_out_4_26), .o(n_1302) );
in01f80 g568996 ( .a(x_out_1_31), .o(n_124) );
in01f80 g568997 ( .a(x_out_41_7), .o(n_544) );
in01f80 g568998 ( .a(x_out_19_33), .o(n_440) );
in01f80 g568999 ( .a(x_out_31_33), .o(n_135) );
in01f80 g569000 ( .a(x_out_43_21), .o(n_802) );
in01f80 g569001 ( .a(x_out_16_20), .o(n_374) );
in01f80 g569002 ( .a(x_out_51_11), .o(n_10) );
in01f80 g569003 ( .a(x_out_7_12), .o(n_458) );
in01f80 g569004 ( .a(x_out_30_33), .o(n_709) );
in01f80 g569005 ( .a(x_out_15_31), .o(n_1800) );
in01f80 g569006 ( .a(x_out_7_9), .o(n_1270) );
in01f80 g569007 ( .a(x_out_24_20), .o(n_388) );
in01f80 g569008 ( .a(x_out_2_19), .o(n_1895) );
in01f80 g569009 ( .a(x_out_29_15), .o(n_55) );
in01f80 g569010 ( .a(x_out_41_0), .o(n_1558) );
in01f80 g569011 ( .a(x_out_9_2), .o(n_1290) );
in01f80 g569012 ( .a(x_out_42_18), .o(n_206) );
in01f80 g569013 ( .a(x_out_34_1), .o(n_9) );
in01f80 g569014 ( .a(x_out_27_21), .o(n_1120) );
in01f80 g569015 ( .a(x_out_61_4), .o(n_1668) );
in01f80 g569016 ( .a(x_out_40_22), .o(n_454) );
in01f80 g569017 ( .a(x_out_21_8), .o(n_11) );
in01f80 g569018 ( .a(x_out_32_4), .o(n_150) );
in01f80 g569019 ( .a(x_out_31_28), .o(n_1597) );
in01f80 g569020 ( .a(x_out_13_1), .o(n_879) );
in01f80 g569021 ( .a(x_out_25_31), .o(n_1042) );
in01f80 g569022 ( .a(x_out_59_9), .o(n_1936) );
in01f80 g569023 ( .a(x_out_35_14), .o(n_793) );
in01f80 g569024 ( .a(x_out_39_23), .o(n_1524) );
in01f80 g569025 ( .a(x_out_55_29), .o(n_1462) );
in01f80 g569026 ( .a(x_out_17_8), .o(n_1211) );
in01f80 g569027 ( .a(x_out_62_18), .o(n_171) );
in01f80 g569028 ( .a(x_out_33_28), .o(n_1237) );
in01f80 g569029 ( .a(x_out_19_12), .o(n_1871) );
in01f80 g569030 ( .a(x_out_50_13), .o(n_203) );
in01f80 g569031 ( .a(x_out_7_19), .o(n_1770) );
in01f80 g569032 ( .a(x_out_41_26), .o(n_955) );
in01f80 g569033 ( .a(x_out_33_32), .o(n_1736) );
in01f80 g569034 ( .a(x_out_36_21), .o(n_160) );
in01f80 g569035 ( .a(x_out_45_30), .o(n_1052) );
in01f80 g569036 ( .a(x_out_14_10), .o(n_1962) );
in01f80 g569037 ( .a(x_out_29_7), .o(n_565) );
in01f80 g569038 ( .a(x_out_16_4), .o(n_144) );
in01f80 g569039 ( .a(x_out_51_14), .o(n_909) );
in01f80 g569040 ( .a(x_out_59_32), .o(n_422) );
in01f80 g569041 ( .a(x_out_51_28), .o(n_806) );
in01f80 g569042 ( .a(x_out_61_10), .o(n_46) );
in01f80 g569043 ( .a(x_out_20_11), .o(n_543) );
in01f80 g569044 ( .a(x_out_63_15), .o(n_835) );
in01f80 g569045 ( .a(x_out_52_3), .o(n_1177) );
in01f80 g569046 ( .a(x_out_28_25), .o(n_575) );
in01f80 g569047 ( .a(x_out_56_5), .o(n_1879) );
in01f80 g569048 ( .a(x_out_59_8), .o(n_1701) );
in01f80 g569049 ( .a(x_out_53_13), .o(n_460) );
in01f80 g569050 ( .a(x_out_28_6), .o(n_357) );
in01f80 g569051 ( .a(x_out_49_1), .o(n_1397) );
in01f80 g569052 ( .a(x_out_56_10), .o(n_649) );
in01f80 g569053 ( .a(x_out_23_6), .o(n_1853) );
in01f80 g569054 ( .a(x_out_7_2), .o(n_1301) );
in01f80 g569055 ( .a(x_out_12_19), .o(n_682) );
in01f80 g569056 ( .a(x_out_36_28), .o(n_908) );
in01f80 g569057 ( .a(x_out_53_11), .o(n_876) );
in01f80 g569058 ( .a(x_out_63_13), .o(n_686) );
in01f80 g569059 ( .a(x_out_60_27), .o(n_1143) );
in01f80 g569060 ( .a(x_out_11_6), .o(n_1443) );
in01f80 g569061 ( .a(x_out_61_24), .o(n_846) );
in01f80 g569062 ( .a(x_out_10_33), .o(n_681) );
in01f80 g569063 ( .a(x_out_56_24), .o(n_1006) );
in01f80 g569064 ( .a(x_out_23_8), .o(n_671) );
in01f80 g569065 ( .a(x_out_37_7), .o(n_632) );
in01f80 g569066 ( .a(x_out_11_29), .o(n_691) );
in01f80 g569067 ( .a(x_out_30_11), .o(n_700) );
in01f80 g569068 ( .a(x_out_37_15), .o(n_429) );
in01f80 g569069 ( .a(x_out_37_18), .o(n_669) );
in01f80 g569070 ( .a(x_out_55_2), .o(n_352) );
in01f80 g569071 ( .a(x_out_6_12), .o(n_1754) );
in01f80 g569072 ( .a(x_out_24_19), .o(n_468) );
in01f80 g569073 ( .a(x_out_23_20), .o(n_641) );
in01f80 g569074 ( .a(x_out_43_15), .o(n_74) );
in01f80 g569075 ( .a(x_out_33_7), .o(n_1227) );
in01f80 g569076 ( .a(x_out_18_33), .o(n_775) );
in01f80 g569077 ( .a(x_out_57_10), .o(n_1408) );
in01f80 g569078 ( .a(x_out_18_3), .o(n_420) );
in01f80 g569079 ( .a(x_out_17_24), .o(n_1748) );
in01f80 g569080 ( .a(x_out_24_28), .o(n_0) );
in01f80 g569081 ( .a(x_out_28_20), .o(n_410) );
in01f80 g569082 ( .a(x_out_51_5), .o(n_333) );
in01f80 g569083 ( .a(x_out_30_1), .o(n_517) );
in01f80 g569084 ( .a(x_out_48_3), .o(n_1897) );
in01f80 g569085 ( .a(x_out_5_6), .o(n_362) );
in01f80 g569086 ( .a(x_out_34_21), .o(n_1740) );
in01f80 g569087 ( .a(x_out_8_32), .o(n_256) );
in01f80 g569088 ( .a(x_out_16_26), .o(n_1068) );
in01f80 g569089 ( .a(x_out_10_2), .o(n_1555) );
in01f80 g569090 ( .a(x_out_13_31), .o(n_1104) );
in01f80 g569091 ( .a(x_out_0_3), .o(n_1960) );
in01f80 g569092 ( .a(x_out_4_0), .o(n_425) );
in01f80 g569093 ( .a(x_out_37_8), .o(n_1842) );
in01f80 g569094 ( .a(x_out_22_31), .o(n_484) );
in01f80 g569095 ( .a(x_out_30_6), .o(n_1235) );
in01f80 g569096 ( .a(x_out_14_21), .o(n_1149) );
in01f80 g569097 ( .a(x_out_57_9), .o(n_1803) );
in01f80 g569098 ( .a(x_out_21_23), .o(n_627) );
in01f80 g569099 ( .a(x_out_5_12), .o(n_169) );
in01f80 g569100 ( .a(x_out_59_5), .o(n_1409) );
in01f80 g569101 ( .a(x_out_52_11), .o(n_1377) );
in01f80 g569102 ( .a(x_out_22_9), .o(n_1583) );
in01f80 g569103 ( .a(x_out_12_14), .o(n_1875) );
in01f80 g569104 ( .a(x_out_23_19), .o(n_225) );
in01f80 g569105 ( .a(x_out_48_30), .o(n_1716) );
in01f80 g569106 ( .a(x_out_20_6), .o(n_1620) );
in01f80 g569107 ( .a(x_out_32_2), .o(n_1673) );
in01f80 g569108 ( .a(x_out_52_9), .o(n_600) );
in01f80 g569109 ( .a(x_out_7_15), .o(n_265) );
in01f80 g569110 ( .a(x_out_8_2), .o(n_1318) );
in01f80 g569111 ( .a(x_out_40_2), .o(n_1679) );
in01f80 g569112 ( .a(x_out_46_10), .o(n_1846) );
in01f80 g569113 ( .a(x_out_17_22), .o(n_1941) );
in01f80 g569114 ( .a(x_out_30_3), .o(n_43) );
in01f80 g569115 ( .a(x_out_28_18), .o(n_471) );
in01f80 g569116 ( .a(x_out_46_28), .o(n_158) );
in01f80 g569117 ( .a(x_out_30_9), .o(n_430) );
in01f80 g569118 ( .a(x_out_10_26), .o(n_557) );
in01f80 g569119 ( .a(x_out_1_24), .o(n_1012) );
in01f80 g569120 ( .a(x_out_31_20), .o(n_520) );
in01f80 g569121 ( .a(x_out_16_3), .o(n_1264) );
in01f80 g569122 ( .a(x_out_8_22), .o(n_1883) );
in01f80 g569123 ( .a(x_out_44_1), .o(n_888) );
in01f80 g569124 ( .a(x_out_20_5), .o(n_1148) );
in01f80 g569125 ( .a(x_out_26_32), .o(n_1422) );
in01f80 g569126 ( .a(x_out_36_3), .o(n_1438) );
in01f80 g569127 ( .a(x_out_23_25), .o(n_1762) );
in01f80 g569128 ( .a(x_out_30_4), .o(n_1258) );
in01f80 g569129 ( .a(x_out_39_25), .o(n_49) );
in01f80 g569130 ( .a(x_out_59_1), .o(n_1607) );
in01f80 g569131 ( .a(x_out_19_1), .o(n_1206) );
in01f80 g569132 ( .a(x_out_2_25), .o(n_788) );
in01f80 g569133 ( .a(x_out_26_11), .o(n_290) );
in01f80 g569134 ( .a(x_out_3_25), .o(n_1779) );
in01f80 g569135 ( .a(x_out_23_15), .o(n_1470) );
in01f80 g569136 ( .a(x_out_8_15), .o(n_1400) );
in01f80 g569137 ( .a(x_out_49_23), .o(n_1287) );
in01f80 g569138 ( .a(x_out_2_9), .o(n_1486) );
in01f80 g569139 ( .a(x_out_58_12), .o(n_1690) );
in01f80 g569140 ( .a(x_out_60_24), .o(n_1666) );
in01f80 g569141 ( .a(x_out_11_0), .o(n_1441) );
in01f80 g569142 ( .a(x_out_61_11), .o(n_500) );
in01f80 g569143 ( .a(x_out_40_8), .o(n_1959) );
in01f80 g569144 ( .a(x_out_41_33), .o(n_1454) );
in01f80 g569145 ( .a(x_out_12_29), .o(n_526) );
in01f80 g569146 ( .a(x_out_35_8), .o(n_1106) );
in01f80 g569147 ( .a(x_out_29_8), .o(n_1531) );
in01f80 g569148 ( .a(x_out_51_23), .o(n_1307) );
in01f80 g569149 ( .a(x_out_28_23), .o(n_102) );
in01f80 g569150 ( .a(x_out_48_21), .o(n_883) );
in01f80 g569151 ( .a(x_out_13_11), .o(n_551) );
in01f80 g569152 ( .a(x_out_6_2), .o(n_797) );
in01f80 g569153 ( .a(x_out_38_24), .o(n_729) );
in01f80 g569154 ( .a(x_out_34_10), .o(n_608) );
in01f80 g569155 ( .a(x_out_12_6), .o(n_1559) );
in01f80 g569156 ( .a(x_out_36_4), .o(n_523) );
in01f80 g569157 ( .a(x_out_19_19), .o(n_976) );
in01f80 g569158 ( .a(x_out_63_10), .o(n_1860) );
in01f80 g569159 ( .a(x_out_9_27), .o(n_493) );
in01f80 g569160 ( .a(x_out_9_9), .o(n_38) );
in01f80 g569161 ( .a(x_out_49_15), .o(n_588) );
in01f80 g569162 ( .a(x_out_56_29), .o(n_318) );
in01f80 g569163 ( .a(x_out_33_12), .o(n_1333) );
in01f80 g569164 ( .a(x_out_3_22), .o(n_1514) );
in01f80 g569165 ( .a(x_out_52_14), .o(n_880) );
in01f80 g569166 ( .a(x_out_26_0), .o(n_108) );
in01f80 g569167 ( .a(x_out_46_22), .o(n_1646) );
in01f80 g569168 ( .a(x_out_44_23), .o(n_1909) );
in01f80 g569169 ( .a(x_out_31_9), .o(n_639) );
in01f80 g569170 ( .a(x_out_47_5), .o(n_1530) );
in01f80 g569171 ( .a(x_out_45_12), .o(n_1628) );
in01f80 g569172 ( .a(x_out_27_15), .o(n_1775) );
in01f80 g569173 ( .a(x_out_57_6), .o(n_312) );
in01f80 g569174 ( .a(x_out_63_1), .o(n_379) );
in01f80 g569175 ( .a(x_out_58_9), .o(n_537) );
in01f80 g569176 ( .a(x_out_8_18), .o(n_1248) );
in01f80 g569177 ( .a(x_out_54_0), .o(n_387) );
in01f80 g569178 ( .a(x_out_2_24), .o(n_1011) );
in01f80 g569179 ( .a(x_out_1_25), .o(n_406) );
in01f80 g569180 ( .a(x_out_6_4), .o(n_683) );
in01f80 g569181 ( .a(x_out_7_11), .o(n_16) );
in01f80 g569182 ( .a(x_out_9_19), .o(n_378) );
in01f80 g569183 ( .a(x_out_10_25), .o(n_1718) );
in01f80 g569184 ( .a(x_out_11_23), .o(n_1179) );
in01f80 g569185 ( .a(x_out_17_31), .o(n_44) );
in01f80 g569186 ( .a(x_out_9_5), .o(n_495) );
in01f80 g569187 ( .a(x_out_24_29), .o(n_12) );
in01f80 g569188 ( .a(x_out_2_14), .o(n_1772) );
in01f80 g569189 ( .a(x_out_37_20), .o(n_439) );
in01f80 g569190 ( .a(x_out_40_5), .o(n_964) );
in01f80 g569191 ( .a(x_out_41_5), .o(n_1578) );
in01f80 g569192 ( .a(x_out_3_24), .o(n_1659) );
in01f80 g569193 ( .a(x_out_57_33), .o(n_1791) );
in01f80 g569194 ( .a(x_out_21_19), .o(n_1548) );
in01f80 g569195 ( .a(x_out_18_32), .o(n_944) );
in01f80 g569196 ( .a(x_out_36_6), .o(n_945) );
in01f80 g569197 ( .a(x_out_36_32), .o(n_847) );
in01f80 g569198 ( .a(x_out_21_25), .o(n_538) );
in01f80 g569199 ( .a(x_out_36_20), .o(n_85) );
in01f80 g569200 ( .a(x_out_21_21), .o(n_1247) );
in01f80 g569201 ( .a(x_out_19_20), .o(n_982) );
in01f80 g569202 ( .a(x_out_63_2), .o(n_1855) );
in01f80 g569203 ( .a(x_out_28_3), .o(n_1109) );
in01f80 g569204 ( .a(x_out_10_14), .o(n_65) );
in01f80 g569205 ( .a(x_out_14_30), .o(n_1088) );
in01f80 g569206 ( .a(x_out_53_1), .o(n_787) );
in01f80 g569207 ( .a(x_out_5_23), .o(n_798) );
in01f80 g569208 ( .a(x_out_31_23), .o(n_1663) );
in01f80 g569209 ( .a(x_out_18_11), .o(n_1510) );
in01f80 g569210 ( .a(x_out_55_10), .o(n_1731) );
in01f80 g569211 ( .a(x_out_63_12), .o(n_651) );
in01f80 g569212 ( .a(x_out_4_29), .o(n_1833) );
in01f80 g569213 ( .a(x_out_44_7), .o(n_1927) );
in01f80 g569214 ( .a(x_out_15_22), .o(n_262) );
in01f80 g569215 ( .a(x_out_56_7), .o(n_1606) );
in01f80 g569216 ( .a(x_out_50_11), .o(n_427) );
in01f80 g569217 ( .a(x_out_36_33), .o(n_1311) );
in01f80 g569218 ( .a(x_out_20_9), .o(n_1940) );
in01f80 g569219 ( .a(x_out_25_8), .o(n_1692) );
in01f80 g569220 ( .a(x_out_10_22), .o(n_1303) );
in01f80 g569221 ( .a(x_out_28_32), .o(n_1378) );
in01f80 g569222 ( .a(x_out_56_15), .o(n_1817) );
in01f80 g569223 ( .a(x_out_42_28), .o(n_585) );
in01f80 g569224 ( .a(x_out_45_13), .o(n_371) );
in01f80 g569225 ( .a(x_out_26_21), .o(n_120) );
in01f80 g569226 ( .a(x_out_41_31), .o(n_1357) );
in01f80 g569227 ( .a(x_out_14_32), .o(n_1949) );
in01f80 g569228 ( .a(x_out_31_24), .o(n_1108) );
in01f80 g569229 ( .a(x_out_35_27), .o(n_643) );
in01f80 g569230 ( .a(x_out_45_1), .o(n_763) );
in01f80 g569231 ( .a(x_out_43_9), .o(n_66) );
in01f80 g569232 ( .a(x_out_18_24), .o(n_1209) );
in01f80 g569233 ( .a(x_out_12_27), .o(n_1033) );
in01f80 g569234 ( .a(x_out_47_0), .o(n_174) );
in01f80 g569235 ( .a(x_out_4_27), .o(n_201) );
in01f80 g569236 ( .a(x_out_2_5), .o(n_912) );
in01f80 g569237 ( .a(x_out_59_19), .o(n_761) );
in01f80 g569238 ( .a(x_out_3_4), .o(n_1798) );
in01f80 g569239 ( .a(x_out_33_2), .o(n_644) );
in01f80 g569240 ( .a(x_out_8_30), .o(n_396) );
in01f80 g569241 ( .a(x_out_60_0), .o(n_1856) );
in01f80 g569242 ( .a(x_out_53_15), .o(n_1815) );
in01f80 g569243 ( .a(x_out_5_18), .o(n_1293) );
in01f80 g569244 ( .a(x_out_43_28), .o(n_723) );
in01f80 g569245 ( .a(x_out_44_25), .o(n_1038) );
in01f80 g569246 ( .a(x_out_44_3), .o(n_1706) );
in01f80 g569247 ( .a(x_out_9_8), .o(n_1345) );
in01f80 g569248 ( .a(x_out_47_13), .o(n_1867) );
in01f80 g569249 ( .a(x_out_4_21), .o(n_236) );
in01f80 g569250 ( .a(x_out_23_23), .o(n_528) );
in01f80 g569251 ( .a(x_out_37_29), .o(n_1271) );
in01f80 g569252 ( .a(x_out_24_13), .o(n_1951) );
in01f80 g569253 ( .a(x_out_33_22), .o(n_234) );
in01f80 g569254 ( .a(x_out_24_3), .o(n_1172) );
in01f80 g569255 ( .a(x_out_43_26), .o(n_1537) );
in01f80 g569256 ( .a(x_out_19_30), .o(n_1816) );
in01f80 g569257 ( .a(x_out_1_12), .o(n_329) );
in01f80 g569258 ( .a(x_out_32_14), .o(n_993) );
in01f80 g569259 ( .a(x_out_31_32), .o(n_1684) );
in01f80 g569260 ( .a(x_out_16_22), .o(n_706) );
in01f80 g569261 ( .a(x_out_5_5), .o(n_614) );
in01f80 g569262 ( .a(x_out_45_6), .o(n_73) );
in01f80 g569263 ( .a(x_out_2_29), .o(n_403) );
in01f80 g569264 ( .a(x_out_49_8), .o(n_781) );
in01f80 g569265 ( .a(x_out_22_28), .o(n_1780) );
in01f80 g569266 ( .a(x_out_45_0), .o(n_578) );
in01f80 g569267 ( .a(x_out_39_31), .o(n_777) );
in01f80 g569268 ( .a(x_out_19_8), .o(n_1685) );
in01f80 g569269 ( .a(x_out_46_21), .o(n_1395) );
in01f80 g569270 ( .a(x_out_47_23), .o(n_1823) );
in01f80 g569271 ( .a(x_out_18_25), .o(n_1847) );
in01f80 g569272 ( .a(x_out_41_25), .o(n_114) );
in01f80 g569273 ( .a(x_out_38_13), .o(n_1445) );
in01f80 g569274 ( .a(x_out_21_29), .o(n_1757) );
in01f80 g569275 ( .a(x_out_54_5), .o(n_1501) );
in01f80 g569276 ( .a(x_out_40_13), .o(n_1826) );
in01f80 g569277 ( .a(x_out_32_6), .o(n_95) );
in01f80 g569278 ( .a(x_out_45_32), .o(n_109) );
in01f80 g569279 ( .a(x_out_2_0), .o(n_674) );
in01f80 g569280 ( .a(x_out_38_28), .o(n_1885) );
in01f80 g569281 ( .a(x_out_60_4), .o(n_347) );
in01f80 g569282 ( .a(x_out_37_6), .o(n_45) );
in01f80 g569283 ( .a(x_out_47_32), .o(n_1952) );
in01f80 g569284 ( .a(x_out_14_1), .o(n_1502) );
in01f80 g569285 ( .a(x_out_35_25), .o(n_1406) );
in01f80 g569286 ( .a(x_out_63_5), .o(n_1243) );
in01f80 g569287 ( .a(x_out_38_15), .o(n_1161) );
in01f80 g569288 ( .a(x_out_46_24), .o(n_153) );
in01f80 g569289 ( .a(x_out_25_12), .o(n_1704) );
in01f80 g569290 ( .a(x_out_42_13), .o(n_1788) );
in01f80 g569291 ( .a(x_out_15_18), .o(n_872) );
in01f80 g569292 ( .a(x_out_60_2), .o(n_394) );
in01f80 g569293 ( .a(x_out_45_11), .o(n_1002) );
in01f80 g569294 ( .a(x_out_26_15), .o(n_672) );
in01f80 g569295 ( .a(x_out_9_24), .o(n_1495) );
in01f80 g569296 ( .a(x_out_31_4), .o(n_1297) );
in01f80 g569297 ( .a(x_out_5_7), .o(n_208) );
in01f80 g569298 ( .a(x_out_32_15), .o(n_663) );
in01f80 g569299 ( .a(x_out_27_4), .o(n_1105) );
in01f80 g569300 ( .a(x_out_23_33), .o(n_1262) );
in01f80 g569301 ( .a(x_out_50_12), .o(n_1928) );
in01f80 g569302 ( .a(x_out_30_20), .o(n_1915) );
in01f80 g569303 ( .a(x_out_48_28), .o(n_1023) );
in01f80 g569304 ( .a(x_out_61_19), .o(n_446) );
in01f80 g569305 ( .a(x_out_53_33), .o(n_1965) );
in01f80 g569306 ( .a(x_out_47_6), .o(n_19) );
in01f80 g569307 ( .a(x_out_47_8), .o(n_831) );
in01f80 g569308 ( .a(x_out_10_24), .o(n_1858) );
in01f80 g569309 ( .a(x_out_39_27), .o(n_1504) );
in01f80 g569310 ( .a(x_out_24_9), .o(n_1232) );
in01f80 g569311 ( .a(x_out_50_6), .o(n_1412) );
in01f80 g569312 ( .a(x_out_26_25), .o(n_26) );
in01f80 g569313 ( .a(x_out_51_7), .o(n_736) );
in01f80 g569314 ( .a(x_out_60_28), .o(n_1187) );
in01f80 g569315 ( .a(x_out_1_6), .o(n_659) );
in01f80 g569316 ( .a(x_out_1_30), .o(n_487) );
in01f80 g569317 ( .a(x_out_26_12), .o(n_1039) );
in01f80 g569318 ( .a(x_out_53_27), .o(n_1475) );
in01f80 g569319 ( .a(x_out_61_33), .o(n_938) );
in01f80 g569320 ( .a(x_out_63_4), .o(n_1000) );
in01f80 g569321 ( .a(x_out_45_28), .o(n_1554) );
in01f80 g569322 ( .a(x_out_3_23), .o(n_1793) );
in01f80 g569323 ( .a(x_out_29_32), .o(n_1334) );
in01f80 g569324 ( .a(x_out_37_28), .o(n_1735) );
in01f80 g569325 ( .a(x_out_8_28), .o(n_348) );
in01f80 g569326 ( .a(x_out_60_33), .o(n_631) );
in01f80 g569327 ( .a(x_out_21_2), .o(n_577) );
in01f80 g569328 ( .a(x_out_58_4), .o(n_712) );
in01f80 g569329 ( .a(x_out_1_10), .o(n_316) );
in01f80 g569330 ( .a(x_out_3_33), .o(n_1608) );
in01f80 g569331 ( .a(x_out_41_29), .o(n_619) );
in01f80 g569332 ( .a(x_out_47_30), .o(n_628) );
in01f80 g569333 ( .a(x_out_46_7), .o(n_464) );
in01f80 g569334 ( .a(x_out_29_1), .o(n_1926) );
in01f80 g569335 ( .a(x_out_18_0), .o(n_1617) );
in01f80 g569336 ( .a(x_out_22_23), .o(n_1263) );
in01f80 g569337 ( .a(x_out_54_6), .o(n_244) );
in01f80 g569338 ( .a(x_out_25_32), .o(n_1821) );
in01f80 g569339 ( .a(x_out_58_3), .o(n_1447) );
in01f80 g569340 ( .a(x_out_63_9), .o(n_381) );
in01f80 g569341 ( .a(x_out_25_0), .o(n_724) );
in01f80 g569342 ( .a(x_out_15_8), .o(n_1222) );
in01f80 g569343 ( .a(x_out_47_29), .o(n_205) );
in01f80 g569344 ( .a(x_out_32_3), .o(n_948) );
in01f80 g569345 ( .a(x_out_61_13), .o(n_1265) );
in01f80 g569346 ( .a(x_out_53_28), .o(n_510) );
in01f80 g569347 ( .a(x_out_16_28), .o(n_1769) );
in01f80 g569348 ( .a(x_out_26_29), .o(n_1352) );
in01f80 g569349 ( .a(x_out_47_24), .o(n_1255) );
in01f80 g569350 ( .a(x_out_49_25), .o(n_366) );
in01f80 g569351 ( .a(x_out_32_13), .o(n_1814) );
in01f80 g569352 ( .a(x_out_13_0), .o(n_419) );
in01f80 g569353 ( .a(x_out_37_25), .o(n_650) );
in01f80 g569354 ( .a(x_out_8_8), .o(n_165) );
in01f80 g569355 ( .a(x_out_29_29), .o(n_1541) );
in01f80 g569356 ( .a(x_out_21_24), .o(n_146) );
in01f80 g569357 ( .a(x_out_31_11), .o(n_1152) );
in01f80 g569358 ( .a(x_out_2_33), .o(n_264) );
in01f80 g569359 ( .a(x_out_51_13), .o(n_1560) );
in01f80 g569360 ( .a(x_out_17_30), .o(n_556) );
in01f80 g569361 ( .a(x_out_8_29), .o(n_1547) );
in01f80 g569362 ( .a(x_out_43_23), .o(n_69) );
in01f80 g569363 ( .a(x_out_57_4), .o(n_1738) );
in01f80 g569364 ( .a(x_out_47_4), .o(n_874) );
in01f80 g569365 ( .a(x_out_28_4), .o(n_1782) );
in01f80 g569366 ( .a(x_out_7_29), .o(n_179) );
in01f80 g569367 ( .a(x_out_56_33), .o(n_989) );
in01f80 g569368 ( .a(x_out_14_31), .o(n_71) );
in01f80 g569369 ( .a(x_out_2_7), .o(n_496) );
in01f80 g569370 ( .a(x_out_61_27), .o(n_676) );
in01f80 g569371 ( .a(x_out_2_8), .o(n_895) );
in01f80 g569372 ( .a(x_out_17_10), .o(n_447) );
in01f80 g569373 ( .a(x_out_46_27), .o(n_266) );
in01f80 g569374 ( .a(x_out_63_26), .o(n_227) );
in01f80 g569375 ( .a(x_out_44_2), .o(n_1089) );
in01f80 g569376 ( .a(x_out_42_11), .o(n_1586) );
in01f80 g569377 ( .a(x_out_44_30), .o(n_112) );
in01f80 g569378 ( .a(x_out_33_26), .o(n_392) );
in01f80 g569379 ( .a(x_out_33_23), .o(n_875) );
in01f80 g569380 ( .a(x_out_21_11), .o(n_224) );
in01f80 g569381 ( .a(x_out_47_21), .o(n_1075) );
in01f80 g569382 ( .a(x_out_27_33), .o(n_1328) );
in01f80 g569383 ( .a(x_out_28_7), .o(n_1683) );
in01f80 g569384 ( .a(x_out_7_4), .o(n_696) );
in01f80 g569385 ( .a(x_out_19_23), .o(n_1697) );
in01f80 g569386 ( .a(x_out_5_15), .o(n_1053) );
in01f80 g569387 ( .a(x_out_61_28), .o(n_1565) );
in01f80 g569388 ( .a(x_out_17_29), .o(n_776) );
in01f80 g569389 ( .a(x_out_14_9), .o(n_477) );
in01f80 g569390 ( .a(x_out_1_1), .o(n_1916) );
in01f80 g569391 ( .a(x_out_51_3), .o(n_1528) );
in01f80 g569392 ( .a(x_out_23_11), .o(n_243) );
in01f80 g569393 ( .a(x_out_45_8), .o(n_752) );
in01f80 g569394 ( .a(x_out_46_33), .o(n_432) );
in01f80 g569395 ( .a(x_out_27_5), .o(n_1641) );
in01f80 g569396 ( .a(x_out_33_6), .o(n_1840) );
in01f80 g569397 ( .a(x_out_45_31), .o(n_1217) );
in01f80 g569398 ( .a(x_out_4_24), .o(n_866) );
in01f80 g569399 ( .a(x_out_50_29), .o(n_1650) );
in01f80 g569400 ( .a(x_out_29_4), .o(n_1512) );
in01f80 g569401 ( .a(x_out_7_25), .o(n_571) );
in01f80 g569402 ( .a(x_out_1_13), .o(n_1183) );
in01f80 g569403 ( .a(x_out_45_19), .o(n_972) );
in01f80 g569404 ( .a(x_out_30_12), .o(n_353) );
in01f80 g569405 ( .a(x_out_55_25), .o(n_670) );
in01f80 g569406 ( .a(x_out_38_14), .o(n_1121) );
in01f80 g569407 ( .a(x_out_36_25), .o(n_465) );
in01f80 g569408 ( .a(x_out_30_26), .o(n_98) );
in01f80 g569409 ( .a(x_out_11_27), .o(n_647) );
in01f80 g569410 ( .a(x_out_11_11), .o(n_1267) );
in01f80 g569411 ( .a(x_out_13_28), .o(n_1642) );
in01f80 g569412 ( .a(x_out_7_27), .o(n_106) );
in01f80 g569413 ( .a(x_out_36_18), .o(n_1375) );
in01f80 g569414 ( .a(x_out_39_20), .o(n_196) );
in01f80 g569415 ( .a(x_out_24_0), .o(n_1527) );
in01f80 g569416 ( .a(x_out_41_18), .o(n_295) );
in01f80 g569417 ( .a(x_out_39_1), .o(n_1568) );
in01f80 g569418 ( .a(x_out_43_33), .o(n_1612) );
in01f80 g569419 ( .a(x_out_18_13), .o(n_967) );
in01f80 g569420 ( .a(x_out_9_23), .o(n_1298) );
in01f80 g569421 ( .a(x_out_29_33), .o(n_325) );
in01f80 g569422 ( .a(x_out_62_33), .o(n_1129) );
in01f80 g569423 ( .a(x_out_48_32), .o(n_1466) );
in01f80 g569424 ( .a(x_out_17_0), .o(n_622) );
in01f80 g569425 ( .a(x_out_59_13), .o(n_488) );
in01f80 g569426 ( .a(x_out_5_2), .o(n_1185) );
in01f80 g569427 ( .a(x_out_38_30), .o(n_1587) );
in01f80 g569428 ( .a(x_out_17_15), .o(n_1571) );
in01f80 g569429 ( .a(x_out_4_10), .o(n_983) );
in01f80 g569430 ( .a(x_out_7_8), .o(n_1682) );
in01f80 g569431 ( .a(x_out_39_33), .o(n_1102) );
in01f80 g569432 ( .a(x_out_54_11), .o(n_1777) );
in01f80 g569433 ( .a(x_out_7_10), .o(n_70) );
in01f80 g569434 ( .a(x_out_61_26), .o(n_1734) );
in01f80 g569435 ( .a(x_out_51_6), .o(n_131) );
in01f80 g569436 ( .a(x_out_42_21), .o(n_539) );
in01f80 g569437 ( .a(x_out_11_3), .o(n_269) );
in01f80 g569438 ( .a(x_out_11_28), .o(n_1212) );
in01f80 g569439 ( .a(x_out_37_27), .o(n_110) );
in01f80 g569440 ( .a(x_out_38_6), .o(n_79) );
in01f80 g569441 ( .a(x_out_19_4), .o(n_906) );
in01f80 g569442 ( .a(x_out_17_5), .o(n_513) );
in01f80 g569443 ( .a(x_out_60_8), .o(n_599) );
in01f80 g569444 ( .a(x_out_53_32), .o(n_339) );
in01f80 g569445 ( .a(x_out_24_4), .o(n_731) );
in01f80 g569446 ( .a(x_out_8_20), .o(n_992) );
in01f80 g569447 ( .a(x_out_14_22), .o(n_1035) );
in01f80 g569448 ( .a(x_out_58_14), .o(n_1463) );
in01f80 g569449 ( .a(x_out_25_14), .o(n_1843) );
in01f80 g569450 ( .a(x_out_34_26), .o(n_572) );
in01f80 g569451 ( .a(x_out_20_12), .o(n_1503) );
in01f80 g569452 ( .a(x_out_5_27), .o(n_1186) );
in01f80 g569453 ( .a(x_out_40_10), .o(n_399) );
in01f80 g569454 ( .a(x_out_7_32), .o(n_355) );
in01f80 g569455 ( .a(x_out_25_19), .o(n_1946) );
in01f80 g569456 ( .a(x_out_15_26), .o(n_1603) );
in01f80 g569457 ( .a(x_out_46_0), .o(n_1046) );
in01f80 g569458 ( .a(x_out_60_30), .o(n_984) );
in01f80 g569459 ( .a(x_out_14_5), .o(n_1082) );
in01f80 g569460 ( .a(x_out_17_12), .o(n_965) );
in01f80 g569461 ( .a(x_out_60_13), .o(n_1496) );
in01f80 g569462 ( .a(x_out_31_2), .o(n_1385) );
in01f80 g569463 ( .a(x_out_63_3), .o(n_185) );
in01f80 g569464 ( .a(x_out_20_14), .o(n_130) );
in01f80 g569465 ( .a(x_out_43_25), .o(n_1100) );
in01f80 g569466 ( .a(x_out_25_18), .o(n_1747) );
in01f80 g569467 ( .a(x_out_8_6), .o(n_1471) );
in01f80 g569468 ( .a(x_out_19_32), .o(n_207) );
in01f80 g569469 ( .a(x_out_60_9), .o(n_1069) );
in01f80 g569470 ( .a(x_out_18_8), .o(n_1894) );
in01f80 g569471 ( .a(x_out_43_13), .o(n_1755) );
in01f80 g569472 ( .a(x_out_9_7), .o(n_1192) );
in01f80 g569473 ( .a(x_out_17_33), .o(n_1181) );
in01f80 g569474 ( .a(x_out_12_24), .o(n_117) );
in01f80 g569475 ( .a(x_out_28_30), .o(n_1356) );
in01f80 g569476 ( .a(x_out_60_19), .o(n_1580) );
in01f80 g569477 ( .a(x_out_6_33), .o(n_1292) );
in01f80 g569478 ( .a(x_out_58_11), .o(n_1931) );
in01f80 g569479 ( .a(x_out_54_18), .o(n_1210) );
in01f80 g569480 ( .a(x_out_0_14), .o(n_451) );
in01f80 g569481 ( .a(x_out_22_18), .o(n_1497) );
in01f80 g569482 ( .a(x_out_19_10), .o(n_1764) );
in01f80 g569483 ( .a(x_out_34_2), .o(n_198) );
in01f80 g569484 ( .a(x_out_34_33), .o(n_301) );
in01f80 g569485 ( .a(x_out_25_11), .o(n_630) );
in01f80 g569486 ( .a(x_out_22_0), .o(n_1329) );
in01f80 g569487 ( .a(x_out_52_5), .o(n_1786) );
in01f80 g569488 ( .a(x_out_0_15), .o(n_1111) );
in01f80 g569489 ( .a(x_out_53_7), .o(n_278) );
in01f80 g569490 ( .a(x_out_60_1), .o(n_283) );
in01f80 g569491 ( .a(x_out_30_29), .o(n_376) );
in01f80 g569492 ( .a(x_out_33_14), .o(n_1935) );
in01f80 g569493 ( .a(x_out_50_2), .o(n_1073) );
in01f80 g569494 ( .a(x_out_12_31), .o(n_1857) );
in01f80 g569495 ( .a(x_out_33_21), .o(n_461) );
in01f80 g569496 ( .a(x_out_15_12), .o(n_902) );
in01f80 g569497 ( .a(x_out_27_22), .o(n_1417) );
in01f80 g569498 ( .a(x_out_48_29), .o(n_1722) );
in01f80 g569499 ( .a(x_out_58_15), .o(n_1925) );
in01f80 g569500 ( .a(x_out_11_7), .o(n_1886) );
in01f80 g569501 ( .a(x_out_34_27), .o(n_218) );
in01f80 g569502 ( .a(x_out_49_21), .o(n_27) );
in01f80 g569503 ( .a(x_out_35_28), .o(n_1094) );
in01f80 g569504 ( .a(x_out_7_28), .o(n_1820) );
in01f80 g569505 ( .a(x_out_28_29), .o(n_143) );
in01f80 g569506 ( .a(x_out_56_3), .o(n_111) );
in01f80 g569507 ( .a(x_out_22_12), .o(n_405) );
in01f80 g569508 ( .a(x_out_38_27), .o(n_830) );
in01f80 g569509 ( .a(x_out_13_14), .o(n_1533) );
in01f80 g569510 ( .a(x_out_34_25), .o(n_917) );
in01f80 g569511 ( .a(x_out_11_13), .o(n_1071) );
in01f80 g569512 ( .a(x_out_10_18), .o(n_861) );
in01f80 g569513 ( .a(x_out_29_22), .o(n_1204) );
in01f80 g569514 ( .a(x_out_5_22), .o(n_1771) );
in01f80 g569515 ( .a(x_out_60_14), .o(n_1889) );
in01f80 g569516 ( .a(x_out_8_19), .o(n_581) );
in01f80 g569517 ( .a(x_out_23_24), .o(n_48) );
in01f80 g569518 ( .a(x_out_38_25), .o(n_560) );
in01f80 g569519 ( .a(x_out_12_9), .o(n_1353) );
in01f80 g569520 ( .a(x_out_57_27), .o(n_303) );
in01f80 g569521 ( .a(x_out_55_12), .o(n_1806) );
in01f80 g569522 ( .a(x_out_4_12), .o(n_957) );
in01f80 g569523 ( .a(x_out_37_11), .o(n_985) );
in01f80 g569524 ( .a(x_out_59_15), .o(n_1368) );
in01f80 g569525 ( .a(x_out_58_18), .o(n_431) );
in01f80 g569526 ( .a(x_out_56_32), .o(n_1966) );
in01f80 g569527 ( .a(x_out_15_4), .o(n_1566) );
in01f80 g569528 ( .a(x_out_54_3), .o(n_1327) );
in01f80 g569529 ( .a(x_out_49_11), .o(n_1621) );
in01f80 g569530 ( .a(x_out_57_18), .o(n_1728) );
in01f80 g569531 ( .a(x_out_35_30), .o(n_52) );
in01f80 g569532 ( .a(x_out_45_10), .o(n_1884) );
in01f80 g569533 ( .a(x_out_43_27), .o(n_78) );
in01f80 g569534 ( .a(x_out_2_13), .o(n_368) );
in01f80 g569535 ( .a(x_out_29_21), .o(n_645) );
in01f80 g569536 ( .a(x_out_11_31), .o(n_903) );
in01f80 g569537 ( .a(x_out_26_8), .o(n_1645) );
in01f80 g569538 ( .a(x_out_2_32), .o(n_1729) );
in01f80 g569539 ( .a(x_out_15_32), .o(n_1550) );
in01f80 g569540 ( .a(x_out_43_5), .o(n_693) );
in01f80 g569541 ( .a(x_out_28_13), .o(n_67) );
in01f80 g569542 ( .a(x_out_14_19), .o(n_707) );
in01f80 g569543 ( .a(x_out_6_6), .o(n_1369) );
in01f80 g569544 ( .a(x_out_11_22), .o(n_1241) );
in01f80 g569545 ( .a(x_out_35_9), .o(n_606) );
in01f80 g569546 ( .a(x_out_42_23), .o(n_408) );
in01f80 g569547 ( .a(x_out_58_19), .o(n_913) );
in01f80 g569548 ( .a(x_out_45_22), .o(n_1154) );
in01f80 g569549 ( .a(x_out_57_28), .o(n_926) );
in01f80 g569550 ( .a(x_out_31_15), .o(n_273) );
in01f80 g569551 ( .a(x_out_54_8), .o(n_1208) );
in01f80 g569552 ( .a(x_out_13_5), .o(n_873) );
in01f80 g569553 ( .a(x_out_26_30), .o(n_300) );
in01f80 g569554 ( .a(x_out_15_25), .o(n_1401) );
in01f80 g569555 ( .a(x_out_13_12), .o(n_1246) );
in01f80 g569556 ( .a(x_out_15_30), .o(n_946) );
in01f80 g569557 ( .a(x_out_45_25), .o(n_1675) );
in01f80 g569558 ( .a(x_out_4_33), .o(n_1415) );
in01f80 g569559 ( .a(x_out_35_22), .o(n_901) );
in01f80 g569560 ( .a(x_out_15_23), .o(n_1478) );
in01f80 g569561 ( .a(x_out_29_20), .o(n_870) );
in01f80 g569562 ( .a(x_out_54_32), .o(n_321) );
in01f80 g569563 ( .a(x_out_19_9), .o(n_634) );
in01f80 g569564 ( .a(x_out_6_14), .o(n_1498) );
in01f80 g569565 ( .a(x_out_6_30), .o(n_1745) );
in01f80 g569566 ( .a(x_out_38_18), .o(n_1920) );
in01f80 g569567 ( .a(x_out_9_25), .o(n_1523) );
in01f80 g569568 ( .a(x_out_54_4), .o(n_1379) );
in01f80 g569569 ( .a(x_out_51_22), .o(n_1910) );
in01f80 g569570 ( .a(x_out_32_11), .o(n_1595) );
in01f80 g569571 ( .a(x_out_14_33), .o(n_1629) );
in01f80 g569572 ( .a(x_out_31_1), .o(n_68) );
in01f80 g569573 ( .a(x_out_57_19), .o(n_230) );
in01f80 g569574 ( .a(x_out_41_23), .o(n_61) );
in01f80 g569575 ( .a(x_out_13_8), .o(n_400) );
in01f80 g569576 ( .a(x_out_36_26), .o(n_535) );
in01f80 g569577 ( .a(x_out_24_12), .o(n_332) );
in01f80 g569578 ( .a(x_out_18_1), .o(n_583) );
in01f80 g569579 ( .a(x_out_54_31), .o(n_327) );
in01f80 g569580 ( .a(x_out_30_23), .o(n_705) );
in01f80 g569581 ( .a(x_out_9_1), .o(n_141) );
in01f80 g569582 ( .a(x_out_52_4), .o(n_1291) );
in01f80 g569583 ( .a(x_out_20_2), .o(n_261) );
in01f80 g569584 ( .a(x_out_11_1), .o(n_925) );
in01f80 g569585 ( .a(x_out_27_20), .o(n_466) );
in01f80 g569586 ( .a(x_out_38_1), .o(n_338) );
in01f80 g569587 ( .a(x_out_19_7), .o(n_418) );
in01f80 g569588 ( .a(x_out_56_27), .o(n_1849) );
in01f80 g569589 ( .a(x_out_1_15), .o(n_164) );
in01f80 g569590 ( .a(x_out_41_8), .o(n_1610) );
in01f80 g569591 ( .a(x_out_48_8), .o(n_1893) );
in01f80 g569592 ( .a(x_out_26_22), .o(n_920) );
in01f80 g569593 ( .a(x_out_55_18), .o(n_1594) );
in01f80 g569594 ( .a(x_out_56_12), .o(n_62) );
in01f80 g569595 ( .a(x_out_9_22), .o(n_1521) );
in01f80 g569596 ( .a(x_out_1_33), .o(n_745) );
in01f80 g569597 ( .a(x_out_39_6), .o(n_297) );
in01f80 g569598 ( .a(x_out_17_14), .o(n_911) );
in01f80 g569599 ( .a(x_out_41_30), .o(n_692) );
in01f80 g569600 ( .a(x_out_0_10), .o(n_485) );
in01f80 g569601 ( .a(x_out_57_15), .o(n_704) );
in01f80 g569602 ( .a(x_out_14_7), .o(n_202) );
in01f80 g569603 ( .a(x_out_4_19), .o(n_1331) );
in01f80 g569604 ( .a(x_out_34_9), .o(n_507) );
in01f80 g569605 ( .a(x_out_12_5), .o(n_1750) );
in01f80 g569606 ( .a(x_out_22_30), .o(n_1758) );
in01f80 g569607 ( .a(x_out_38_20), .o(n_545) );
in01f80 g569608 ( .a(x_out_47_27), .o(n_1157) );
in01f80 g569609 ( .a(x_out_25_6), .o(n_1538) );
in01f80 g569610 ( .a(x_out_35_7), .o(n_1876) );
in01f80 g569611 ( .a(x_out_24_25), .o(n_580) );
in01f80 g569612 ( .a(x_out_49_33), .o(n_509) );
in01f80 g569613 ( .a(x_out_1_29), .o(n_773) );
in01f80 g569614 ( .a(x_out_21_18), .o(n_1083) );
in01f80 g569615 ( .a(x_out_57_13), .o(n_40) );
in01f80 g569616 ( .a(x_out_63_30), .o(n_1549) );
in01f80 g569617 ( .a(x_out_25_3), .o(n_1567) );
in01f80 g569618 ( .a(x_out_26_9), .o(n_1859) );
in01f80 g569619 ( .a(x_out_1_7), .o(n_878) );
in01f80 g569620 ( .a(x_out_19_14), .o(n_1174) );
in01f80 g569621 ( .a(x_out_45_33), .o(n_287) );
in01f80 g569622 ( .a(x_out_22_4), .o(n_754) );
in01f80 g569623 ( .a(x_out_35_2), .o(n_624) );
in01f80 g569624 ( .a(x_out_47_28), .o(n_1199) );
in01f80 g569625 ( .a(x_out_9_21), .o(n_152) );
in01f80 g569626 ( .a(x_out_8_26), .o(n_380) );
in01f80 g569627 ( .a(x_out_46_11), .o(n_1170) );
in01f80 g569628 ( .a(x_out_30_31), .o(n_1097) );
in01f80 g569629 ( .a(x_out_12_33), .o(n_689) );
in01f80 g569630 ( .a(x_out_35_24), .o(n_76) );
in01f80 g569631 ( .a(x_out_63_6), .o(n_282) );
in01f80 g569632 ( .a(x_out_30_15), .o(n_675) );
in01f80 g569633 ( .a(x_out_8_21), .o(n_519) );
in01f80 g569634 ( .a(x_out_15_9), .o(n_1534) );
in01f80 g569635 ( .a(x_out_13_10), .o(n_715) );
in01f80 g569636 ( .a(x_out_48_4), .o(n_1090) );
in01f80 g569637 ( .a(x_out_18_14), .o(n_1114) );
in01f80 g569638 ( .a(x_out_49_2), .o(n_869) );
in01f80 g569639 ( .a(x_out_4_8), .o(n_637) );
in01f80 g569640 ( .a(x_out_3_31), .o(n_1604) );
in01f80 g569641 ( .a(x_out_20_3), .o(n_618) );
in01f80 g569642 ( .a(x_out_40_27), .o(n_1488) );
in01f80 g569643 ( .a(x_out_40_26), .o(n_1955) );
in01f80 g569644 ( .a(x_out_10_30), .o(n_1382) );
in01f80 g569645 ( .a(x_out_28_10), .o(n_281) );
in01f80 g569646 ( .a(x_out_13_15), .o(n_341) );
in01f80 g569647 ( .a(x_out_39_9), .o(n_1932) );
in01f80 g569648 ( .a(x_out_40_30), .o(n_783) );
in01f80 g569649 ( .a(x_out_44_9), .o(n_270) );
in01f80 g569650 ( .a(x_out_9_6), .o(n_1310) );
in01f80 g569651 ( .a(x_out_62_22), .o(n_666) );
in01f80 g569652 ( .a(x_out_59_29), .o(n_302) );
in01f80 g569653 ( .a(x_out_48_0), .o(n_654) );
in01f80 g569654 ( .a(x_out_45_2), .o(n_594) );
in01f80 g569655 ( .a(x_out_16_27), .o(n_1655) );
in01f80 g569656 ( .a(x_out_26_7), .o(n_951) );
in01f80 g569657 ( .a(x_out_50_7), .o(n_1516) );
in01f80 g569658 ( .a(x_out_43_4), .o(n_1215) );
in01f80 g569659 ( .a(x_out_50_10), .o(n_1044) );
in01f80 g569660 ( .a(x_out_32_5), .o(n_923) );
in01f80 g569661 ( .a(x_out_34_32), .o(n_1939) );
in01f80 g569662 ( .a(x_out_30_8), .o(n_1254) );
in01f80 g569663 ( .a(x_out_40_28), .o(n_661) );
in01f80 g569664 ( .a(x_out_48_7), .o(n_1838) );
in01f80 g569665 ( .a(x_out_42_7), .o(n_175) );
in01f80 g569666 ( .a(x_out_16_8), .o(n_1286) );
in01f80 g569667 ( .a(x_out_57_12), .o(n_1119) );
in01f80 g569668 ( .a(x_out_4_13), .o(n_949) );
in01f80 g569669 ( .a(x_out_5_0), .o(n_710) );
in01f80 g569670 ( .a(x_out_14_29), .o(n_126) );
in01f80 g569671 ( .a(x_out_29_27), .o(n_1322) );
in01f80 g569672 ( .a(x_out_10_1), .o(n_139) );
in01f80 g569673 ( .a(x_out_12_23), .o(n_975) );
in01f80 g569674 ( .a(x_out_45_20), .o(n_1031) );
in01f80 g569675 ( .a(x_out_40_4), .o(n_950) );
in01f80 g569676 ( .a(x_out_26_6), .o(n_304) );
in01f80 g569677 ( .a(x_out_23_7), .o(n_803) );
in01f80 g569678 ( .a(x_out_63_19), .o(n_882) );
in01f80 g569679 ( .a(x_out_55_26), .o(n_1446) );
in01f80 g569680 ( .a(x_out_17_3), .o(n_148) );
in01f80 g569681 ( .a(x_out_63_22), .o(n_145) );
in01f80 g569682 ( .a(x_out_39_3), .o(n_424) );
in01f80 g569683 ( .a(x_out_16_12), .o(n_1929) );
in01f80 g569684 ( .a(x_out_60_7), .o(n_1691) );
in01f80 g569685 ( .a(x_out_14_24), .o(n_1742) );
in01f80 g569686 ( .a(x_out_13_6), .o(n_501) );
in01f80 g569687 ( .a(x_out_40_1), .o(n_308) );
in01f80 g569688 ( .a(x_out_53_0), .o(n_286) );
in01f80 g569689 ( .a(x_out_6_20), .o(n_1829) );
in01f80 g569690 ( .a(x_out_50_9), .o(n_239) );
in01f80 g569691 ( .a(x_out_23_30), .o(n_815) );
in01f80 g569692 ( .a(x_out_9_13), .o(n_105) );
in01f80 g569693 ( .a(x_out_12_30), .o(n_542) );
in01f80 g569694 ( .a(x_out_7_33), .o(n_836) );
in01f80 g569695 ( .a(x_out_0_8), .o(n_881) );
in01f80 g569696 ( .a(x_out_31_6), .o(n_1866) );
in01f80 g569697 ( .a(x_out_18_6), .o(n_4) );
in01f80 g569698 ( .a(x_out_21_15), .o(n_486) );
in01f80 g569699 ( .a(x_out_16_1), .o(n_99) );
in01f80 g569700 ( .a(x_out_29_19), .o(n_1151) );
in01f80 g569701 ( .a(x_out_49_20), .o(n_1834) );
in01f80 g569702 ( .a(x_out_28_21), .o(n_1948) );
in01f80 g569703 ( .a(x_out_56_18), .o(n_1223) );
in01f80 g569704 ( .a(x_out_32_0), .o(n_223) );
in01f80 g569705 ( .a(x_out_23_4), .o(n_23) );
in01f80 g569706 ( .a(x_out_46_14), .o(n_732) );
in01f80 g569707 ( .a(x_out_19_24), .o(n_1197) );
in01f80 g569708 ( .a(x_out_55_22), .o(n_441) );
in01f80 g569709 ( .a(x_out_2_20), .o(n_1633) );
in01f80 g569710 ( .a(x_out_28_12), .o(n_1971) );
in01f80 g569711 ( .a(x_out_52_6), .o(n_1781) );
in01f80 g569712 ( .a(x_out_24_24), .o(n_1008) );
in01f80 g569713 ( .a(x_out_43_10), .o(n_1231) );
in01f80 g569714 ( .a(x_out_54_20), .o(n_1600) );
in01f80 g569715 ( .a(x_out_14_2), .o(n_1491) );
in01f80 g569716 ( .a(x_out_41_10), .o(n_1440) );
in01f80 g569717 ( .a(x_out_48_6), .o(n_1067) );
in01f80 g569718 ( .a(x_out_10_32), .o(n_1726) );
in01f80 g569719 ( .a(x_out_33_3), .o(n_811) );
in01f80 g569720 ( .a(x_out_43_0), .o(n_1155) );
in01f80 g569721 ( .a(x_out_24_31), .o(n_1427) );
in01f80 g569722 ( .a(x_out_8_12), .o(n_1741) );
in01f80 g569723 ( .a(x_out_13_32), .o(n_204) );
in01f80 g569724 ( .a(x_out_56_20), .o(n_1562) );
in01f80 g569725 ( .a(x_out_58_7), .o(n_1236) );
in01f80 g569726 ( .a(x_out_56_14), .o(n_1901) );
in01f80 g569727 ( .a(x_out_6_10), .o(n_1805) );
in01f80 g569728 ( .a(x_out_10_11), .o(n_433) );
in01f80 g569729 ( .a(x_out_52_7), .o(n_505) );
in01f80 g569730 ( .a(x_out_54_14), .o(n_1041) );
in01f80 g569731 ( .a(x_out_4_20), .o(n_1593) );
in01f80 g569732 ( .a(x_out_49_10), .o(n_276) );
in01f80 g569733 ( .a(x_out_23_10), .o(n_753) );
in01f80 g569734 ( .a(x_out_59_26), .o(n_1315) );
in01f80 g569735 ( .a(x_out_53_18), .o(n_685) );
in01f80 g569736 ( .a(x_out_58_1), .o(n_1224) );
in01f80 g569737 ( .a(x_out_29_5), .o(n_193) );
in01f80 g569738 ( .a(x_out_0_13), .o(n_1967) );
in01f80 g569739 ( .a(x_out_6_32), .o(n_536) );
in01f80 g569740 ( .a(x_out_15_15), .o(n_242) );
in01f80 g569741 ( .a(x_out_18_22), .o(n_1086) );
in01f80 g569742 ( .a(x_out_12_12), .o(n_305) );
in01f80 g569743 ( .a(x_out_31_12), .o(n_228) );
in01f80 g569744 ( .a(x_out_33_29), .o(n_860) );
in01f80 g569745 ( .a(x_out_16_15), .o(n_1831) );
in01f80 g569746 ( .a(x_out_24_14), .o(n_1325) );
in01f80 g569747 ( .a(x_out_51_0), .o(n_822) );
in01f80 g569748 ( .a(x_out_13_33), .o(n_1483) );
in01f80 g569749 ( .a(x_out_47_22), .o(n_772) );
in01f80 g569750 ( .a(x_out_44_27), .o(n_1436) );
in01f80 g569751 ( .a(x_out_61_14), .o(n_1469) );
in01f80 g569752 ( .a(x_out_12_10), .o(n_1317) );
in01f80 g569753 ( .a(x_out_9_12), .o(n_1413) );
in01f80 g569754 ( .a(x_out_43_24), .o(n_1272) );
in01f80 g569755 ( .a(x_out_51_31), .o(n_1308) );
in01f80 g569756 ( .a(x_out_27_2), .o(n_936) );
in01f80 g569757 ( .a(x_out_15_29), .o(n_1717) );
in01f80 g569758 ( .a(x_out_12_11), .o(n_559) );
in01f80 g569759 ( .a(x_out_12_28), .o(n_1126) );
in01f80 g569760 ( .a(x_out_58_6), .o(n_1370) );
in01f80 g569761 ( .a(x_out_50_22), .o(n_887) );
in01f80 g569762 ( .a(x_out_25_20), .o(n_1839) );
in01f80 g569763 ( .a(x_out_30_10), .o(n_1947) );
in01f80 g569764 ( .a(x_out_42_14), .o(n_1030) );
in01f80 g569765 ( .a(x_out_24_8), .o(n_819) );
in01f80 g569766 ( .a(x_out_62_26), .o(n_369) );
in01f80 g569767 ( .a(x_out_3_18), .o(n_758) );
in01f80 g569768 ( .a(x_out_34_15), .o(n_697) );
in01f80 g569769 ( .a(x_out_9_32), .o(n_698) );
in01f80 g569770 ( .a(x_out_61_30), .o(n_97) );
in01f80 g569771 ( .a(x_out_19_18), .o(n_364) );
in01f80 g569772 ( .a(x_out_4_5), .o(n_974) );
in01f80 g569773 ( .a(x_out_17_11), .o(n_843) );
in01f80 g569774 ( .a(x_out_0_6), .o(n_1147) );
in01f80 g569775 ( .a(x_out_54_33), .o(n_796) );
in01f80 g569776 ( .a(x_out_22_32), .o(n_765) );
in01f80 g569777 ( .a(x_out_34_28), .o(n_899) );
in01f80 g569778 ( .a(x_out_30_19), .o(n_1732) );
in01f80 g569779 ( .a(x_out_27_3), .o(n_383) );
in01f80 g569780 ( .a(x_out_57_24), .o(n_1481) );
in01f80 g569781 ( .a(x_out_40_11), .o(n_640) );
in01f80 g569782 ( .a(x_out_4_30), .o(n_1045) );
in01f80 g569783 ( .a(x_out_37_24), .o(n_832) );
in01f80 g569784 ( .a(x_out_58_2), .o(n_764) );
in01f80 g569785 ( .a(x_out_24_7), .o(n_1047) );
in01f80 g569786 ( .a(x_out_52_15), .o(n_932) );
in01f80 g569787 ( .a(x_out_44_22), .o(n_1160) );
in01f80 g569788 ( .a(x_out_7_6), .o(n_91) );
in01f80 g569789 ( .a(x_out_25_26), .o(n_1459) );
in01f80 g569790 ( .a(x_out_28_1), .o(n_1634) );
in01f80 g569791 ( .a(x_out_62_0), .o(n_1431) );
in01f80 g569792 ( .a(x_out_9_33), .o(n_981) );
in01f80 g569793 ( .a(x_out_21_3), .o(n_1713) );
in01f80 g569794 ( .a(x_out_44_6), .o(n_1249) );
in01f80 g569795 ( .a(x_out_57_3), .o(n_718) );
in01f80 g569796 ( .a(x_out_7_18), .o(n_3) );
in01f80 g569797 ( .a(x_out_35_6), .o(n_747) );
in01f80 g569798 ( .a(x_out_53_4), .o(n_1242) );
in01f80 g569799 ( .a(x_out_40_12), .o(n_612) );
in01f80 g569800 ( .a(x_out_34_18), .o(n_1585) );
in01f80 g569801 ( .a(x_out_37_14), .o(n_1018) );
in01f80 g569802 ( .a(x_out_5_31), .o(n_1709) );
in01f80 g569803 ( .a(x_out_9_31), .o(n_1372) );
in01f80 g569804 ( .a(x_out_38_5), .o(n_845) );
in01f80 g569805 ( .a(x_out_53_9), .o(n_837) );
in01f80 g569806 ( .a(x_out_42_6), .o(n_33) );
in01f80 g569807 ( .a(x_out_48_25), .o(n_437) );
in01f80 g569808 ( .a(x_out_10_7), .o(n_1694) );
in01f80 g569809 ( .a(x_out_63_28), .o(n_1384) );
in01f80 g569810 ( .a(x_out_44_5), .o(n_1783) );
in01f80 g569811 ( .a(x_out_62_27), .o(n_930) );
in01f80 g569812 ( .a(x_out_62_29), .o(n_1813) );
in01f80 g569813 ( .a(x_out_53_26), .o(n_1877) );
in01f80 g569814 ( .a(x_out_62_8), .o(n_512) );
in01f80 g569815 ( .a(x_out_26_23), .o(n_1970) );
in01f80 g569816 ( .a(x_out_51_9), .o(n_1376) );
in01f80 g569817 ( .a(x_out_42_33), .o(n_1825) );
in01f80 g569818 ( .a(x_out_29_10), .o(n_1708) );
in01f80 g569819 ( .a(x_out_27_13), .o(n_789) );
in01f80 g569820 ( .a(x_out_56_23), .o(n_1828) );
in01f80 g569821 ( .a(x_out_17_9), .o(n_1647) );
in01f80 g569822 ( .a(x_out_27_32), .o(n_1652) );
in01f80 g569823 ( .a(x_out_17_1), .o(n_1880) );
in01f80 g569824 ( .a(x_out_19_28), .o(n_1797) );
in01f80 g569825 ( .a(x_out_18_19), .o(n_1077) );
in01f80 g569826 ( .a(x_out_22_10), .o(n_1579) );
in01f80 g569827 ( .a(x_out_31_5), .o(n_1040) );
in01f80 g569828 ( .a(x_out_56_21), .o(n_636) );
in01f80 g569829 ( .a(x_out_34_29), .o(n_176) );
in01f80 g569830 ( .a(x_out_33_24), .o(n_1085) );
in01f80 g569831 ( .a(x_out_35_10), .o(n_1342) );
in01f80 g569832 ( .a(x_out_46_15), .o(n_1693) );
in01f80 g569833 ( .a(x_out_25_2), .o(n_1116) );
in01f80 g569834 ( .a(x_out_15_2), .o(n_1205) );
in01f80 g569835 ( .a(x_out_49_5), .o(n_138) );
in01f80 g569836 ( .a(x_out_3_26), .o(n_1028) );
in01f80 g569837 ( .a(x_out_48_13), .o(n_22) );
in01f80 g569838 ( .a(x_out_5_4), .o(n_1338) );
in01f80 g569839 ( .a(x_out_45_27), .o(n_1651) );
in01f80 g569840 ( .a(x_out_19_27), .o(n_319) );
in01f80 g569841 ( .a(x_out_39_0), .o(n_313) );
in01f80 g569842 ( .a(x_out_58_10), .o(n_1416) );
in01f80 g569843 ( .a(x_out_20_0), .o(n_147) );
in01f80 g569844 ( .a(x_out_50_33), .o(n_217) );
in01f80 g569845 ( .a(x_out_21_31), .o(n_1801) );
in01f80 g569846 ( .a(x_out_49_0), .o(n_527) );
in01f80 g569847 ( .a(x_out_16_13), .o(n_251) );
in01f80 g569848 ( .a(x_out_4_6), .o(n_210) );
in01f80 g569849 ( .a(x_out_23_0), .o(n_1622) );
in01f80 g569850 ( .a(x_out_60_12), .o(n_459) );
in01f80 g569851 ( .a(x_out_63_11), .o(n_853) );
in01f80 g569852 ( .a(x_out_43_31), .o(n_1702) );
in01f80 g569853 ( .a(x_out_52_0), .o(n_272) );
in01f80 g569854 ( .a(x_out_22_1), .o(n_1917) );
in01f80 g569855 ( .a(x_out_43_18), .o(n_921) );
in01f80 g569856 ( .a(x_out_63_8), .o(n_258) );
in01f80 g569857 ( .a(x_out_38_23), .o(n_1677) );
in01f80 g569858 ( .a(x_out_49_3), .o(n_1457) );
in01f80 g569859 ( .a(x_out_43_20), .o(n_1712) );
in01f80 g569860 ( .a(x_out_41_21), .o(n_586) );
in01f80 g569861 ( .a(x_out_48_26), .o(n_1835) );
in01f80 g569862 ( .a(x_out_50_21), .o(n_928) );
in01f80 g569863 ( .a(x_out_59_14), .o(n_1134) );
in01f80 g569864 ( .a(x_out_10_31), .o(n_219) );
in01f80 g569865 ( .a(x_out_9_30), .o(n_1048) );
in01f80 g569866 ( .a(x_out_30_14), .o(n_1364) );
in01f80 g569867 ( .a(x_out_61_9), .o(n_1316) );
in01f80 g569868 ( .a(x_out_14_28), .o(n_1526) );
in01f80 g569869 ( .a(x_out_50_23), .o(n_407) );
in01f80 g569870 ( .a(x_out_18_10), .o(n_1244) );
in01f80 g569871 ( .a(x_out_14_3), .o(n_1627) );
in01f80 g569872 ( .a(x_out_1_9), .o(n_979) );
in01f80 g569873 ( .a(x_out_33_20), .o(n_939) );
in01f80 g569874 ( .a(x_out_48_14), .o(n_1451) );
in01f80 g569875 ( .a(x_out_24_11), .o(n_1542) );
in01f80 g569876 ( .a(x_out_31_31), .o(n_1280) );
in01f80 g569877 ( .a(x_out_58_32), .o(n_1163) );
in01f80 g569878 ( .a(x_out_21_27), .o(n_1630) );
in01f80 g569879 ( .a(x_out_10_20), .o(n_727) );
in01f80 g569880 ( .a(x_out_46_32), .o(n_1321) );
in01f80 g569881 ( .a(x_out_46_30), .o(n_229) );
in01f80 g569882 ( .a(x_out_50_31), .o(n_372) );
in01f80 g569883 ( .a(x_out_62_7), .o(n_1269) );
in01f80 g569884 ( .a(x_out_34_0), .o(n_221) );
in01f80 g569885 ( .a(x_out_51_21), .o(n_1117) );
in01f80 g569886 ( .a(x_out_22_19), .o(n_978) );
in01f80 g569887 ( .a(x_out_40_7), .o(n_215) );
in01f80 g569888 ( .a(x_out_5_8), .o(n_1275) );
in01f80 g569889 ( .a(x_out_25_7), .o(n_1874) );
in01f80 g569890 ( .a(x_out_36_1), .o(n_1214) );
in01f80 g569891 ( .a(x_out_43_2), .o(n_1010) );
in01f80 g569892 ( .a(x_out_40_31), .o(n_309) );
in01f80 g569893 ( .a(x_out_49_24), .o(n_1553) );
in01f80 g569894 ( .a(x_out_49_14), .o(n_1625) );
in01f80 g569895 ( .a(x_out_7_5), .o(n_728) );
in01f80 g569896 ( .a(x_out_12_22), .o(n_1284) );
in01f80 g569897 ( .a(x_out_51_27), .o(n_136) );
in01f80 g569898 ( .a(x_out_34_11), .o(n_1127) );
in01f80 g569899 ( .a(x_out_50_24), .o(n_529) );
in01f80 g569900 ( .a(x_out_3_11), .o(n_1153) );
in01f80 g569901 ( .a(x_out_37_13), .o(n_296) );
in01f80 g569902 ( .a(x_out_54_12), .o(n_1911) );
in01f80 g569903 ( .a(x_out_8_14), .o(n_655) );
in01f80 g569904 ( .a(x_out_0_9), .o(n_1404) );
in01f80 g569905 ( .a(x_out_28_26), .o(n_958) );
in01f80 g569906 ( .a(x_out_42_29), .o(n_849) );
in01f80 g569907 ( .a(x_out_62_15), .o(n_17) );
in01f80 g569908 ( .a(x_out_9_29), .o(n_1145) );
in01f80 g569909 ( .a(x_out_16_18), .o(n_1115) );
in01f80 g569910 ( .a(x_out_23_32), .o(n_1330) );
in01f80 g569911 ( .a(x_out_6_11), .o(n_1508) );
in01f80 g569912 ( .a(x_out_53_31), .o(n_397) );
in01f80 g569913 ( .a(x_out_10_12), .o(n_563) );
in01f80 g569914 ( .a(x_out_16_7), .o(n_1907) );
in01f80 g569915 ( .a(x_out_22_15), .o(n_1563) );
in01f80 g569916 ( .a(x_out_63_0), .o(n_1107) );
in01f80 g569917 ( .a(x_out_21_33), .o(n_1219) );
in01f80 g569918 ( .a(x_out_56_0), .o(n_200) );
in01f80 g569919 ( .a(x_out_62_19), .o(n_162) );
in01f80 g569920 ( .a(x_out_52_10), .o(n_57) );
in01f80 g569921 ( .a(x_out_27_29), .o(n_1421) );
in01f80 g569922 ( .a(x_out_20_13), .o(n_717) );
in01f80 g569923 ( .a(x_out_29_12), .o(n_814) );
in01f80 g569924 ( .a(x_out_13_3), .o(n_827) );
in01f80 g569925 ( .a(x_out_5_1), .o(n_660) );
in01f80 g569926 ( .a(x_out_16_10), .o(n_250) );
in01f80 g569927 ( .a(x_out_16_0), .o(n_714) );
in01f80 g569928 ( .a(x_out_25_10), .o(n_1794) );
in01f80 g569929 ( .a(x_out_23_13), .o(n_86) );
in01f80 g569930 ( .a(x_out_29_23), .o(n_744) );
in01f80 g569931 ( .a(x_out_12_15), .o(n_1898) );
in01f80 g569932 ( .a(x_out_37_2), .o(n_605) );
in01f80 g569933 ( .a(x_out_39_4), .o(n_1309) );
in01f80 g569934 ( .a(x_out_32_8), .o(n_893) );
in01f80 g569935 ( .a(x_out_6_23), .o(n_615) );
in01f80 g569936 ( .a(x_out_37_30), .o(n_785) );
in01f80 g569937 ( .a(x_out_53_25), .o(n_83) );
in01f80 g569938 ( .a(x_out_2_27), .o(n_582) );
in01f80 g569939 ( .a(x_out_21_0), .o(n_241) );
in01f80 g569940 ( .a(x_out_2_11), .o(n_1492) );
in01f80 g569941 ( .a(x_out_13_18), .o(n_498) );
in01f80 g569942 ( .a(x_out_47_9), .o(n_730) );
in01f80 g569943 ( .a(x_out_10_28), .o(n_255) );
in01f80 g569944 ( .a(x_out_37_26), .o(n_1296) );
in01f80 g569945 ( .a(x_out_45_15), .o(n_664) );
in01f80 g569946 ( .a(x_out_23_31), .o(n_1337) );
in01f80 g569947 ( .a(x_out_0_1), .o(n_1392) );
in01f80 g569948 ( .a(x_out_61_3), .o(n_1476) );
in01f80 g569949 ( .a(x_out_55_7), .o(n_39) );
in01f80 g569950 ( .a(x_out_43_8), .o(n_298) );
in01f80 g569951 ( .a(x_out_5_30), .o(n_1020) );
in01f80 g569952 ( .a(x_out_9_18), .o(n_1490) );
in01f80 g569953 ( .a(x_out_29_11), .o(n_1306) );
in01f80 g569954 ( .a(x_out_12_26), .o(n_30) );
in01f80 g569955 ( .a(x_out_3_10), .o(n_1374) );
in01f80 g569956 ( .a(x_out_31_10), .o(n_1854) );
in01f80 g569957 ( .a(x_out_31_14), .o(n_716) );
in01f80 g569958 ( .a(x_out_50_14), .o(n_568) );
in01f80 g569959 ( .a(x_out_44_26), .o(n_415) );
in01f80 g569960 ( .a(x_out_19_31), .o(n_167) );
in01f80 g569961 ( .a(x_out_39_14), .o(n_474) );
in01f80 g569962 ( .a(x_out_41_11), .o(n_567) );
in01f80 g569963 ( .a(x_out_58_27), .o(n_214) );
in01f80 g569964 ( .a(x_out_23_14), .o(n_757) );
in01f80 g569965 ( .a(x_out_4_9), .o(n_1003) );
in01f80 g569966 ( .a(x_out_46_12), .o(n_947) );
in01f80 g569967 ( .a(x_out_48_11), .o(n_1795) );
in01f80 g569968 ( .a(x_out_12_20), .o(n_910) );
in01f80 g569969 ( .a(x_out_17_6), .o(n_534) );
in01f80 g569970 ( .a(x_out_2_30), .o(n_668) );
in01f80 g569971 ( .a(x_out_38_3), .o(n_871) );
in01f80 g569972 ( .a(x_out_41_1), .o(n_416) );
in01f80 g569973 ( .a(x_out_57_5), .o(n_851) );
in01f80 g569974 ( .a(x_out_34_5), .o(n_323) );
in01f80 g569975 ( .a(x_out_63_27), .o(n_1013) );
in01f80 g569976 ( .a(x_out_3_15), .o(n_1776) );
in01f80 g569977 ( .a(x_out_17_19), .o(n_1144) );
in01f80 g569978 ( .a(x_out_6_27), .o(n_695) );
in01f80 g569979 ( .a(x_out_35_3), .o(n_1954) );
in01f80 g569980 ( .a(x_out_19_15), .o(n_1546) );
in01f80 g569981 ( .a(x_out_21_9), .o(n_1092) );
in01f80 g569982 ( .a(x_out_36_12), .o(n_620) );
in01f80 g569983 ( .a(x_out_49_31), .o(n_1283) );
in01f80 g569984 ( .a(x_out_34_13), .o(n_404) );
in01f80 g569985 ( .a(x_out_54_19), .o(n_1513) );
in01f80 g569986 ( .a(x_out_7_26), .o(n_336) );
in01f80 g569987 ( .a(x_out_42_5), .o(n_1596) );
in01f80 g569988 ( .a(x_out_12_25), .o(n_658) );
in01f80 g569989 ( .a(x_out_5_32), .o(n_800) );
in01f80 g569990 ( .a(x_out_28_24), .o(n_1150) );
in01f80 g569991 ( .a(x_out_55_1), .o(n_548) );
in01f80 g569992 ( .a(x_out_29_13), .o(n_1194) );
in01f80 g569993 ( .a(x_out_3_3), .o(n_1424) );
in01f80 g569994 ( .a(x_out_39_30), .o(n_1660) );
in01f80 g569995 ( .a(x_out_43_1), .o(n_986) );
in01f80 g569996 ( .a(x_out_45_26), .o(n_310) );
in01f80 g569997 ( .a(x_out_6_18), .o(n_390) );
in01f80 g569998 ( .a(x_out_0_5), .o(n_1428) );
in01f80 g569999 ( .a(x_out_63_20), .o(n_1574) );
in01f80 g570000 ( .a(x_out_15_19), .o(n_1930) );
in01f80 g570001 ( .a(x_out_45_9), .o(n_1964) );
in01f80 g570002 ( .a(x_out_28_5), .o(n_1500) );
in01f80 g570003 ( .a(x_out_26_27), .o(n_1973) );
in01f80 g570004 ( .a(x_out_28_28), .o(n_1009) );
in01f80 g570005 ( .a(x_out_48_22), .o(n_934) );
in01f80 g570006 ( .a(x_out_38_4), .o(n_314) );
in01f80 g570007 ( .a(x_out_37_3), .o(n_1590) );
in01f80 g570008 ( .a(x_out_37_12), .o(n_361) );
in01f80 g570009 ( .a(x_out_55_28), .o(n_56) );
in01f80 g570010 ( .a(x_out_46_29), .o(n_32) );
in01f80 g570011 ( .a(x_out_9_20), .o(n_587) );
in01f80 g570012 ( .a(x_out_48_1), .o(n_1371) );
in01f80 g570013 ( .a(x_out_0_11), .o(n_929) );
in01f80 g570014 ( .a(x_out_33_15), .o(n_1945) );
in01f80 g570015 ( .a(x_out_8_24), .o(n_629) );
in01f80 g570016 ( .a(x_out_19_2), .o(n_824) );
in01f80 g570017 ( .a(x_out_14_4), .o(n_342) );
in01f80 g570018 ( .a(x_out_56_11), .o(n_966) );
in01f80 g570019 ( .a(x_out_13_27), .o(n_1638) );
in01f80 g570020 ( .a(x_out_50_0), .o(n_190) );
in01f80 g570021 ( .a(x_out_48_20), .o(n_51) );
in01f80 g570022 ( .a(x_out_55_13), .o(n_1944) );
in01f80 g570023 ( .a(x_out_13_23), .o(n_393) );
in01f80 g570024 ( .a(x_out_8_4), .o(n_1656) );
in01f80 g570025 ( .a(x_out_50_26), .o(n_1201) );
in01f80 g570026 ( .a(x_out_11_33), .o(n_1517) );
in01f80 g570027 ( .a(x_out_23_18), .o(n_994) );
in01f80 g570028 ( .a(x_out_31_18), .o(n_15) );
in01f80 g570029 ( .a(x_out_29_25), .o(n_101) );
in01f80 g570030 ( .a(x_out_15_3), .o(n_708) );
in01f80 g570031 ( .a(x_out_55_15), .o(n_838) );
in01f80 g570032 ( .a(x_out_36_23), .o(n_657) );
in01f80 g570033 ( .a(x_out_58_26), .o(n_621) );
in01f80 g570034 ( .a(x_out_53_19), .o(n_546) );
in01f80 g570035 ( .a(x_out_33_13), .o(n_1637) );
in01f80 g570036 ( .a(x_out_10_29), .o(n_1632) );
in01f80 g570037 ( .a(x_out_38_9), .o(n_417) );
in01f80 g570038 ( .a(x_out_26_5), .o(n_1257) );
in01f80 g570039 ( .a(x_out_31_25), .o(n_626) );
in01f80 g570040 ( .a(x_out_46_5), .o(n_133) );
in01f80 g570041 ( .a(x_out_6_15), .o(n_566) );
in01f80 g570042 ( .a(x_out_42_26), .o(n_31) );
in01f80 g570043 ( .a(x_out_17_26), .o(n_596) );
in01f80 g570044 ( .a(x_out_30_22), .o(n_1892) );
in01f80 g570045 ( .a(x_out_54_10), .o(n_561) );
in01f80 g570046 ( .a(x_out_1_21), .o(n_554) );
in01f80 g570047 ( .a(x_out_35_15), .o(n_1785) );
in01f80 g570048 ( .a(x_out_30_7), .o(n_1943) );
in01f80 g570049 ( .a(x_out_61_22), .o(n_1557) );
in01f80 g570050 ( .a(x_out_21_14), .o(n_1037) );
in01f80 g570051 ( .a(x_out_12_18), .o(n_1022) );
in01f80 g570052 ( .a(x_out_15_21), .o(n_59) );
in01f80 g570053 ( .a(x_out_55_6), .o(n_391) );
in01f80 g570054 ( .a(x_out_9_28), .o(n_603) );
in01f80 g570055 ( .a(x_out_8_25), .o(n_750) );
in01f80 g570056 ( .a(x_out_39_13), .o(n_199) );
in01f80 g570057 ( .a(x_out_1_26), .o(n_722) );
in01f80 g570058 ( .a(x_out_2_31), .o(n_343) );
in01f80 g570059 ( .a(x_out_21_7), .o(n_820) );
in01f80 g570060 ( .a(x_out_11_15), .o(n_638) );
in01f80 g570061 ( .a(x_out_61_6), .o(n_1200) );
in01f80 g570062 ( .a(x_out_40_18), .o(n_593) );
in01f80 g570063 ( .a(x_out_37_5), .o(n_1341) );
in01f80 g570064 ( .a(x_out_24_6), .o(n_1351) );
in01f80 g570065 ( .a(x_out_50_5), .o(n_569) );
in01f80 g570066 ( .a(x_out_46_18), .o(n_479) );
in01f80 g570067 ( .a(x_out_49_28), .o(n_1968) );
in01f80 g570068 ( .a(x_out_13_30), .o(n_100) );
in01f80 g570069 ( .a(x_out_15_33), .o(n_249) );
in01f80 g570070 ( .a(x_out_55_33), .o(n_1678) );
in01f80 g570071 ( .a(x_out_52_12), .o(n_1176) );
in01f80 g570072 ( .a(x_out_33_8), .o(n_1869) );
in01f80 g570073 ( .a(x_out_14_13), .o(n_941) );
in01f80 g570074 ( .a(x_out_0_4), .o(n_810) );
in01f80 g570075 ( .a(x_out_26_26), .o(n_970) );
in01f80 g570076 ( .a(x_out_12_21), .o(n_987) );
in01f80 g570077 ( .a(x_out_1_27), .o(n_1477) );
in01f80 g570078 ( .a(x_out_63_24), .o(n_1576) );
in01f80 g570079 ( .a(x_out_26_1), .o(n_1461) );
in01f80 g570080 ( .a(x_out_50_15), .o(n_741) );
in01f80 g570081 ( .a(x_out_58_20), .o(n_1636) );
in01f80 g570082 ( .a(x_out_17_13), .o(n_444) );
in01f80 g570083 ( .a(x_out_30_24), .o(n_1458) );
in01f80 g570084 ( .a(x_out_53_3), .o(n_1366) );
in01f80 g570085 ( .a(x_out_45_18), .o(n_1189) );
in01f80 g570086 ( .a(x_out_9_15), .o(n_1506) );
in01f80 g570087 ( .a(x_out_17_28), .o(n_1689) );
in01f80 g570088 ( .a(x_out_5_25), .o(n_991) );
in01f80 g570089 ( .a(x_out_11_25), .o(n_779) );
in01f80 g570090 ( .a(x_out_3_7), .o(n_667) );
in01f80 g570091 ( .a(x_out_16_25), .o(n_192) );
in01f80 g570092 ( .a(x_out_50_4), .o(n_1091) );
in01f80 g570093 ( .a(x_out_48_10), .o(n_1015) );
in01f80 g570094 ( .a(x_out_19_21), .o(n_1613) );
in01f80 g570095 ( .a(x_out_25_28), .o(n_1582) );
in01f80 g570096 ( .a(x_out_45_5), .o(n_1676) );
in01f80 g570097 ( .a(x_out_19_22), .o(n_1278) );
in01f80 g570098 ( .a(x_out_40_33), .o(n_1700) );
in01f80 g570099 ( .a(x_out_40_21), .o(n_574) );
in01f80 g570100 ( .a(x_out_29_3), .o(n_1358) );
in01f80 g570101 ( .a(x_out_13_21), .o(n_642) );
in01f80 g570102 ( .a(x_out_10_23), .o(n_1556) );
in01f80 g570103 ( .a(x_out_61_32), .o(n_799) );
in01f80 g570104 ( .a(x_out_1_32), .o(n_968) );
in01f80 g570105 ( .a(x_out_3_1), .o(n_1564) );
in01f80 g570106 ( .a(x_out_36_9), .o(n_897) );
in01f80 g570107 ( .a(x_out_34_14), .o(n_480) );
in01f80 g570108 ( .a(x_out_50_20), .o(n_191) );
in01f80 g570109 ( .a(x_out_20_4), .o(n_864) );
in01f80 g570110 ( .a(x_out_48_2), .o(n_953) );
in01f80 g570111 ( .a(x_out_24_32), .o(n_1435) );
in01f80 g570112 ( .a(x_out_29_2), .o(n_1605) );
in01f80 g570113 ( .a(x_out_38_26), .o(n_1180) );
in01f80 g570114 ( .a(x_out_33_9), .o(n_1850) );
in01f80 g570115 ( .a(x_out_14_0), .o(n_1277) );
in01f80 g570116 ( .a(x_out_57_7), .o(n_990) );
in01f80 g570117 ( .a(x_out_52_2), .o(n_1113) );
in01f80 g570118 ( .a(x_out_5_13), .o(n_1078) );
in01f80 g570119 ( .a(x_out_41_3), .o(n_1361) );
in01f80 g570120 ( .a(x_out_47_3), .o(n_1494) );
in01f80 g570121 ( .a(x_out_6_8), .o(n_508) );
in01f80 g570122 ( .a(x_out_39_26), .o(n_825) );
in01f80 g570123 ( .a(x_out_62_1), .o(n_1509) );
in01f80 g570124 ( .a(x_out_1_4), .o(n_1056) );
in01f80 g570125 ( .a(x_out_21_5), .o(n_1207) );
in01f80 g570126 ( .a(x_out_59_6), .o(n_475) );
in01f80 g570127 ( .a(x_out_19_3), .o(n_962) );
in01f80 g570128 ( .a(x_out_43_7), .o(n_1203) );
in01f80 g570129 ( .a(x_out_36_0), .o(n_195) );
in01f80 g570130 ( .a(x_out_31_0), .o(n_679) );
in01f80 g570131 ( .a(x_out_24_2), .o(n_1584) );
in01f80 g570132 ( .a(x_out_8_7), .o(n_1285) );
in01f80 g570133 ( .a(x_in_6_14), .o(n_1489) );
in01f80 g570134 ( .a(x_in_25_7), .o(n_3132) );
in01f80 g570135 ( .a(x_in_35_14), .o(n_2752) );
in01f80 g570136 ( .a(x_in_49_3), .o(n_3238) );
in01f80 g570137 ( .a(x_in_47_7), .o(n_7901) );
in01f80 g570138 ( .a(x_in_27_13), .o(n_7229) );
in01f80 g570139 ( .a(x_in_62_0), .o(n_11644) );
in01f80 g570140 ( .a(x_in_47_4), .o(n_3445) );
in01f80 g570141 ( .a(x_in_19_6), .o(n_5326) );
in01f80 g570142 ( .a(x_in_13_9), .o(n_2521) );
in01f80 g570143 ( .a(x_in_53_9), .o(n_2550) );
in01f80 g570144 ( .a(x_in_12_7), .o(n_1863) );
in01f80 g570145 ( .a(x_in_41_9), .o(n_9329) );
in01f80 g570146 ( .a(x_in_13_12), .o(n_5926) );
in01f80 g570147 ( .a(x_in_4_12), .o(n_2112) );
in01f80 g570148 ( .a(x_in_49_5), .o(n_5095) );
in01f80 g570149 ( .a(x_in_21_10), .o(n_5869) );
in01f80 g570150 ( .a(x_in_37_14), .o(n_2419) );
in01f80 g570151 ( .a(x_in_43_5), .o(n_3176) );
in01f80 g570152 ( .a(x_in_11_11), .o(n_7818) );
in01f80 g570153 ( .a(x_in_36_1), .o(n_17497) );
in01f80 g570154 ( .a(x_in_29_15), .o(n_2327) );
in01f80 g570155 ( .a(x_in_43_9), .o(n_7268) );
in01f80 g570156 ( .a(x_in_49_11), .o(n_3186) );
in01f80 g570157 ( .a(x_in_21_2), .o(n_7434) );
in01f80 g570158 ( .a(x_in_32_1), .o(n_16224) );
in01f80 g570159 ( .a(x_in_50_0), .o(n_1616) );
in01f80 g570160 ( .a(x_in_37_0), .o(n_3126) );
in01f80 g570161 ( .a(x_in_8_0), .o(n_7982) );
in01f80 g570162 ( .a(x_in_29_5), .o(n_3470) );
in01f80 g570163 ( .a(x_in_61_9), .o(n_4914) );
in01f80 g570164 ( .a(x_in_9_1), .o(n_5848) );
in01f80 g570165 ( .a(x_in_9_7), .o(n_2289) );
in01f80 g570166 ( .a(x_in_33_11), .o(n_12178) );
in01f80 g570167 ( .a(x_in_28_15), .o(n_463) );
in01f80 g570168 ( .a(x_in_51_10), .o(n_5283) );
in01f80 g570169 ( .a(x_in_43_3), .o(n_2541) );
in01f80 g570170 ( .a(x_in_24_14), .o(n_24029) );
in01f80 g570171 ( .a(x_in_39_13), .o(n_7213) );
in01f80 g570172 ( .a(x_in_55_7), .o(n_7905) );
in01f80 g570173 ( .a(x_in_4_15), .o(n_2608) );
in01f80 g570174 ( .a(x_in_53_2), .o(n_2231) );
in01f80 g570175 ( .a(x_in_35_10), .o(n_2652) );
in01f80 g570176 ( .a(x_in_51_7), .o(n_5331) );
in01f80 g570177 ( .a(x_in_35_15), .o(n_1388) );
in01f80 g570178 ( .a(x_in_11_6), .o(n_5309) );
in01f80 g570179 ( .a(x_in_25_10), .o(n_2743) );
in01f80 g570180 ( .a(x_in_25_15), .o(n_2546) );
in01f80 g570181 ( .a(x_in_17_6), .o(n_5362) );
in01f80 g570182 ( .a(x_in_17_2), .o(n_4687) );
in01f80 g570183 ( .a(x_in_5_11), .o(n_5754) );
in01f80 g570184 ( .a(x_in_41_3), .o(n_2424) );
in01f80 g570185 ( .a(x_in_49_10), .o(n_3187) );
in01f80 g570186 ( .a(x_in_5_0), .o(n_742) );
in01f80 g570187 ( .a(x_in_25_6), .o(n_3771) );
in01f80 g570188 ( .a(x_in_15_5), .o(n_4746) );
in01f80 g570189 ( .a(x_in_37_4), .o(n_2240) );
in01f80 g570190 ( .a(x_in_56_1), .o(n_13769) );
in01f80 g570191 ( .a(x_in_57_5), .o(n_4668) );
in01f80 g570192 ( .a(x_in_59_12), .o(n_4992) );
in01f80 g570193 ( .a(x_in_27_6), .o(n_5677) );
in01f80 g570194 ( .a(x_in_23_1), .o(n_2646) );
in01f80 g570195 ( .a(x_in_53_5), .o(n_2626) );
in01f80 g570196 ( .a(x_in_25_11), .o(n_3189) );
in01f80 g570197 ( .a(x_in_57_8), .o(n_2627) );
in01f80 g570198 ( .a(x_in_19_4), .o(n_5939) );
in01f80 g570199 ( .a(x_in_43_12), .o(n_7263) );
in01f80 g570200 ( .a(x_in_43_2), .o(n_2349) );
in01f80 g570201 ( .a(x_in_15_15), .o(n_5368) );
in01f80 g570202 ( .a(x_in_29_0), .o(n_491) );
in01f80 g570203 ( .a(x_in_21_14), .o(n_3043) );
in01f80 g570204 ( .a(x_in_43_14), .o(n_7311) );
in01f80 g570205 ( .a(x_in_13_3), .o(n_2516) );
in01f80 g570206 ( .a(x_in_51_1), .o(n_4932) );
in01f80 g570207 ( .a(x_in_16_1), .o(n_15444) );
in01f80 g570208 ( .a(x_in_53_11), .o(n_2870) );
in01f80 g570209 ( .a(x_in_1_6), .o(n_521) );
in01f80 g570210 ( .a(x_in_33_8), .o(n_12175) );
in01f80 g570211 ( .a(x_in_63_1), .o(n_2603) );
in01f80 g570212 ( .a(x_in_14_7), .o(n_1848) );
in01f80 g570213 ( .a(x_in_37_2), .o(n_3011) );
in01f80 g570214 ( .a(x_in_37_12), .o(n_5849) );
in01f80 g570215 ( .a(x_in_55_11), .o(n_7332) );
in01f80 g570216 ( .a(x_in_53_4), .o(n_3038) );
in01f80 g570217 ( .a(x_in_33_9), .o(n_8884) );
in01f80 g570218 ( .a(x_in_53_14), .o(n_2762) );
in01f80 g570219 ( .a(x_in_41_1), .o(n_533) );
in01f80 g570220 ( .a(x_in_38_0), .o(n_1439) );
in01f80 g570221 ( .a(x_in_61_10), .o(n_3833) );
in01f80 g570222 ( .a(x_in_48_1), .o(n_16221) );
in01f80 g570223 ( .a(x_in_21_1), .o(n_3746) );
in01f80 g570224 ( .a(x_in_57_14), .o(n_442) );
in01f80 g570225 ( .a(x_in_7_2), .o(n_2699) );
in01f80 g570226 ( .a(x_in_21_3), .o(n_6781) );
in01f80 g570227 ( .a(x_in_63_10), .o(n_11696) );
in01f80 g570228 ( .a(x_in_20_1), .o(n_17498) );
in01f80 g570229 ( .a(x_in_3_11), .o(n_6380) );
in01f80 g570230 ( .a(x_in_60_13), .o(n_27562) );
in01f80 g570231 ( .a(x_in_37_1), .o(n_4376) );
in01f80 g570232 ( .a(x_in_27_4), .o(n_5679) );
in01f80 g570233 ( .a(x_in_43_1), .o(n_2664) );
in01f80 g570234 ( .a(x_in_11_12), .o(n_5025) );
in01f80 g570235 ( .a(x_in_57_7), .o(n_4055) );
in01f80 g570236 ( .a(x_in_3_0), .o(n_2139) );
in01f80 g570237 ( .a(x_in_39_3), .o(n_2537) );
in01f80 g570238 ( .a(x_in_17_14), .o(n_4794) );
in01f80 g570239 ( .a(x_in_3_10), .o(n_5666) );
in01f80 g570240 ( .a(x_in_1_4), .o(n_247) );
in01f80 g570241 ( .a(x_in_59_14), .o(n_2422) );
in01f80 g570242 ( .a(x_in_21_7), .o(n_3036) );
in01f80 g570243 ( .a(x_in_37_10), .o(n_5745) );
in01f80 g570244 ( .a(x_in_49_8), .o(n_3188) );
in01f80 g570245 ( .a(x_in_57_13), .o(n_3560) );
in01f80 g570246 ( .a(x_in_21_0), .o(n_2066) );
in01f80 g570247 ( .a(x_in_19_11), .o(n_7765) );
in01f80 g570248 ( .a(x_in_21_4), .o(n_8557) );
in01f80 g570249 ( .a(x_in_4_0), .o(n_63) );
in01f80 g570250 ( .a(x_in_20_0), .o(n_1599) );
in01f80 g570251 ( .a(x_in_33_10), .o(n_12634) );
in01f80 g570252 ( .a(x_in_59_1), .o(n_2509) );
in01f80 g570253 ( .a(x_in_27_11), .o(n_8513) );
in01f80 g570254 ( .a(x_in_15_3), .o(n_2780) );
in01f80 g570255 ( .a(x_in_59_4), .o(n_5271) );
in01f80 g570256 ( .a(x_in_63_9), .o(n_10916) );
in01f80 g570257 ( .a(x_in_37_7), .o(n_3318) );
in01f80 g570258 ( .a(x_in_1_12), .o(n_1808) );
in01f80 g570259 ( .a(x_in_23_2), .o(n_5430) );
in01f80 g570260 ( .a(x_in_45_13), .o(n_7216) );
in01f80 g570261 ( .a(x_in_24_15), .o(n_2545) );
in01f80 g570262 ( .a(x_in_53_12), .o(n_2548) );
in01f80 g570263 ( .a(x_in_25_14), .o(n_2492) );
in01f80 g570264 ( .a(x_in_51_11), .o(n_8420) );
in01f80 g570265 ( .a(x_in_23_9), .o(n_10918) );
in01f80 g570266 ( .a(x_in_3_7), .o(n_5757) );
in01f80 g570267 ( .a(x_in_39_9), .o(n_4514) );
in01f80 g570268 ( .a(x_in_41_7), .o(n_9327) );
in01f80 g570269 ( .a(x_in_61_12), .o(n_2353) );
in01f80 g570270 ( .a(x_in_63_11), .o(n_7308) );
in01f80 g570271 ( .a(x_in_60_0), .o(n_16010) );
in01f80 g570272 ( .a(x_in_19_13), .o(n_5556) );
in01f80 g570273 ( .a(x_in_51_2), .o(n_2490) );
in01f80 g570274 ( .a(x_in_35_9), .o(n_5098) );
in01f80 g570275 ( .a(x_in_45_3), .o(n_2439) );
in01f80 g570276 ( .a(x_in_28_1), .o(n_8438) );
in01f80 g570277 ( .a(x_in_55_8), .o(n_7315) );
in01f80 g570278 ( .a(x_in_19_3), .o(n_5252) );
in01f80 g570279 ( .a(x_in_59_15), .o(n_4409) );
in01f80 g570280 ( .a(x_in_63_3), .o(n_2828) );
in01f80 g570281 ( .a(x_in_37_3), .o(n_4654) );
in01f80 g570282 ( .a(x_in_47_5), .o(n_4737) );
in01f80 g570283 ( .a(x_in_55_9), .o(n_10915) );
in01f80 g570284 ( .a(x_in_31_11), .o(n_7298) );
in01f80 g570285 ( .a(x_in_56_15), .o(n_818) );
in01f80 g570286 ( .a(x_in_23_13), .o(n_6488) );
in01f80 g570287 ( .a(x_in_41_8), .o(n_9612) );
in01f80 g570288 ( .a(x_in_11_5), .o(n_2430) );
in01f80 g570289 ( .a(x_in_33_3), .o(n_2329) );
in01f80 g570290 ( .a(x_in_55_14), .o(n_16156) );
in01f80 g570291 ( .a(x_in_35_13), .o(n_5245) );
in01f80 g570292 ( .a(x_in_49_1), .o(n_448) );
in01f80 g570293 ( .a(x_in_51_14), .o(n_2269) );
in01f80 g570294 ( .a(x_in_5_9), .o(n_6000) );
in01f80 g570295 ( .a(x_in_51_4), .o(n_5979) );
in01f80 g570296 ( .a(x_in_25_8), .o(n_3129) );
in01f80 g570297 ( .a(x_in_56_0), .o(n_20) );
in01f80 g570298 ( .a(x_in_11_8), .o(n_5352) );
in01f80 g570299 ( .a(x_in_29_3), .o(n_3591) );
in01f80 g570300 ( .a(x_in_6_1), .o(n_16928) );
in01f80 g570301 ( .a(x_in_12_0), .o(n_11650) );
in01f80 g570302 ( .a(x_in_53_13), .o(n_5988) );
in01f80 g570303 ( .a(x_in_8_1), .o(n_12312) );
in01f80 g570304 ( .a(x_in_47_12), .o(n_7247) );
in01f80 g570305 ( .a(x_in_12_1), .o(n_15678) );
in01f80 g570306 ( .a(x_in_47_2), .o(n_5365) );
in01f80 g570307 ( .a(x_in_54_0), .o(n_738) );
in01f80 g570308 ( .a(x_in_45_12), .o(n_10486) );
in01f80 g570309 ( .a(x_in_51_5), .o(n_3792) );
in01f80 g570310 ( .a(x_in_47_10), .o(n_11034) );
in01f80 g570311 ( .a(x_in_41_4), .o(n_5381) );
in01f80 g570312 ( .a(x_in_57_3), .o(n_2526) );
in01f80 g570313 ( .a(x_in_49_12), .o(n_2737) );
in01f80 g570314 ( .a(x_in_52_13), .o(n_280) );
in01f80 g570315 ( .a(x_in_53_10), .o(n_2653) );
in01f80 g570316 ( .a(x_in_9_13), .o(n_6726) );
in01f80 g570317 ( .a(x_in_23_11), .o(n_7296) );
in01f80 g570318 ( .a(x_in_31_15), .o(n_5355) );
in01f80 g570319 ( .a(x_in_43_8), .o(n_5501) );
in01f80 g570320 ( .a(x_in_45_9), .o(n_2428) );
in01f80 g570321 ( .a(x_in_21_11), .o(n_5872) );
in01f80 g570322 ( .a(x_in_7_8), .o(n_7304) );
in01f80 g570323 ( .a(x_in_57_2), .o(n_2222) );
in01f80 g570324 ( .a(x_in_39_1), .o(n_2607) );
in01f80 g570325 ( .a(x_in_7_12), .o(n_7340) );
in01f80 g570326 ( .a(x_in_51_9), .o(n_5332) );
in01f80 g570327 ( .a(x_in_27_10), .o(n_7417) );
in01f80 g570328 ( .a(x_in_17_5), .o(n_9646) );
in01f80 g570329 ( .a(x_in_61_11), .o(n_4529) );
in01f80 g570330 ( .a(x_in_25_12), .o(n_5317) );
in01f80 g570331 ( .a(x_in_59_3), .o(n_3260) );
in01f80 g570332 ( .a(x_in_52_14), .o(n_616) );
in01f80 g570333 ( .a(x_in_24_1), .o(n_12572) );
in01f80 g570334 ( .a(x_in_53_7), .o(n_2525) );
in01f80 g570335 ( .a(x_in_17_11), .o(n_5418) );
in01f80 g570336 ( .a(x_in_19_5), .o(n_3174) );
in01f80 g570337 ( .a(x_in_32_7), .o(n_22508) );
in01f80 g570338 ( .a(x_in_31_7), .o(n_7902) );
in01f80 g570339 ( .a(x_in_25_13), .o(n_5311) );
in01f80 g570340 ( .a(x_in_25_3), .o(n_5703) );
in01f80 g570341 ( .a(x_in_17_13), .o(n_10477) );
in01f80 g570342 ( .a(x_in_27_2), .o(n_2478) );
in01f80 g570343 ( .a(x_in_27_8), .o(n_7287) );
in01f80 g570344 ( .a(x_in_5_10), .o(n_5388) );
in01f80 g570345 ( .a(x_in_33_12), .o(n_12635) );
in01f80 g570346 ( .a(x_in_37_13), .o(n_4343) );
in01f80 g570347 ( .a(x_in_61_8), .o(n_4937) );
in01f80 g570348 ( .a(x_in_26_1), .o(n_16007) );
in01f80 g570349 ( .a(x_in_3_12), .o(n_5247) );
in01f80 g570350 ( .a(x_in_29_9), .o(n_2597) );
in01f80 g570351 ( .a(x_in_11_1), .o(n_2365) );
in01f80 g570352 ( .a(x_in_9_12), .o(n_8957) );
in01f80 g570353 ( .a(x_in_63_14), .o(n_2606) );
in01f80 g570354 ( .a(x_in_31_2), .o(n_5373) );
in01f80 g570355 ( .a(x_in_63_12), .o(n_8206) );
in01f80 g570356 ( .a(x_in_9_14), .o(n_2376) );
in01f80 g570357 ( .a(x_in_47_8), .o(n_7241) );
in01f80 g570358 ( .a(x_in_61_6), .o(n_5761) );
in01f80 g570359 ( .a(x_in_61_15), .o(n_2655) );
in01f80 g570360 ( .a(x_in_55_1), .o(n_2618) );
in01f80 g570361 ( .a(x_in_51_3), .o(n_5180) );
in01f80 g570362 ( .a(x_in_17_10), .o(n_5359) );
in01f80 g570363 ( .a(x_in_22_0), .o(n_1511) );
in01f80 g570364 ( .a(x_in_27_9), .o(n_7289) );
in01f80 g570365 ( .a(x_in_13_13), .o(n_2834) );
in01f80 g570366 ( .a(x_in_17_8), .o(n_5360) );
in01f80 g570367 ( .a(x_in_39_12), .o(n_2036) );
in01f80 g570368 ( .a(x_in_3_13), .o(n_6746) );
in01f80 g570369 ( .a(x_in_17_3), .o(n_2520) );
in01f80 g570370 ( .a(x_in_19_0), .o(n_2039) );
in01f80 g570371 ( .a(x_in_43_4), .o(n_5293) );
in01f80 g570372 ( .a(x_in_2_1), .o(n_16026) );
in01f80 g570373 ( .a(x_in_33_4), .o(n_5281) );
in01f80 g570374 ( .a(x_in_45_6), .o(n_2513) );
in01f80 g570375 ( .a(x_in_55_12), .o(n_7278) );
in01f80 g570376 ( .a(x_in_40_0), .o(n_1790) );
in01f80 g570377 ( .a(x_in_29_2), .o(n_4592) );
in01f80 g570378 ( .a(x_in_50_15), .o(n_2) );
in01f80 g570379 ( .a(x_in_34_1), .o(n_16351) );
in01f80 g570380 ( .a(x_in_5_5), .o(n_5296) );
in01f80 g570381 ( .a(x_in_63_4), .o(n_3737) );
in01f80 g570382 ( .a(x_in_55_4), .o(n_3742) );
in01f80 g570383 ( .a(x_in_17_12), .o(n_5415) );
in01f80 g570384 ( .a(x_in_3_1), .o(n_4419) );
in01f80 g570385 ( .a(x_in_9_9), .o(n_2248) );
in01f80 g570386 ( .a(x_in_13_6), .o(n_2506) );
in01f80 g570387 ( .a(x_in_59_7), .o(n_5699) );
in01f80 g570388 ( .a(x_in_11_3), .o(n_2431) );
in01f80 g570389 ( .a(x_in_13_11), .o(n_482) );
in01f80 g570390 ( .a(x_in_18_0), .o(n_503) );
in01f80 g570391 ( .a(x_in_1_0), .o(n_2235) );
in01f80 g570392 ( .a(x_in_4_1), .o(n_2567) );
in01f80 g570393 ( .a(x_in_22_1), .o(n_15720) );
in01f80 g570394 ( .a(x_in_39_5), .o(n_4338) );
in01f80 g570395 ( .a(x_in_35_12), .o(n_5032) );
in01f80 g570396 ( .a(x_in_52_7), .o(n_22222) );
in01f80 g570397 ( .a(x_in_59_5), .o(n_3259) );
in01f80 g570398 ( .a(x_in_2_0), .o(n_884) );
in01f80 g570399 ( .a(x_in_29_12), .o(n_1164) );
in01f80 g570400 ( .a(x_in_59_11), .o(n_8482) );
in01f80 g570401 ( .a(x_in_24_0), .o(n_1300) );
in01f80 g570402 ( .a(x_in_23_10), .o(n_11041) );
in01f80 g570403 ( .a(x_in_5_3), .o(n_2540) );
in01f80 g570404 ( .a(x_in_45_5), .o(n_2438) );
in01f80 g570405 ( .a(x_in_23_6), .o(n_6689) );
in01f80 g570406 ( .a(x_in_14_0), .o(n_900) );
in01f80 g570407 ( .a(x_in_49_4), .o(n_2234) );
in01f80 g570408 ( .a(x_in_7_5), .o(n_5256) );
in01f80 g570409 ( .a(x_in_19_2), .o(n_2440) );
in01f80 g570410 ( .a(x_in_29_6), .o(n_3390) );
in01f80 g570411 ( .a(x_in_27_3), .o(n_2421) );
in01f80 g570412 ( .a(x_in_7_7), .o(n_6494) );
in01f80 g570413 ( .a(x_in_31_3), .o(n_2721) );
in01f80 g570414 ( .a(x_in_45_10), .o(n_2134) );
in01f80 g570415 ( .a(x_in_61_0), .o(n_2605) );
in01f80 g570416 ( .a(x_in_39_8), .o(n_8133) );
in01f80 g570417 ( .a(x_in_32_13), .o(n_27151) );
in01f80 g570418 ( .a(x_in_5_7), .o(n_2645) );
in01f80 g570419 ( .a(x_in_37_15), .o(n_3241) );
in01f80 g570420 ( .a(x_in_1_8), .o(n_1072) );
in01f80 g570421 ( .a(x_in_41_12), .o(n_9608) );
in01f80 g570422 ( .a(x_in_3_15), .o(n_123) );
in01f80 g570423 ( .a(x_in_19_10), .o(n_3020) );
in01f80 g570424 ( .a(x_in_61_14), .o(n_4847) );
in01f80 g570425 ( .a(x_in_57_10), .o(n_3409) );
in01f80 g570426 ( .a(x_in_35_6), .o(n_5369) );
in01f80 g570427 ( .a(x_in_51_6), .o(n_6350) );
in01f80 g570428 ( .a(x_in_23_5), .o(n_4744) );
in01f80 g570429 ( .a(x_in_61_2), .o(n_4143) );
in01f80 g570430 ( .a(x_in_63_5), .o(n_4745) );
in01f80 g570431 ( .a(x_in_51_15), .o(n_558) );
in01f80 g570432 ( .a(x_in_45_14), .o(n_2326) );
in01f80 g570433 ( .a(x_in_45_8), .o(n_2527) );
in01f80 g570434 ( .a(x_in_20_15), .o(n_1140) );
in01f80 g570435 ( .a(x_in_15_2), .o(n_4946) );
in01f80 g570436 ( .a(x_in_59_2), .o(n_2445) );
in01f80 g570437 ( .a(x_in_15_1), .o(n_2593) );
in01f80 g570438 ( .a(x_in_45_15), .o(n_1720) );
in01f80 g570439 ( .a(x_in_21_13), .o(n_2310) );
in01f80 g570440 ( .a(x_in_29_1), .o(n_2409) );
in01f80 g570441 ( .a(x_in_33_15), .o(n_2538) );
in01f80 g570442 ( .a(x_in_39_14), .o(n_2343) );
in01f80 g570443 ( .a(x_in_45_7), .o(n_2528) );
in01f80 g570444 ( .a(x_in_62_1), .o(n_16012) );
in01f80 g570445 ( .a(x_in_52_0), .o(n_119) );
in01f80 g570446 ( .a(x_in_42_0), .o(n_1903) );
in01f80 g570447 ( .a(x_in_46_1), .o(n_15810) );
in01f80 g570448 ( .a(x_in_15_8), .o(n_6492) );
in01f80 g570449 ( .a(x_in_11_13), .o(n_2681) );
in01f80 g570450 ( .a(x_in_15_10), .o(n_11037) );
in01f80 g570451 ( .a(x_in_58_0), .o(n_13729) );
in01f80 g570452 ( .a(x_in_1_10), .o(n_260) );
in01f80 g570453 ( .a(x_in_5_4), .o(n_2517) );
in01f80 g570454 ( .a(x_in_51_0), .o(n_610) );
in01f80 g570455 ( .a(x_in_13_5), .o(n_2505) );
in01f80 g570456 ( .a(x_in_59_9), .o(n_2363) );
in01f80 g570457 ( .a(x_in_15_6), .o(n_6687) );
in01f80 g570458 ( .a(x_in_17_0), .o(n_1) );
in01f80 g570459 ( .a(x_in_24_2), .o(n_13487) );
in01f80 g570460 ( .a(x_in_33_2), .o(n_2451) );
in01f80 g570461 ( .a(x_in_23_4), .o(n_3744) );
in01f80 g570462 ( .a(x_in_57_9), .o(n_3245) );
in01f80 g570463 ( .a(x_in_53_6), .o(n_2651) );
in01f80 g570464 ( .a(x_in_5_13), .o(n_13241) );
in01f80 g570465 ( .a(x_in_43_15), .o(n_2394) );
in01f80 g570466 ( .a(x_in_45_2), .o(n_5986) );
in01f80 g570467 ( .a(x_in_57_4), .o(n_2601) );
in01f80 g570468 ( .a(x_in_31_4), .o(n_3739) );
in01f80 g570469 ( .a(x_in_39_2), .o(n_2037) );
in01f80 g570470 ( .a(x_in_31_10), .o(n_11698) );
in01f80 g570471 ( .a(x_in_31_13), .o(n_7291) );
in01f80 g570472 ( .a(x_in_58_1), .o(n_15723) );
in01f80 g570473 ( .a(FE_OFN37_n_17184), .o(n_15183) );
in01f80 g570474 ( .a(n_17184), .o(n_13676) );
in01f80 g570476 ( .a(FE_OFN1115_rst), .o(n_28682) );
in01f80 g570477 ( .a(FE_OFN1115_rst), .o(n_28597) );
in01f80 g570484 ( .a(FE_OFN1115_rst), .o(n_17184) );
in01f80 g570513 ( .a(FE_OFN1108_rst), .o(n_26609) );
in01f80 g570521 ( .a(n_26609), .o(n_29617) );
in01f80 g570522 ( .a(n_26609), .o(n_27452) );
in01f80 g570527 ( .a(n_26609), .o(n_29204) );
in01f80 g570528 ( .a(n_26609), .o(n_29068) );
in01f80 g570549 ( .a(n_2022), .o(n_16289) );
in01f80 g570550 ( .a(n_2022), .o(n_16909) );
in01f80 g570596 ( .a(n_16909), .o(n_28303) );
in01f80 g570598 ( .a(FE_OFN1115_rst), .o(n_2022) );
in01f80 g570602 ( .a(FE_OFN349_n_4860), .o(n_16028) );
in01f80 g570603 ( .a(FE_OFN324_n_4860), .o(n_16893) );
in01f80 g570605 ( .a(FE_OFN347_n_4860), .o(n_16656) );
in01f80 g570610 ( .a(FE_OFN349_n_4860), .o(n_27400) );
in01f80 g570638 ( .a(n_26312), .o(n_27012) );
in01f80 g570735 ( .a(n_26312), .o(n_27449) );
in01f80 g570736 ( .a(n_5003), .o(n_29264) );
in01f80 g570737 ( .a(FE_OFN1162_n_5003), .o(n_25680) );
in01f80 g570745 ( .a(FE_OFN1162_n_5003), .o(n_27709) );
in01f80 g570746 ( .a(n_5003), .o(n_29261) );
in01f80 g570754 ( .a(n_5003), .o(n_29104) );
in01f80 g570755 ( .a(n_5003), .o(n_28928) );
in01f80 g570773 ( .a(n_5003), .o(n_28607) );
in01f80 g570774 ( .a(n_5003), .o(n_28362) );
in01f80 g570775 ( .a(n_4860), .o(n_5003) );
in01f80 g570791 ( .a(FE_OFN331_n_4860), .o(n_28771) );
in01f80 g570797 ( .a(FE_OFN324_n_4860), .o(n_29269) );
in01f80 g570800 ( .a(FE_OFN349_n_4860), .o(n_27681) );
in01f80 g570803 ( .a(FE_OFN349_n_4860), .o(n_22615) );
in01f80 g570806 ( .a(FE_OFN349_n_4860), .o(n_29687) );
in01f80 g570807 ( .a(FE_OFN329_n_4860), .o(n_26454) );
in01f80 g570809 ( .a(FE_OFN349_n_4860), .o(n_23315) );
in01f80 g570810 ( .a(n_4860), .o(n_26184) );
in01f80 g570813 ( .a(FE_OFN349_n_4860), .o(n_29496) );
in01f80 g570818 ( .a(n_4860), .o(n_4162) );
in01f80 g570821 ( .a(FE_OFN331_n_4860), .o(n_4280) );
in01f80 g570841 ( .a(FE_OFN303_n_3069), .o(n_29266) );
in01f80 g570847 ( .a(n_4276), .o(n_29046) );
in01f80 g570848 ( .a(n_4276), .o(n_29683) );
in01f80 g570849 ( .a(FE_OFN293_n_3069), .o(n_4276) );
in01f80 g570853 ( .a(n_4276), .o(n_29691) );
in01f80 g570854 ( .a(n_4276), .o(n_29698) );
in01f80 g570856 ( .a(n_4276), .o(n_27933) );
in01f80 g570857 ( .a(n_4276), .o(n_23813) );
in01f80 g570910 ( .a(FE_OFN293_n_3069), .o(n_27194) );
in01f80 g570912 ( .a(n_4270), .o(n_21076) );
in01f80 g570916 ( .a(FE_OFN292_n_3069), .o(n_4270) );
in01f80 g570917 ( .a(n_4270), .o(n_29033) );
in01f80 g570919 ( .a(n_4270), .o(n_29664) );
in01f80 g570920 ( .a(n_4270), .o(n_21988) );
in01f80 g570927 ( .a(n_4270), .o(n_28608) );
in01f80 g570930 ( .a(n_4270), .o(n_22019) );
in01f80 g570932 ( .a(n_4270), .o(n_23291) );
in01f80 g570933 ( .a(n_4270), .o(n_22960) );
in01f80 g570943 ( .a(n_26312), .o(n_4860) );
in01f80 g570944 ( .a(FE_OFN1118_rst), .o(n_26312) );
in01f80 g570945 ( .a(x_in_36_0), .o(n_1914) );
in01f80 g570946 ( .a(x_in_7_3), .o(n_5272) );
in01f80 g570947 ( .a(x_in_7_11), .o(n_7336) );
in01f80 g570948 ( .a(x_in_39_10), .o(n_8851) );
in01f80 g570949 ( .a(x_in_4_14), .o(n_2403) );
in01f80 g570950 ( .a(x_in_49_13), .o(n_2691) );
in01f80 g570951 ( .a(x_in_5_8), .o(n_5291) );
in01f80 g570952 ( .a(x_in_20_13), .o(n_28222) );
in01f80 g570953 ( .a(x_in_27_1), .o(n_2420) );
in01f80 g570954 ( .a(x_in_48_0), .o(n_1810) );
in01f80 g570955 ( .a(x_in_30_0), .o(n_11647) );
in01f80 g570956 ( .a(x_in_40_1), .o(n_16438) );
in01f80 g570957 ( .a(x_in_37_6), .o(n_5884) );
in01f80 g570958 ( .a(x_in_2_15), .o(n_1029) );
in01f80 g570959 ( .a(x_in_27_14), .o(n_14997) );
in01f80 g570960 ( .a(x_in_55_6), .o(n_6685) );
in01f80 g570961 ( .a(x_in_19_14), .o(n_4057) );
in01f80 g570962 ( .a(x_in_29_13), .o(n_1250) );
in01f80 g570963 ( .a(x_in_41_13), .o(n_2214) );
in01f80 g570964 ( .a(x_in_49_9), .o(n_3191) );
in01f80 g570965 ( .a(x_in_42_1), .o(n_15877) );
in01f80 g570966 ( .a(x_in_3_2), .o(n_2272) );
in01f80 g570967 ( .a(x_in_41_14), .o(n_8032) );
in01f80 g570968 ( .a(x_in_11_14), .o(n_2124) );
in01f80 g570969 ( .a(x_in_16_0), .o(n_844) );
in01f80 g570970 ( .a(x_in_35_2), .o(n_2061) );
in01f80 g570971 ( .a(x_in_29_14), .o(n_3736) );
in01f80 g570972 ( .a(x_in_37_8), .o(n_5881) );
in01f80 g570973 ( .a(x_in_31_12), .o(n_6753) );
in01f80 g570974 ( .a(x_in_47_6), .o(n_6683) );
in01f80 g570975 ( .a(x_in_13_7), .o(n_2657) );
in01f80 g570976 ( .a(x_in_25_1), .o(n_289) );
in01f80 g570977 ( .a(x_in_59_10), .o(n_2668) );
in01f80 g570978 ( .a(x_in_19_1), .o(n_3763) );
in01f80 g570979 ( .a(x_in_15_14), .o(n_2574) );
in01f80 g570980 ( .a(x_in_54_1), .o(n_15717) );
in01f80 g570981 ( .a(x_in_46_0), .o(n_11653) );
in01f80 g570982 ( .a(x_in_47_15), .o(n_5363) );
in01f80 g570983 ( .a(x_in_35_3), .o(n_5390) );
in01f80 g570984 ( .a(x_in_23_14), .o(n_16158) );
in01f80 g570985 ( .a(x_in_25_0), .o(n_1021) );
in01f80 g570986 ( .a(x_in_41_6), .o(n_9610) );
in01f80 g570987 ( .a(x_in_1_14), .o(n_892) );
in01f80 g570988 ( .a(x_in_37_11), .o(n_4180) );
in01f80 g570989 ( .a(x_in_13_10), .o(n_2673) );
in01f80 g570990 ( .a(x_in_7_10), .o(n_8165) );
in01f80 g570991 ( .a(x_in_0_1), .o(n_2434) );
in01f80 g570992 ( .a(x_in_33_5), .o(n_11297) );
in01f80 g570993 ( .a(x_in_19_12), .o(n_5244) );
in01f80 g570994 ( .a(x_in_15_9), .o(n_10917) );
in01f80 g570995 ( .a(x_in_44_0), .o(n_11640) );
in01f80 g570996 ( .a(x_in_55_15), .o(n_5376) );
in01f80 g570997 ( .a(x_in_5_15), .o(n_23944) );
in01f80 g570998 ( .a(x_in_55_10), .o(n_11040) );
in01f80 g570999 ( .a(x_in_9_15), .o(n_2643) );
in01f80 g571000 ( .a(x_in_3_3), .o(n_5825) );
in01f80 g571001 ( .a(x_in_51_13), .o(n_5689) );
in01f80 g571002 ( .a(x_in_29_7), .o(n_3035) );
in01f80 g571003 ( .a(x_in_55_3), .o(n_3079) );
in01f80 g571004 ( .a(x_in_47_13), .o(n_2448) );
in01f80 g571005 ( .a(x_in_61_3), .o(n_3608) );
in01f80 g571006 ( .a(x_in_19_8), .o(n_5554) );
in01f80 g571007 ( .a(x_in_41_2), .o(n_5435) );
in01f80 g571008 ( .a(x_in_56_12), .o(n_246) );
in01f80 g571009 ( .a(x_in_3_5), .o(n_5963) );
in01f80 g571010 ( .a(x_in_21_15), .o(n_2309) );
in01f80 g571011 ( .a(x_in_53_1), .o(n_4825) );
in01f80 g571012 ( .a(x_in_11_4), .o(n_5387) );
in01f80 g571013 ( .a(x_in_55_2), .o(n_5336) );
in01f80 g571014 ( .a(x_in_33_7), .o(n_8885) );
in01f80 g571015 ( .a(x_in_23_3), .o(n_3075) );
in01f80 g571016 ( .a(x_in_47_9), .o(n_10913) );
in01f80 g571017 ( .a(x_in_55_13), .o(n_7231) );
in01f80 g571018 ( .a(x_in_21_6), .o(n_5914) );
in01f80 g571019 ( .a(x_in_10_1), .o(n_15988) );
in01f80 g571020 ( .a(x_in_28_0), .o(n_1449) );
in01f80 g571021 ( .a(x_in_60_1), .o(n_17191) );
in01f80 g571022 ( .a(x_in_17_7), .o(n_9651) );
in01f80 g571023 ( .a(x_in_6_7), .o(n_467) );
in01f80 g571024 ( .a(x_in_35_8), .o(n_4939) );
in01f80 g571025 ( .a(x_in_29_11), .o(n_2875) );
in01f80 g571026 ( .a(x_in_47_3), .o(n_2747) );
in01f80 g571027 ( .a(x_in_25_5), .o(n_4593) );
in01f80 g571028 ( .a(x_in_19_7), .o(n_5940) );
in01f80 g571029 ( .a(x_in_13_14), .o(n_3077) );
in01f80 g571030 ( .a(x_in_0_0), .o(n_699) );
in01f80 g571031 ( .a(x_in_4_11), .o(n_1168) );
in01f80 g571032 ( .a(x_in_33_6), .o(n_12172) );
in01f80 g571033 ( .a(x_in_47_11), .o(n_7245) );
in01f80 g571034 ( .a(x_in_49_15), .o(n_1624) );
in01f80 g571035 ( .a(x_in_39_11), .o(n_7317) );
in01f80 g571036 ( .a(x_in_3_4), .o(n_5931) );
in01f80 g571037 ( .a(x_in_13_15), .o(n_2354) );
in01f80 g571038 ( .a(x_in_11_2), .o(n_2332) );
in01f80 g571039 ( .a(x_in_11_7), .o(n_5089) );
in01f80 g571040 ( .a(x_in_10_0), .o(n_373) );
in01f80 g571041 ( .a(x_in_7_1), .o(n_2408) );
in01f80 g571042 ( .a(x_in_61_13), .o(n_2518) );
in01f80 g571043 ( .a(x_in_13_8), .o(n_2522) );
in01f80 g571044 ( .a(x_in_27_5), .o(n_3747) );
in01f80 g571045 ( .a(x_in_55_5), .o(n_4329) );
in01f80 g571046 ( .a(x_in_33_14), .o(n_2052) );
in01f80 g571047 ( .a(x_in_31_8), .o(n_8200) );
in01f80 g571048 ( .a(x_in_23_7), .o(n_7906) );
in01f80 g571049 ( .a(x_in_27_15), .o(n_2536) );
in01f80 g571050 ( .a(x_in_31_9), .o(n_10914) );
in01f80 g571051 ( .a(x_in_21_12), .o(n_5977) );
in01f80 g571052 ( .a(x_in_34_15), .o(n_1125) );
in01f80 g571053 ( .a(x_in_49_2), .o(n_1913) );
in01f80 g571054 ( .a(x_in_51_12), .o(n_6420) );
in01f80 g571055 ( .a(x_in_45_11), .o(n_2049) );
in01f80 g571056 ( .a(x_in_63_13), .o(n_2523) );
in01f80 g571057 ( .a(x_in_15_12), .o(n_7338) );
in01f80 g571058 ( .a(x_in_45_4), .o(n_2442) );
in01f80 g571059 ( .a(x_in_36_7), .o(n_22395) );
in01f80 g571060 ( .a(x_in_30_1), .o(n_16013) );
in01f80 g571061 ( .a(x_in_39_6), .o(n_6500) );
in01f80 g571062 ( .a(x_in_17_1), .o(n_3363) );
in01f80 g571063 ( .a(x_in_29_4), .o(n_3724) );
in01f80 g571064 ( .a(x_in_57_15), .o(n_3641) );
in01f80 g571065 ( .a(x_in_59_6), .o(n_5275) );
in01f80 g571066 ( .a(x_in_63_8), .o(n_7272) );
in01f80 g571067 ( .a(x_in_47_14), .o(n_2558) );
in01f80 g571068 ( .a(x_in_13_4), .o(n_2433) );
in01f80 g571069 ( .a(x_in_48_13), .o(n_27547) );
in01f80 g571070 ( .a(x_in_9_6), .o(n_2230) );
in01f80 g571071 ( .a(x_in_49_6), .o(n_2588) );
in01f80 g571072 ( .a(x_in_17_9), .o(n_9654) );
in01f80 g571073 ( .a(x_in_57_6), .o(n_2512) );
in01f80 g571074 ( .a(x_in_15_11), .o(n_7334) );
in01f80 g571075 ( .a(x_in_39_4), .o(n_3107) );
in01f80 g571076 ( .a(x_in_36_14), .o(n_29194) );
in01f80 g571077 ( .a(x_in_5_6), .o(n_3568) );
in01f80 g571078 ( .a(x_in_53_0), .o(n_4042) );
in01f80 g571079 ( .a(x_in_43_7), .o(n_5519) );
in01f80 g571080 ( .a(x_in_44_1), .o(n_15992) );
in01f80 g571081 ( .a(x_in_7_15), .o(n_2624) );
in01f80 g571082 ( .a(x_in_61_4), .o(n_8929) );
in01f80 g571083 ( .a(x_in_7_14), .o(n_15590) );
in01f80 g571084 ( .a(x_in_51_8), .o(n_6351) );
in01f80 g571085 ( .a(x_in_43_6), .o(n_5327) );
in01f80 g571086 ( .a(x_in_41_0), .o(n_2534) );
in01f80 g571087 ( .a(x_in_61_1), .o(n_3237) );
in01f80 g571088 ( .a(x_in_26_0), .o(n_497) );
in01f80 g571089 ( .a(x_in_49_7), .o(n_2589) );
in01f80 g571090 ( .a(x_in_7_4), .o(n_8522) );
in01f80 g571091 ( .a(x_in_7_13), .o(n_7285) );
in01f80 g571092 ( .a(x_in_25_9), .o(n_2581) );
in01f80 g571093 ( .a(x_in_31_5), .o(n_4738) );
in01f80 g571094 ( .a(x_in_36_15), .o(n_27230) );
in01f80 g571095 ( .a(x_in_35_11), .o(n_8524) );
in01f80 g571096 ( .a(x_in_41_5), .o(n_2583) );
in01f80 g571097 ( .a(x_in_8_15), .o(n_1942) );
in01f80 g571098 ( .a(x_in_9_4), .o(n_1480) );
in01f80 g571099 ( .a(x_in_7_9), .o(n_7320) );
in01f80 g571100 ( .a(x_in_45_1), .o(n_2385) );
in01f80 g571101 ( .a(x_in_41_11), .o(n_11409) );
in01f80 g571102 ( .a(x_in_27_7), .o(n_5680) );
in01f80 g571103 ( .a(x_in_23_15), .o(n_5371) );
in01f80 g571104 ( .a(x_in_59_13), .o(n_2635) );
in01f80 g571105 ( .a(x_in_43_11), .o(n_8443) );
in01f80 g571106 ( .a(x_in_3_9), .o(n_5905) );
in01f80 g571107 ( .a(x_in_34_0), .o(n_1266) );
in01f80 g571108 ( .a(x_in_5_12), .o(n_5888) );
in01f80 g571109 ( .a(x_in_35_4), .o(n_5987) );
in01f80 g571110 ( .a(x_in_33_13), .o(n_2533) );
in01f80 g571111 ( .a(x_in_38_1), .o(n_8847) );
in01f80 g571112 ( .a(x_in_4_13), .o(n_96) );
in01f80 g571113 ( .a(x_in_9_11), .o(n_2488) );
in01f80 g571114 ( .a(x_in_63_6), .o(n_6711) );
in01f80 g571115 ( .a(x_in_32_0), .o(n_1705) );
in01f80 g571116 ( .a(x_in_9_8), .o(n_2060) );
in01f80 g571117 ( .a(x_in_5_2), .o(n_2413) );
in01f80 g571118 ( .a(x_in_9_2), .o(n_5216) );
in01f80 g571119 ( .a(x_in_59_8), .o(n_5691) );
in01f80 g571120 ( .a(x_in_15_4), .o(n_3482) );
in01f80 g571121 ( .a(x_in_39_7), .o(n_7325) );
in01f80 g571122 ( .a(x_in_61_5), .o(n_5242) );
in01f80 g571123 ( .a(x_in_49_14), .o(n_9118) );
in01f80 g571124 ( .a(x_in_33_0), .o(n_2636) );
in01f80 g571125 ( .a(x_in_35_7), .o(n_4942) );
in01f80 g571126 ( .a(x_in_23_12), .o(n_7323) );
in01f80 g571127 ( .a(x_in_29_8), .o(n_2864) );
in01f80 g571128 ( .a(x_in_29_10), .o(n_8537) );
in01f80 g571129 ( .a(x_in_6_0), .o(n_784) );
in01f80 g571130 ( .a(x_in_3_14), .o(n_2317) );
in01f80 g571131 ( .a(x_in_31_14), .o(n_16154) );
in01f80 g571132 ( .a(x_in_19_9), .o(n_5537) );
in01f80 g571133 ( .a(x_in_53_15), .o(n_3193) );
in01f80 g571134 ( .a(x_in_11_10), .o(n_3229) );
in01f80 g571135 ( .a(x_in_31_6), .o(n_6483) );
in01f80 g571136 ( .a(x_in_35_1), .o(n_5156) );
in01f80 g571137 ( .a(x_in_35_5), .o(n_2377) );
in01f80 g571138 ( .a(x_in_3_6), .o(n_5515) );
in01f80 g571139 ( .a(x_in_23_8), .o(n_7270) );
in01f80 g571140 ( .a(x_in_14_1), .o(n_15724) );
in01f80 g571141 ( .a(x_in_37_5), .o(n_5742) );
in01f80 g571142 ( .a(x_in_63_15), .o(n_5042) );
in01f80 g571143 ( .a(x_in_9_10), .o(n_2285) );
in01f80 g571144 ( .a(x_in_15_13), .o(n_2575) );
in01f80 g571145 ( .a(x_in_27_12), .o(n_7402) );
in01f80 g571146 ( .a(x_in_37_9), .o(n_5962) );
in01f80 g571147 ( .a(x_in_31_1), .o(n_2660) );
in01f80 g571148 ( .a(x_in_61_7), .o(n_5839) );
in01f80 g571149 ( .a(x_in_21_8), .o(n_5860) );
in01f80 g571150 ( .a(x_in_1_1), .o(n_2395) );
in01f80 g571151 ( .a(x_in_43_13), .o(n_7274) );
in01f80 g571152 ( .a(x_in_17_15), .o(n_2549) );
in01f80 g571153 ( .a(x_in_18_1), .o(n_16354) );
in01f80 g571154 ( .a(x_in_53_8), .o(n_2654) );
in01f80 g571155 ( .a(x_in_63_7), .o(n_7903) );
in01f80 g571156 ( .a(x_in_63_2), .o(n_5351) );
in01f80 g571157 ( .a(x_in_3_8), .o(n_5524) );
in01f80 g571158 ( .a(x_in_17_4), .o(n_4021) );
in01f80 g571159 ( .a(x_in_7_6), .o(n_5968) );
in01f80 g571160 ( .a(x_in_5_1), .o(n_2539) );
in01f80 g571161 ( .a(x_in_19_15), .o(n_149) );
in01f80 g571162 ( .a(x_in_41_10), .o(n_7915) );
in01f80 g571163 ( .a(x_in_21_9), .o(n_3887) );
in01f80 g571164 ( .a(x_in_50_1), .o(n_16031) );
in01f80 g571165 ( .a(x_in_13_1), .o(n_2707) );
in01f80 g571166 ( .a(x_in_57_11), .o(n_5313) );
in01f80 g571167 ( .a(x_in_11_9), .o(n_5310) );
in01f80 g571168 ( .a(x_in_25_4), .o(n_2554) );
in01f80 g571169 ( .a(x_in_47_1), .o(n_2616) );
in01f80 g571170 ( .a(x_in_41_15), .o(n_1175) );
in01f80 g571171 ( .a(x_in_32_15), .o(n_1383) );
in01f80 g571172 ( .a(x_in_25_2), .o(n_2535) );
in01f80 g571173 ( .a(x_in_57_12), .o(n_5302) );
in01f80 g571174 ( .a(x_in_53_3), .o(n_5827) );
in01f80 g571175 ( .a(x_in_52_1), .o(n_16227) );
in01f80 g571176 ( .a(x_in_1_2), .o(n_1036) );
in01f80 g571177 ( .a(x_in_21_5), .o(n_5900) );
in01f80 g571178 ( .a(x_in_15_7), .o(n_7904) );
in01f80 g571179 ( .a(x_in_33_1), .o(n_2452) );
in01f80 g571180 ( .a(x_in_43_10), .o(n_6496) );
in01f80 g571181 ( .a(x_in_5_14), .o(n_3169) );
in01f80 g573176 ( .a(n_3918), .o(n_32729) );
in01f80 g573177 ( .a(n_6330), .o(n_32730) );
in01f80 g573178 ( .a(n_4332), .o(n_32731) );
no02f80 g573179 ( .a(n_9798), .b(n_9796), .o(n_32733) );
no02f80 g573180 ( .a(n_8015), .b(n_8014), .o(n_32734) );
oa12f80 g573181 ( .a(n_5396), .b(n_5357), .c(x_in_17_13), .o(n_32735) );
no02f80 g573182 ( .a(FE_OFN931_n_4898), .b(n_5283), .o(n_32736) );
no02f80 g573183 ( .a(n_2596), .b(x_in_31_15), .o(n_32737) );
no02f80 g573184 ( .a(n_3872), .b(x_in_15_15), .o(n_32738) );
no02f80 g573185 ( .a(n_3870), .b(x_in_47_15), .o(n_32739) );
no02f80 g573186 ( .a(n_2401), .b(x_in_23_15), .o(n_32740) );
no02f80 g573187 ( .a(n_2532), .b(x_in_55_15), .o(n_32741) );
no02f80 g573188 ( .a(n_3793), .b(n_3792), .o(n_32742) );
no02f80 g573189 ( .a(n_3504), .b(x_in_63_15), .o(n_32743) );
ms00f80 x_out_0_reg_0_ ( .ck(ispd_clk), .d(n_7222), .o(x_out_0_0) );
ms00f80 x_out_0_reg_10_ ( .ck(ispd_clk), .d(n_22107), .o(x_out_0_10) );
ms00f80 x_out_0_reg_11_ ( .ck(ispd_clk), .d(n_23370), .o(x_out_0_11) );
ms00f80 x_out_0_reg_12_ ( .ck(ispd_clk), .d(n_24666), .o(x_out_0_12) );
ms00f80 x_out_0_reg_13_ ( .ck(ispd_clk), .d(n_25934), .o(x_out_0_13) );
ms00f80 x_out_0_reg_14_ ( .ck(ispd_clk), .d(n_26847), .o(x_out_0_14) );
ms00f80 x_out_0_reg_15_ ( .ck(ispd_clk), .d(n_27748), .o(x_out_0_15) );
ms00f80 x_out_0_reg_1_ ( .ck(ispd_clk), .d(n_7998), .o(x_out_0_1) );
ms00f80 x_out_0_reg_2_ ( .ck(ispd_clk), .d(n_10124), .o(x_out_0_2) );
ms00f80 x_out_0_reg_3_ ( .ck(ispd_clk), .d(n_12240), .o(x_out_0_3) );
ms00f80 x_out_0_reg_4_ ( .ck(ispd_clk), .d(n_14426), .o(x_out_0_4) );
ms00f80 x_out_0_reg_5_ ( .ck(ispd_clk), .d(n_15978), .o(x_out_0_5) );
ms00f80 x_out_0_reg_6_ ( .ck(ispd_clk), .d(n_17114), .o(x_out_0_6) );
ms00f80 x_out_0_reg_7_ ( .ck(ispd_clk), .d(n_18322), .o(x_out_0_7) );
ms00f80 x_out_0_reg_8_ ( .ck(ispd_clk), .d(n_19557), .o(x_out_0_8) );
ms00f80 x_out_0_reg_9_ ( .ck(ispd_clk), .d(n_21007), .o(x_out_0_9) );
ms00f80 x_out_10_reg_0_ ( .ck(ispd_clk), .d(n_17243), .o(x_out_10_0) );
ms00f80 x_out_10_reg_10_ ( .ck(ispd_clk), .d(n_28397), .o(x_out_10_10) );
ms00f80 x_out_10_reg_11_ ( .ck(ispd_clk), .d(n_28770), .o(x_out_10_11) );
ms00f80 x_out_10_reg_12_ ( .ck(ispd_clk), .d(n_29106), .o(x_out_10_12) );
ms00f80 x_out_10_reg_13_ ( .ck(ispd_clk), .d(n_29454), .o(x_out_10_13) );
ms00f80 x_out_10_reg_14_ ( .ck(ispd_clk), .d(n_29622), .o(x_out_10_14) );
ms00f80 x_out_10_reg_15_ ( .ck(ispd_clk), .d(n_29669), .o(x_out_10_15) );
ms00f80 x_out_10_reg_18_ ( .ck(ispd_clk), .d(n_14625), .o(x_out_10_18) );
ms00f80 x_out_10_reg_19_ ( .ck(ispd_clk), .d(n_15201), .o(x_out_10_19) );
ms00f80 x_out_10_reg_1_ ( .ck(ispd_clk), .d(n_19746), .o(x_out_10_1) );
ms00f80 x_out_10_reg_20_ ( .ck(ispd_clk), .d(n_15933), .o(x_out_10_20) );
ms00f80 x_out_10_reg_21_ ( .ck(ispd_clk), .d(n_17076), .o(x_out_10_21) );
ms00f80 x_out_10_reg_22_ ( .ck(ispd_clk), .d(n_17773), .o(x_out_10_22) );
ms00f80 x_out_10_reg_23_ ( .ck(ispd_clk), .d(n_18983), .o(x_out_10_23) );
ms00f80 x_out_10_reg_24_ ( .ck(ispd_clk), .d(n_19650), .o(x_out_10_24) );
ms00f80 x_out_10_reg_25_ ( .ck(ispd_clk), .d(n_20796), .o(x_out_10_25) );
ms00f80 x_out_10_reg_26_ ( .ck(ispd_clk), .d(n_21543), .o(x_out_10_26) );
ms00f80 x_out_10_reg_27_ ( .ck(ispd_clk), .d(n_22854), .o(x_out_10_27) );
ms00f80 x_out_10_reg_28_ ( .ck(ispd_clk), .d(n_23551), .o(x_out_10_28) );
ms00f80 x_out_10_reg_29_ ( .ck(ispd_clk), .d(n_24497), .o(x_out_10_29) );
ms00f80 x_out_10_reg_2_ ( .ck(ispd_clk), .d(n_20893), .o(x_out_10_2) );
ms00f80 x_out_10_reg_30_ ( .ck(ispd_clk), .d(n_25255), .o(x_out_10_30) );
ms00f80 x_out_10_reg_31_ ( .ck(ispd_clk), .d(n_26460), .o(x_out_10_31) );
ms00f80 x_out_10_reg_32_ ( .ck(ispd_clk), .d(n_27790), .o(x_out_10_32) );
ms00f80 x_out_10_reg_33_ ( .ck(ispd_clk), .d(n_27732), .o(x_out_10_33) );
ms00f80 x_out_10_reg_3_ ( .ck(ispd_clk), .d(n_21269), .o(x_out_10_3) );
ms00f80 x_out_10_reg_4_ ( .ck(ispd_clk), .d(n_22313), .o(x_out_10_4) );
ms00f80 x_out_10_reg_5_ ( .ck(ispd_clk), .d(n_23614), .o(x_out_10_5) );
ms00f80 x_out_10_reg_6_ ( .ck(ispd_clk), .d(n_24923), .o(x_out_10_6) );
ms00f80 x_out_10_reg_7_ ( .ck(ispd_clk), .d(n_26141), .o(x_out_10_7) );
ms00f80 x_out_10_reg_8_ ( .ck(ispd_clk), .d(n_27028), .o(x_out_10_8) );
ms00f80 x_out_10_reg_9_ ( .ck(ispd_clk), .d(n_27866), .o(x_out_10_9) );
ms00f80 x_out_11_reg_0_ ( .ck(ispd_clk), .d(n_16802), .o(x_out_11_0) );
ms00f80 x_out_11_reg_10_ ( .ck(ispd_clk), .d(n_27934), .o(x_out_11_10) );
ms00f80 x_out_11_reg_11_ ( .ck(ispd_clk), .d(n_28366), .o(x_out_11_11) );
ms00f80 x_out_11_reg_12_ ( .ck(ispd_clk), .d(n_28748), .o(x_out_11_12) );
ms00f80 x_out_11_reg_13_ ( .ck(ispd_clk), .d(n_29101), .o(x_out_11_13) );
ms00f80 x_out_11_reg_14_ ( .ck(ispd_clk), .d(n_29415), .o(x_out_11_14) );
ms00f80 x_out_11_reg_15_ ( .ck(ispd_clk), .d(n_29580), .o(x_out_11_15) );
ms00f80 x_out_11_reg_18_ ( .ck(ispd_clk), .d(n_17226), .o(x_out_11_18) );
ms00f80 x_out_11_reg_19_ ( .ck(ispd_clk), .d(n_17398), .o(x_out_11_19) );
ms00f80 x_out_11_reg_1_ ( .ck(ispd_clk), .d(n_18284), .o(x_out_11_1) );
ms00f80 x_out_11_reg_20_ ( .ck(ispd_clk), .d(n_18016), .o(x_out_11_20) );
ms00f80 x_out_11_reg_21_ ( .ck(ispd_clk), .d(n_18645), .o(x_out_11_21) );
ms00f80 x_out_11_reg_22_ ( .ck(ispd_clk), .d(n_19995), .o(x_out_11_22) );
ms00f80 x_out_11_reg_23_ ( .ck(ispd_clk), .d(n_20441), .o(x_out_11_23) );
ms00f80 x_out_11_reg_24_ ( .ck(ispd_clk), .d(n_21905), .o(x_out_11_24) );
ms00f80 x_out_11_reg_25_ ( .ck(ispd_clk), .d(n_22553), .o(x_out_11_25) );
ms00f80 x_out_11_reg_26_ ( .ck(ispd_clk), .d(n_23812), .o(x_out_11_26) );
ms00f80 x_out_11_reg_27_ ( .ck(ispd_clk), .d(n_24179), .o(x_out_11_27) );
ms00f80 x_out_11_reg_28_ ( .ck(ispd_clk), .d(n_25523), .o(x_out_11_28) );
ms00f80 x_out_11_reg_29_ ( .ck(ispd_clk), .d(n_26170), .o(x_out_11_29) );
ms00f80 x_out_11_reg_2_ ( .ck(ispd_clk), .d(n_19837), .o(x_out_11_2) );
ms00f80 x_out_11_reg_30_ ( .ck(ispd_clk), .d(n_27154), .o(x_out_11_30) );
ms00f80 x_out_11_reg_31_ ( .ck(ispd_clk), .d(n_27458), .o(x_out_11_31) );
ms00f80 x_out_11_reg_32_ ( .ck(ispd_clk), .d(n_28261), .o(x_out_11_32) );
ms00f80 x_out_11_reg_33_ ( .ck(ispd_clk), .d(n_28759), .o(x_out_11_33) );
ms00f80 x_out_11_reg_3_ ( .ck(ispd_clk), .d(n_21266), .o(x_out_11_3) );
ms00f80 x_out_11_reg_4_ ( .ck(ispd_clk), .d(n_21770), .o(x_out_11_4) );
ms00f80 x_out_11_reg_5_ ( .ck(ispd_clk), .d(n_23051), .o(x_out_11_5) );
ms00f80 x_out_11_reg_6_ ( .ck(ispd_clk), .d(n_24298), .o(x_out_11_6) );
ms00f80 x_out_11_reg_7_ ( .ck(ispd_clk), .d(n_25667), .o(x_out_11_7) );
ms00f80 x_out_11_reg_8_ ( .ck(ispd_clk), .d(n_26234), .o(x_out_11_8) );
ms00f80 x_out_11_reg_9_ ( .ck(ispd_clk), .d(n_27153), .o(x_out_11_9) );
ms00f80 x_out_12_reg_0_ ( .ck(ispd_clk), .d(n_14362), .o(x_out_12_0) );
ms00f80 x_out_12_reg_10_ ( .ck(ispd_clk), .d(n_27350), .o(x_out_12_10) );
ms00f80 x_out_12_reg_11_ ( .ck(ispd_clk), .d(n_28086), .o(x_out_12_11) );
ms00f80 x_out_12_reg_12_ ( .ck(ispd_clk), .d(n_28481), .o(x_out_12_12) );
ms00f80 x_out_12_reg_13_ ( .ck(ispd_clk), .d(n_28822), .o(x_out_12_13) );
ms00f80 x_out_12_reg_14_ ( .ck(ispd_clk), .d(n_29208), .o(x_out_12_14) );
ms00f80 x_out_12_reg_15_ ( .ck(ispd_clk), .d(n_29495), .o(x_out_12_15) );
ms00f80 x_out_12_reg_18_ ( .ck(ispd_clk), .d(n_6046), .o(x_out_12_18) );
ms00f80 x_out_12_reg_19_ ( .ck(ispd_clk), .d(n_7437), .o(x_out_12_19) );
ms00f80 x_out_12_reg_1_ ( .ck(ispd_clk), .d(n_17921), .o(x_out_12_1) );
ms00f80 x_out_12_reg_20_ ( .ck(ispd_clk), .d(n_7997), .o(x_out_12_20) );
ms00f80 x_out_12_reg_21_ ( .ck(ispd_clk), .d(n_11677), .o(x_out_12_21) );
ms00f80 x_out_12_reg_22_ ( .ck(ispd_clk), .d(n_11675), .o(x_out_12_22) );
ms00f80 x_out_12_reg_23_ ( .ck(ispd_clk), .d(n_12855), .o(x_out_12_23) );
ms00f80 x_out_12_reg_24_ ( .ck(ispd_clk), .d(n_13762), .o(x_out_12_24) );
ms00f80 x_out_12_reg_25_ ( .ck(ispd_clk), .d(n_15637), .o(x_out_12_25) );
ms00f80 x_out_12_reg_26_ ( .ck(ispd_clk), .d(n_16350), .o(x_out_12_26) );
ms00f80 x_out_12_reg_27_ ( .ck(ispd_clk), .d(n_17493), .o(x_out_12_27) );
ms00f80 x_out_12_reg_28_ ( .ck(ispd_clk), .d(n_18098), .o(x_out_12_28) );
ms00f80 x_out_12_reg_29_ ( .ck(ispd_clk), .d(n_19389), .o(x_out_12_29) );
ms00f80 x_out_12_reg_2_ ( .ck(ispd_clk), .d(n_18283), .o(x_out_12_2) );
ms00f80 x_out_12_reg_30_ ( .ck(ispd_clk), .d(n_19724), .o(x_out_12_30) );
ms00f80 x_out_12_reg_31_ ( .ck(ispd_clk), .d(n_21191), .o(x_out_12_31) );
ms00f80 x_out_12_reg_32_ ( .ck(ispd_clk), .d(n_22882), .o(x_out_12_32) );
ms00f80 x_out_12_reg_33_ ( .ck(ispd_clk), .d(n_22928), .o(x_out_12_33) );
ms00f80 x_out_12_reg_3_ ( .ck(ispd_clk), .d(n_20883), .o(x_out_12_3) );
ms00f80 x_out_12_reg_4_ ( .ck(ispd_clk), .d(n_20963), .o(x_out_12_4) );
ms00f80 x_out_12_reg_5_ ( .ck(ispd_clk), .d(n_22058), .o(x_out_12_5) );
ms00f80 x_out_12_reg_6_ ( .ck(ispd_clk), .d(n_23300), .o(x_out_12_6) );
ms00f80 x_out_12_reg_7_ ( .ck(ispd_clk), .d(n_24604), .o(x_out_12_7) );
ms00f80 x_out_12_reg_8_ ( .ck(ispd_clk), .d(n_25663), .o(x_out_12_8) );
ms00f80 x_out_12_reg_9_ ( .ck(ispd_clk), .d(n_26229), .o(x_out_12_9) );
ms00f80 x_out_13_reg_0_ ( .ck(ispd_clk), .d(n_14666), .o(x_out_13_0) );
ms00f80 x_out_13_reg_10_ ( .ck(ispd_clk), .d(n_27461), .o(x_out_13_10) );
ms00f80 x_out_13_reg_11_ ( .ck(ispd_clk), .d(n_28126), .o(x_out_13_11) );
ms00f80 x_out_13_reg_12_ ( .ck(ispd_clk), .d(n_28528), .o(x_out_13_12) );
ms00f80 x_out_13_reg_13_ ( .ck(ispd_clk), .d(n_28945), .o(x_out_13_13) );
ms00f80 x_out_13_reg_14_ ( .ck(ispd_clk), .d(n_29304), .o(x_out_13_14) );
ms00f80 x_out_13_reg_15_ ( .ck(ispd_clk), .d(n_29556), .o(x_out_13_15) );
ms00f80 x_out_13_reg_18_ ( .ck(ispd_clk), .d(n_11772), .o(x_out_13_18) );
ms00f80 x_out_13_reg_19_ ( .ck(ispd_clk), .d(n_15719), .o(x_out_13_19) );
ms00f80 x_out_13_reg_1_ ( .ck(ispd_clk), .d(n_17918), .o(x_out_13_1) );
ms00f80 x_out_13_reg_20_ ( .ck(ispd_clk), .d(n_15932), .o(x_out_13_20) );
ms00f80 x_out_13_reg_21_ ( .ck(ispd_clk), .d(n_16608), .o(x_out_13_21) );
ms00f80 x_out_13_reg_22_ ( .ck(ispd_clk), .d(n_18145), .o(x_out_13_22) );
ms00f80 x_out_13_reg_23_ ( .ck(ispd_clk), .d(n_18847), .o(x_out_13_23) );
ms00f80 x_out_13_reg_24_ ( .ck(ispd_clk), .d(n_19830), .o(x_out_13_24) );
ms00f80 x_out_13_reg_25_ ( .ck(ispd_clk), .d(n_20661), .o(x_out_13_25) );
ms00f80 x_out_13_reg_26_ ( .ck(ispd_clk), .d(n_22018), .o(x_out_13_26) );
ms00f80 x_out_13_reg_27_ ( .ck(ispd_clk), .d(n_22374), .o(x_out_13_27) );
ms00f80 x_out_13_reg_28_ ( .ck(ispd_clk), .d(n_23653), .o(x_out_13_28) );
ms00f80 x_out_13_reg_29_ ( .ck(ispd_clk), .d(n_24021), .o(x_out_13_29) );
ms00f80 x_out_13_reg_2_ ( .ck(ispd_clk), .d(n_18281), .o(x_out_13_2) );
ms00f80 x_out_13_reg_30_ ( .ck(ispd_clk), .d(n_25023), .o(x_out_13_30) );
ms00f80 x_out_13_reg_31_ ( .ck(ispd_clk), .d(n_25726), .o(x_out_13_31) );
ms00f80 x_out_13_reg_32_ ( .ck(ispd_clk), .d(n_27169), .o(x_out_13_32) );
ms00f80 x_out_13_reg_33_ ( .ck(ispd_clk), .d(n_27167), .o(x_out_13_33) );
ms00f80 x_out_13_reg_3_ ( .ck(ispd_clk), .d(n_19513), .o(x_out_13_3) );
ms00f80 x_out_13_reg_4_ ( .ck(ispd_clk), .d(n_20908), .o(x_out_13_4) );
ms00f80 x_out_13_reg_5_ ( .ck(ispd_clk), .d(n_22285), .o(x_out_13_5) );
ms00f80 x_out_13_reg_6_ ( .ck(ispd_clk), .d(n_22959), .o(x_out_13_6) );
ms00f80 x_out_13_reg_7_ ( .ck(ispd_clk), .d(n_24206), .o(x_out_13_7) );
ms00f80 x_out_13_reg_8_ ( .ck(ispd_clk), .d(n_25547), .o(x_out_13_8) );
ms00f80 x_out_13_reg_9_ ( .ck(ispd_clk), .d(n_26680), .o(x_out_13_9) );
ms00f80 x_out_14_reg_0_ ( .ck(ispd_clk), .d(n_8642), .o(x_out_14_0) );
ms00f80 x_out_14_reg_10_ ( .ck(ispd_clk), .d(n_26451), .o(x_out_14_10) );
ms00f80 x_out_14_reg_11_ ( .ck(ispd_clk), .d(n_27264), .o(x_out_14_11) );
ms00f80 x_out_14_reg_12_ ( .ck(ispd_clk), .d(n_28012), .o(x_out_14_12) );
ms00f80 x_out_14_reg_13_ ( .ck(ispd_clk), .d(n_28425), .o(x_out_14_13) );
ms00f80 x_out_14_reg_14_ ( .ck(ispd_clk), .d(n_28868), .o(x_out_14_14) );
ms00f80 x_out_14_reg_15_ ( .ck(ispd_clk), .d(n_29207), .o(x_out_14_15) );
ms00f80 x_out_14_reg_18_ ( .ck(ispd_clk), .d(n_11494), .o(x_out_14_18) );
ms00f80 x_out_14_reg_19_ ( .ck(ispd_clk), .d(n_16367), .o(x_out_14_19) );
ms00f80 x_out_14_reg_1_ ( .ck(ispd_clk), .d(n_13355), .o(x_out_14_1) );
ms00f80 x_out_14_reg_20_ ( .ck(ispd_clk), .d(n_15182), .o(x_out_14_20) );
ms00f80 x_out_14_reg_21_ ( .ck(ispd_clk), .d(n_16220), .o(x_out_14_21) );
ms00f80 x_out_14_reg_22_ ( .ck(ispd_clk), .d(n_17367), .o(x_out_14_22) );
ms00f80 x_out_14_reg_23_ ( .ck(ispd_clk), .d(n_18009), .o(x_out_14_23) );
ms00f80 x_out_14_reg_24_ ( .ck(ispd_clk), .d(n_19279), .o(x_out_14_24) );
ms00f80 x_out_14_reg_25_ ( .ck(ispd_clk), .d(n_19990), .o(x_out_14_25) );
ms00f80 x_out_14_reg_26_ ( .ck(ispd_clk), .d(n_21078), .o(x_out_14_26) );
ms00f80 x_out_14_reg_27_ ( .ck(ispd_clk), .d(n_21898), .o(x_out_14_27) );
ms00f80 x_out_14_reg_28_ ( .ck(ispd_clk), .d(n_23131), .o(x_out_14_28) );
ms00f80 x_out_14_reg_29_ ( .ck(ispd_clk), .d(n_23806), .o(x_out_14_29) );
ms00f80 x_out_14_reg_2_ ( .ck(ispd_clk), .d(n_14128), .o(x_out_14_2) );
ms00f80 x_out_14_reg_30_ ( .ck(ispd_clk), .d(n_25093), .o(x_out_14_30) );
ms00f80 x_out_14_reg_31_ ( .ck(ispd_clk), .d(n_26310), .o(x_out_14_31) );
ms00f80 x_out_14_reg_32_ ( .ck(ispd_clk), .d(n_25141), .o(x_out_14_32) );
ms00f80 x_out_14_reg_33_ ( .ck(ispd_clk), .d(n_25140), .o(x_out_14_33) );
ms00f80 x_out_14_reg_3_ ( .ck(ispd_clk), .d(n_18793), .o(x_out_14_3) );
ms00f80 x_out_14_reg_4_ ( .ck(ispd_clk), .d(n_19151), .o(x_out_14_4) );
ms00f80 x_out_14_reg_5_ ( .ck(ispd_clk), .d(n_20222), .o(x_out_14_5) );
ms00f80 x_out_14_reg_6_ ( .ck(ispd_clk), .d(n_21639), .o(x_out_14_6) );
ms00f80 x_out_14_reg_7_ ( .ck(ispd_clk), .d(n_22643), .o(x_out_14_7) );
ms00f80 x_out_14_reg_8_ ( .ck(ispd_clk), .d(n_23938), .o(x_out_14_8) );
ms00f80 x_out_14_reg_9_ ( .ck(ispd_clk), .d(n_25283), .o(x_out_14_9) );
ms00f80 x_out_15_reg_0_ ( .ck(ispd_clk), .d(n_17521), .o(x_out_15_0) );
ms00f80 x_out_15_reg_10_ ( .ck(ispd_clk), .d(n_28294), .o(x_out_15_10) );
ms00f80 x_out_15_reg_11_ ( .ck(ispd_clk), .d(n_28693), .o(x_out_15_11) );
ms00f80 x_out_15_reg_12_ ( .ck(ispd_clk), .d(n_29047), .o(x_out_15_12) );
ms00f80 x_out_15_reg_13_ ( .ck(ispd_clk), .d(n_29347), .o(x_out_15_13) );
ms00f80 x_out_15_reg_14_ ( .ck(ispd_clk), .d(n_29533), .o(x_out_15_14) );
ms00f80 x_out_15_reg_15_ ( .ck(ispd_clk), .d(n_29652), .o(x_out_15_15) );
ms00f80 x_out_15_reg_18_ ( .ck(ispd_clk), .d(n_15756), .o(x_out_15_18) );
ms00f80 x_out_15_reg_19_ ( .ck(ispd_clk), .d(n_17228), .o(x_out_15_19) );
ms00f80 x_out_15_reg_1_ ( .ck(ispd_clk), .d(n_19441), .o(x_out_15_1) );
ms00f80 x_out_15_reg_20_ ( .ck(ispd_clk), .d(n_17082), .o(x_out_15_20) );
ms00f80 x_out_15_reg_21_ ( .ck(ispd_clk), .d(n_18285), .o(x_out_15_21) );
ms00f80 x_out_15_reg_22_ ( .ck(ispd_clk), .d(n_18990), .o(x_out_15_22) );
ms00f80 x_out_15_reg_23_ ( .ck(ispd_clk), .d(n_20320), .o(x_out_15_23) );
ms00f80 x_out_15_reg_24_ ( .ck(ispd_clk), .d(n_20803), .o(x_out_15_24) );
ms00f80 x_out_15_reg_25_ ( .ck(ispd_clk), .d(n_22159), .o(x_out_15_25) );
ms00f80 x_out_15_reg_26_ ( .ck(ispd_clk), .d(n_22852), .o(x_out_15_26) );
ms00f80 x_out_15_reg_27_ ( .ck(ispd_clk), .d(n_24090), .o(x_out_15_27) );
ms00f80 x_out_15_reg_28_ ( .ck(ispd_clk), .d(n_24495), .o(x_out_15_28) );
ms00f80 x_out_15_reg_29_ ( .ck(ispd_clk), .d(n_25799), .o(x_out_15_29) );
ms00f80 x_out_15_reg_2_ ( .ck(ispd_clk), .d(n_20187), .o(x_out_15_2) );
ms00f80 x_out_15_reg_30_ ( .ck(ispd_clk), .d(n_26452), .o(x_out_15_30) );
ms00f80 x_out_15_reg_31_ ( .ck(ispd_clk), .d(n_27372), .o(x_out_15_31) );
ms00f80 x_out_15_reg_32_ ( .ck(ispd_clk), .d(n_27694), .o(x_out_15_32) );
ms00f80 x_out_15_reg_33_ ( .ck(ispd_clk), .d(n_27693), .o(x_out_15_33) );
ms00f80 x_out_15_reg_3_ ( .ck(ispd_clk), .d(n_21267), .o(x_out_15_3) );
ms00f80 x_out_15_reg_4_ ( .ck(ispd_clk), .d(n_22067), .o(x_out_15_4) );
ms00f80 x_out_15_reg_5_ ( .ck(ispd_clk), .d(n_23319), .o(x_out_15_5) );
ms00f80 x_out_15_reg_6_ ( .ck(ispd_clk), .d(n_24617), .o(x_out_15_6) );
ms00f80 x_out_15_reg_7_ ( .ck(ispd_clk), .d(n_25897), .o(x_out_15_7) );
ms00f80 x_out_15_reg_8_ ( .ck(ispd_clk), .d(n_26808), .o(x_out_15_8) );
ms00f80 x_out_15_reg_9_ ( .ck(ispd_clk), .d(n_27710), .o(x_out_15_9) );
ms00f80 x_out_16_reg_0_ ( .ck(ispd_clk), .d(n_15555), .o(x_out_16_0) );
ms00f80 x_out_16_reg_10_ ( .ck(ispd_clk), .d(n_27708), .o(x_out_16_10) );
ms00f80 x_out_16_reg_11_ ( .ck(ispd_clk), .d(n_28314), .o(x_out_16_11) );
ms00f80 x_out_16_reg_12_ ( .ck(ispd_clk), .d(n_28686), .o(x_out_16_12) );
ms00f80 x_out_16_reg_13_ ( .ck(ispd_clk), .d(n_29037), .o(x_out_16_13) );
ms00f80 x_out_16_reg_14_ ( .ck(ispd_clk), .d(n_29340), .o(x_out_16_14) );
ms00f80 x_out_16_reg_15_ ( .ck(ispd_clk), .d(n_29619), .o(x_out_16_15) );
ms00f80 x_out_16_reg_18_ ( .ck(ispd_clk), .d(n_11490), .o(x_out_16_18) );
ms00f80 x_out_16_reg_19_ ( .ck(ispd_clk), .d(n_16079), .o(x_out_16_19) );
ms00f80 x_out_16_reg_1_ ( .ck(ispd_clk), .d(n_18150), .o(x_out_16_1) );
ms00f80 x_out_16_reg_20_ ( .ck(ispd_clk), .d(n_16036), .o(x_out_16_20) );
ms00f80 x_out_16_reg_21_ ( .ck(ispd_clk), .d(n_15941), .o(x_out_16_21) );
ms00f80 x_out_16_reg_22_ ( .ck(ispd_clk), .d(n_16925), .o(x_out_16_22) );
ms00f80 x_out_16_reg_23_ ( .ck(ispd_clk), .d(n_17702), .o(x_out_16_23) );
ms00f80 x_out_16_reg_24_ ( .ck(ispd_clk), .d(n_18852), .o(x_out_16_24) );
ms00f80 x_out_16_reg_25_ ( .ck(ispd_clk), .d(n_19560), .o(x_out_16_25) );
ms00f80 x_out_16_reg_26_ ( .ck(ispd_clk), .d(n_21010), .o(x_out_16_26) );
ms00f80 x_out_16_reg_27_ ( .ck(ispd_clk), .d(n_21454), .o(x_out_16_27) );
ms00f80 x_out_16_reg_28_ ( .ck(ispd_clk), .d(n_22753), .o(x_out_16_28) );
ms00f80 x_out_16_reg_29_ ( .ck(ispd_clk), .d(n_23454), .o(x_out_16_29) );
ms00f80 x_out_16_reg_2_ ( .ck(ispd_clk), .d(n_18529), .o(x_out_16_2) );
ms00f80 x_out_16_reg_30_ ( .ck(ispd_clk), .d(n_24713), .o(x_out_16_30) );
ms00f80 x_out_16_reg_31_ ( .ck(ispd_clk), .d(n_25745), .o(x_out_16_31) );
ms00f80 x_out_16_reg_32_ ( .ck(ispd_clk), .d(n_26955), .o(x_out_16_32) );
ms00f80 x_out_16_reg_33_ ( .ck(ispd_clk), .d(n_26954), .o(x_out_16_33) );
ms00f80 x_out_16_reg_3_ ( .ck(ispd_clk), .d(n_20184), .o(x_out_16_3) );
ms00f80 x_out_16_reg_4_ ( .ck(ispd_clk), .d(n_20970), .o(x_out_16_4) );
ms00f80 x_out_16_reg_5_ ( .ck(ispd_clk), .d(n_22069), .o(x_out_16_5) );
ms00f80 x_out_16_reg_6_ ( .ck(ispd_clk), .d(n_23308), .o(x_out_16_6) );
ms00f80 x_out_16_reg_7_ ( .ck(ispd_clk), .d(n_24612), .o(x_out_16_7) );
ms00f80 x_out_16_reg_8_ ( .ck(ispd_clk), .d(n_25892), .o(x_out_16_8) );
ms00f80 x_out_16_reg_9_ ( .ck(ispd_clk), .d(n_26796), .o(x_out_16_9) );
ms00f80 x_out_17_reg_0_ ( .ck(ispd_clk), .d(n_16375), .o(x_out_17_0) );
ms00f80 x_out_17_reg_10_ ( .ck(ispd_clk), .d(n_27989), .o(x_out_17_10) );
ms00f80 x_out_17_reg_11_ ( .ck(ispd_clk), .d(n_28513), .o(x_out_17_11) );
ms00f80 x_out_17_reg_12_ ( .ck(ispd_clk), .d(n_28848), .o(x_out_17_12) );
ms00f80 x_out_17_reg_13_ ( .ck(ispd_clk), .d(n_29179), .o(x_out_17_13) );
ms00f80 x_out_17_reg_14_ ( .ck(ispd_clk), .d(n_29522), .o(x_out_17_14) );
ms00f80 x_out_17_reg_15_ ( .ck(ispd_clk), .d(n_29654), .o(x_out_17_15) );
ms00f80 x_out_17_reg_18_ ( .ck(ispd_clk), .d(n_16646), .o(x_out_17_18) );
ms00f80 x_out_17_reg_19_ ( .ck(ispd_clk), .d(n_17255), .o(x_out_17_19) );
ms00f80 x_out_17_reg_1_ ( .ck(ispd_clk), .d(n_18148), .o(x_out_17_1) );
ms00f80 x_out_17_reg_20_ ( .ck(ispd_clk), .d(n_17846), .o(x_out_17_20) );
ms00f80 x_out_17_reg_21_ ( .ck(ispd_clk), .d(n_18523), .o(x_out_17_21) );
ms00f80 x_out_17_reg_22_ ( .ck(ispd_clk), .d(n_19836), .o(x_out_17_22) );
ms00f80 x_out_17_reg_23_ ( .ck(ispd_clk), .d(n_20663), .o(x_out_17_23) );
ms00f80 x_out_17_reg_24_ ( .ck(ispd_clk), .d(n_21769), .o(x_out_17_24) );
ms00f80 x_out_17_reg_25_ ( .ck(ispd_clk), .d(n_22429), .o(x_out_17_25) );
ms00f80 x_out_17_reg_26_ ( .ck(ispd_clk), .d(n_23693), .o(x_out_17_26) );
ms00f80 x_out_17_reg_27_ ( .ck(ispd_clk), .d(n_24362), .o(x_out_17_27) );
ms00f80 x_out_17_reg_28_ ( .ck(ispd_clk), .d(n_25403), .o(x_out_17_28) );
ms00f80 x_out_17_reg_29_ ( .ck(ispd_clk), .d(n_26012), .o(x_out_17_29) );
ms00f80 x_out_17_reg_2_ ( .ck(ispd_clk), .d(n_18799), .o(x_out_17_2) );
ms00f80 x_out_17_reg_30_ ( .ck(ispd_clk), .d(n_27433), .o(x_out_17_30) );
ms00f80 x_out_17_reg_31_ ( .ck(ispd_clk), .d(n_27756), .o(x_out_17_31) );
ms00f80 x_out_17_reg_32_ ( .ck(ispd_clk), .d(n_27755), .o(x_out_17_32) );
ms00f80 x_out_17_reg_33_ ( .ck(ispd_clk), .d(n_27753), .o(x_out_17_33) );
ms00f80 x_out_17_reg_3_ ( .ck(ispd_clk), .d(n_20183), .o(x_out_17_3) );
ms00f80 x_out_17_reg_4_ ( .ck(ispd_clk), .d(n_21603), .o(x_out_17_4) );
ms00f80 x_out_17_reg_5_ ( .ck(ispd_clk), .d(n_22611), .o(x_out_17_5) );
ms00f80 x_out_17_reg_6_ ( .ck(ispd_clk), .d(n_23921), .o(x_out_17_6) );
ms00f80 x_out_17_reg_7_ ( .ck(ispd_clk), .d(n_25256), .o(x_out_17_7) );
ms00f80 x_out_17_reg_8_ ( .ck(ispd_clk), .d(n_26397), .o(x_out_17_8) );
ms00f80 x_out_17_reg_9_ ( .ck(ispd_clk), .d(n_27248), .o(x_out_17_9) );
ms00f80 x_out_18_reg_0_ ( .ck(ispd_clk), .d(n_15214), .o(x_out_18_0) );
ms00f80 x_out_18_reg_10_ ( .ck(ispd_clk), .d(n_27548), .o(x_out_18_10) );
ms00f80 x_out_18_reg_11_ ( .ck(ispd_clk), .d(n_28208), .o(x_out_18_11) );
ms00f80 x_out_18_reg_12_ ( .ck(ispd_clk), .d(n_28601), .o(x_out_18_12) );
ms00f80 x_out_18_reg_13_ ( .ck(ispd_clk), .d(n_28911), .o(x_out_18_13) );
ms00f80 x_out_18_reg_14_ ( .ck(ispd_clk), .d(n_29336), .o(x_out_18_14) );
ms00f80 x_out_18_reg_15_ ( .ck(ispd_clk), .d(n_29559), .o(x_out_18_15) );
ms00f80 x_out_18_reg_18_ ( .ck(ispd_clk), .d(n_13852), .o(x_out_18_18) );
ms00f80 x_out_18_reg_19_ ( .ck(ispd_clk), .d(n_16369), .o(x_out_18_19) );
ms00f80 x_out_18_reg_1_ ( .ck(ispd_clk), .d(n_18147), .o(x_out_18_1) );
ms00f80 x_out_18_reg_20_ ( .ck(ispd_clk), .d(n_16226), .o(x_out_18_20) );
ms00f80 x_out_18_reg_21_ ( .ck(ispd_clk), .d(n_17375), .o(x_out_18_21) );
ms00f80 x_out_18_reg_22_ ( .ck(ispd_clk), .d(n_18014), .o(x_out_18_22) );
ms00f80 x_out_18_reg_23_ ( .ck(ispd_clk), .d(n_19283), .o(x_out_18_23) );
ms00f80 x_out_18_reg_24_ ( .ck(ispd_clk), .d(n_19994), .o(x_out_18_24) );
ms00f80 x_out_18_reg_25_ ( .ck(ispd_clk), .d(n_21082), .o(x_out_18_25) );
ms00f80 x_out_18_reg_26_ ( .ck(ispd_clk), .d(n_21904), .o(x_out_18_26) );
ms00f80 x_out_18_reg_27_ ( .ck(ispd_clk), .d(n_23135), .o(x_out_18_27) );
ms00f80 x_out_18_reg_28_ ( .ck(ispd_clk), .d(n_23811), .o(x_out_18_28) );
ms00f80 x_out_18_reg_29_ ( .ck(ispd_clk), .d(n_24821), .o(x_out_18_29) );
ms00f80 x_out_18_reg_2_ ( .ck(ispd_clk), .d(n_18797), .o(x_out_18_2) );
ms00f80 x_out_18_reg_30_ ( .ck(ispd_clk), .d(n_26022), .o(x_out_18_30) );
ms00f80 x_out_18_reg_31_ ( .ck(ispd_clk), .d(n_27052), .o(x_out_18_31) );
ms00f80 x_out_18_reg_32_ ( .ck(ispd_clk), .d(n_27054), .o(x_out_18_32) );
ms00f80 x_out_18_reg_33_ ( .ck(ispd_clk), .d(n_27050), .o(x_out_18_33) );
ms00f80 x_out_18_reg_3_ ( .ck(ispd_clk), .d(n_19834), .o(x_out_18_3) );
ms00f80 x_out_18_reg_4_ ( .ck(ispd_clk), .d(n_20662), .o(x_out_18_4) );
ms00f80 x_out_18_reg_5_ ( .ck(ispd_clk), .d(n_21766), .o(x_out_18_5) );
ms00f80 x_out_18_reg_6_ ( .ck(ispd_clk), .d(n_23049), .o(x_out_18_6) );
ms00f80 x_out_18_reg_7_ ( .ck(ispd_clk), .d(n_24296), .o(x_out_18_7) );
ms00f80 x_out_18_reg_8_ ( .ck(ispd_clk), .d(n_25664), .o(x_out_18_8) );
ms00f80 x_out_18_reg_9_ ( .ck(ispd_clk), .d(n_26522), .o(x_out_18_9) );
ms00f80 x_out_19_reg_0_ ( .ck(ispd_clk), .d(n_15818), .o(x_out_19_0) );
ms00f80 x_out_19_reg_10_ ( .ck(ispd_clk), .d(n_27695), .o(x_out_19_10) );
ms00f80 x_out_19_reg_11_ ( .ck(ispd_clk), .d(n_28302), .o(x_out_19_11) );
ms00f80 x_out_19_reg_12_ ( .ck(ispd_clk), .d(n_28677), .o(x_out_19_12) );
ms00f80 x_out_19_reg_13_ ( .ck(ispd_clk), .d(n_29029), .o(x_out_19_13) );
ms00f80 x_out_19_reg_14_ ( .ck(ispd_clk), .d(n_29403), .o(x_out_19_14) );
ms00f80 x_out_19_reg_15_ ( .ck(ispd_clk), .d(n_29603), .o(x_out_19_15) );
ms00f80 x_out_19_reg_18_ ( .ck(ispd_clk), .d(n_17223), .o(x_out_19_18) );
ms00f80 x_out_19_reg_19_ ( .ck(ispd_clk), .d(n_17396), .o(x_out_19_19) );
ms00f80 x_out_19_reg_1_ ( .ck(ispd_clk), .d(n_18146), .o(x_out_19_1) );
ms00f80 x_out_19_reg_20_ ( .ck(ispd_clk), .d(n_18012), .o(x_out_19_20) );
ms00f80 x_out_19_reg_21_ ( .ck(ispd_clk), .d(n_19280), .o(x_out_19_21) );
ms00f80 x_out_19_reg_22_ ( .ck(ispd_clk), .d(n_19992), .o(x_out_19_22) );
ms00f80 x_out_19_reg_23_ ( .ck(ispd_clk), .d(n_21079), .o(x_out_19_23) );
ms00f80 x_out_19_reg_24_ ( .ck(ispd_clk), .d(n_21901), .o(x_out_19_24) );
ms00f80 x_out_19_reg_25_ ( .ck(ispd_clk), .d(n_23132), .o(x_out_19_25) );
ms00f80 x_out_19_reg_26_ ( .ck(ispd_clk), .d(n_23808), .o(x_out_19_26) );
ms00f80 x_out_19_reg_27_ ( .ck(ispd_clk), .d(n_24817), .o(x_out_19_27) );
ms00f80 x_out_19_reg_28_ ( .ck(ispd_clk), .d(n_25797), .o(x_out_19_28) );
ms00f80 x_out_19_reg_29_ ( .ck(ispd_clk), .d(n_27237), .o(x_out_19_29) );
ms00f80 x_out_19_reg_2_ ( .ck(ispd_clk), .d(n_18520), .o(x_out_19_2) );
ms00f80 x_out_19_reg_30_ ( .ck(ispd_clk), .d(n_27907), .o(x_out_19_30) );
ms00f80 x_out_19_reg_31_ ( .ck(ispd_clk), .d(n_27905), .o(x_out_19_31) );
ms00f80 x_out_19_reg_32_ ( .ck(ispd_clk), .d(n_27903), .o(x_out_19_32) );
ms00f80 x_out_19_reg_33_ ( .ck(ispd_clk), .d(n_27901), .o(x_out_19_33) );
ms00f80 x_out_19_reg_3_ ( .ck(ispd_clk), .d(n_19514), .o(x_out_19_3) );
ms00f80 x_out_19_reg_4_ ( .ck(ispd_clk), .d(n_20962), .o(x_out_19_4) );
ms00f80 x_out_19_reg_5_ ( .ck(ispd_clk), .d(n_22057), .o(x_out_19_5) );
ms00f80 x_out_19_reg_6_ ( .ck(ispd_clk), .d(n_23298), .o(x_out_19_6) );
ms00f80 x_out_19_reg_7_ ( .ck(ispd_clk), .d(n_24603), .o(x_out_19_7) );
ms00f80 x_out_19_reg_8_ ( .ck(ispd_clk), .d(n_25886), .o(x_out_19_8) );
ms00f80 x_out_19_reg_9_ ( .ck(ispd_clk), .d(n_26774), .o(x_out_19_9) );
ms00f80 x_out_1_reg_0_ ( .ck(ispd_clk), .d(n_16790), .o(x_out_1_0) );
ms00f80 x_out_1_reg_10_ ( .ck(ispd_clk), .d(n_27930), .o(x_out_1_10) );
ms00f80 x_out_1_reg_11_ ( .ck(ispd_clk), .d(n_28363), .o(x_out_1_11) );
ms00f80 x_out_1_reg_12_ ( .ck(ispd_clk), .d(n_28740), .o(x_out_1_12) );
ms00f80 x_out_1_reg_13_ ( .ck(ispd_clk), .d(n_29171), .o(x_out_1_13) );
ms00f80 x_out_1_reg_14_ ( .ck(ispd_clk), .d(n_29350), .o(x_out_1_14) );
ms00f80 x_out_1_reg_15_ ( .ck(ispd_clk), .d(n_29583), .o(x_out_1_15) );
ms00f80 x_out_1_reg_18_ ( .ck(ispd_clk), .d(n_14207), .o(x_out_1_18) );
ms00f80 x_out_1_reg_19_ ( .ck(ispd_clk), .d(n_16077), .o(x_out_1_19) );
ms00f80 x_out_1_reg_1_ ( .ck(ispd_clk), .d(n_18282), .o(x_out_1_1) );
ms00f80 x_out_1_reg_20_ ( .ck(ispd_clk), .d(n_16223), .o(x_out_1_20) );
ms00f80 x_out_1_reg_21_ ( .ck(ispd_clk), .d(n_16609), .o(x_out_1_21) );
ms00f80 x_out_1_reg_22_ ( .ck(ispd_clk), .d(n_17775), .o(x_out_1_22) );
ms00f80 x_out_1_reg_23_ ( .ck(ispd_clk), .d(n_18368), .o(x_out_1_23) );
ms00f80 x_out_1_reg_24_ ( .ck(ispd_clk), .d(n_19652), .o(x_out_1_24) );
ms00f80 x_out_1_reg_25_ ( .ck(ispd_clk), .d(n_20085), .o(x_out_1_25) );
ms00f80 x_out_1_reg_26_ ( .ck(ispd_clk), .d(n_21539), .o(x_out_1_26) );
ms00f80 x_out_1_reg_27_ ( .ck(ispd_clk), .d(n_22250), .o(x_out_1_27) );
ms00f80 x_out_1_reg_28_ ( .ck(ispd_clk), .d(n_23546), .o(x_out_1_28) );
ms00f80 x_out_1_reg_29_ ( .ck(ispd_clk), .d(n_23884), .o(x_out_1_29) );
ms00f80 x_out_1_reg_2_ ( .ck(ispd_clk), .d(n_19831), .o(x_out_1_2) );
ms00f80 x_out_1_reg_30_ ( .ck(ispd_clk), .d(n_25537), .o(x_out_1_30) );
ms00f80 x_out_1_reg_31_ ( .ck(ispd_clk), .d(n_26258), .o(x_out_1_31) );
ms00f80 x_out_1_reg_32_ ( .ck(ispd_clk), .d(n_26257), .o(x_out_1_32) );
ms00f80 x_out_1_reg_33_ ( .ck(ispd_clk), .d(n_26255), .o(x_out_1_33) );
ms00f80 x_out_1_reg_3_ ( .ck(ispd_clk), .d(n_21600), .o(x_out_1_3) );
ms00f80 x_out_1_reg_4_ ( .ck(ispd_clk), .d(n_21765), .o(x_out_1_4) );
ms00f80 x_out_1_reg_5_ ( .ck(ispd_clk), .d(n_23047), .o(x_out_1_5) );
ms00f80 x_out_1_reg_6_ ( .ck(ispd_clk), .d(n_24292), .o(x_out_1_6) );
ms00f80 x_out_1_reg_7_ ( .ck(ispd_clk), .d(n_25658), .o(x_out_1_7) );
ms00f80 x_out_1_reg_8_ ( .ck(ispd_clk), .d(n_26223), .o(x_out_1_8) );
ms00f80 x_out_1_reg_9_ ( .ck(ispd_clk), .d(n_27149), .o(x_out_1_9) );
ms00f80 x_out_20_reg_0_ ( .ck(ispd_clk), .d(n_15791), .o(x_out_20_0) );
ms00f80 x_out_20_reg_10_ ( .ck(ispd_clk), .d(n_27691), .o(x_out_20_10) );
ms00f80 x_out_20_reg_11_ ( .ck(ispd_clk), .d(n_28299), .o(x_out_20_11) );
ms00f80 x_out_20_reg_12_ ( .ck(ispd_clk), .d(n_28674), .o(x_out_20_12) );
ms00f80 x_out_20_reg_13_ ( .ck(ispd_clk), .d(n_29026), .o(x_out_20_13) );
ms00f80 x_out_20_reg_14_ ( .ck(ispd_clk), .d(n_29400), .o(x_out_20_14) );
ms00f80 x_out_20_reg_15_ ( .ck(ispd_clk), .d(n_29589), .o(x_out_20_15) );
ms00f80 x_out_20_reg_1_ ( .ck(ispd_clk), .d(n_17916), .o(x_out_20_1) );
ms00f80 x_out_20_reg_2_ ( .ck(ispd_clk), .d(n_18795), .o(x_out_20_2) );
ms00f80 x_out_20_reg_3_ ( .ck(ispd_clk), .d(n_19829), .o(x_out_20_3) );
ms00f80 x_out_20_reg_4_ ( .ck(ispd_clk), .d(n_20960), .o(x_out_20_4) );
ms00f80 x_out_20_reg_5_ ( .ck(ispd_clk), .d(n_22054), .o(x_out_20_5) );
ms00f80 x_out_20_reg_6_ ( .ck(ispd_clk), .d(n_23296), .o(x_out_20_6) );
ms00f80 x_out_20_reg_7_ ( .ck(ispd_clk), .d(n_24600), .o(x_out_20_7) );
ms00f80 x_out_20_reg_8_ ( .ck(ispd_clk), .d(n_25883), .o(x_out_20_8) );
ms00f80 x_out_20_reg_9_ ( .ck(ispd_clk), .d(n_26767), .o(x_out_20_9) );
ms00f80 x_out_21_reg_0_ ( .ck(ispd_clk), .d(n_15854), .o(x_out_21_0) );
ms00f80 x_out_21_reg_10_ ( .ck(ispd_clk), .d(n_27686), .o(x_out_21_10) );
ms00f80 x_out_21_reg_11_ ( .ck(ispd_clk), .d(n_28297), .o(x_out_21_11) );
ms00f80 x_out_21_reg_12_ ( .ck(ispd_clk), .d(n_28670), .o(x_out_21_12) );
ms00f80 x_out_21_reg_13_ ( .ck(ispd_clk), .d(n_29023), .o(x_out_21_13) );
ms00f80 x_out_21_reg_14_ ( .ck(ispd_clk), .d(n_29398), .o(x_out_21_14) );
ms00f80 x_out_21_reg_15_ ( .ck(ispd_clk), .d(n_29588), .o(x_out_21_15) );
ms00f80 x_out_21_reg_18_ ( .ck(ispd_clk), .d(n_8060), .o(x_out_21_18) );
ms00f80 x_out_21_reg_19_ ( .ck(ispd_clk), .d(n_6491), .o(x_out_21_19) );
ms00f80 x_out_21_reg_1_ ( .ck(ispd_clk), .d(n_17913), .o(x_out_21_1) );
ms00f80 x_out_21_reg_20_ ( .ck(ispd_clk), .d(n_7307), .o(x_out_21_20) );
ms00f80 x_out_21_reg_21_ ( .ck(ispd_clk), .d(n_7303), .o(x_out_21_21) );
ms00f80 x_out_21_reg_22_ ( .ck(ispd_clk), .d(n_7253), .o(x_out_21_22) );
ms00f80 x_out_21_reg_23_ ( .ck(ispd_clk), .d(n_7269), .o(x_out_21_23) );
ms00f80 x_out_21_reg_24_ ( .ck(ispd_clk), .d(n_6497), .o(x_out_21_24) );
ms00f80 x_out_21_reg_25_ ( .ck(ispd_clk), .d(n_7266), .o(x_out_21_25) );
ms00f80 x_out_21_reg_26_ ( .ck(ispd_clk), .d(n_7264), .o(x_out_21_26) );
ms00f80 x_out_21_reg_27_ ( .ck(ispd_clk), .d(n_7275), .o(x_out_21_27) );
ms00f80 x_out_21_reg_28_ ( .ck(ispd_clk), .d(n_7312), .o(x_out_21_28) );
ms00f80 x_out_21_reg_29_ ( .ck(ispd_clk), .d(n_6428), .o(x_out_21_29) );
ms00f80 x_out_21_reg_2_ ( .ck(ispd_clk), .d(n_18794), .o(x_out_21_2) );
ms00f80 x_out_21_reg_30_ ( .ck(ispd_clk), .d(n_5733), .o(x_out_21_30) );
ms00f80 x_out_21_reg_31_ ( .ck(ispd_clk), .d(n_7243), .o(x_out_21_31) );
ms00f80 x_out_21_reg_32_ ( .ck(ispd_clk), .d(n_8189), .o(x_out_21_32) );
ms00f80 x_out_21_reg_33_ ( .ck(ispd_clk), .d(n_7369), .o(x_out_21_33) );
ms00f80 x_out_21_reg_3_ ( .ck(ispd_clk), .d(n_19827), .o(x_out_21_3) );
ms00f80 x_out_21_reg_4_ ( .ck(ispd_clk), .d(n_20959), .o(x_out_21_4) );
ms00f80 x_out_21_reg_5_ ( .ck(ispd_clk), .d(n_22052), .o(x_out_21_5) );
ms00f80 x_out_21_reg_6_ ( .ck(ispd_clk), .d(n_23294), .o(x_out_21_6) );
ms00f80 x_out_21_reg_7_ ( .ck(ispd_clk), .d(n_24596), .o(x_out_21_7) );
ms00f80 x_out_21_reg_8_ ( .ck(ispd_clk), .d(n_25880), .o(x_out_21_8) );
ms00f80 x_out_21_reg_9_ ( .ck(ispd_clk), .d(n_26765), .o(x_out_21_9) );
ms00f80 x_out_22_reg_0_ ( .ck(ispd_clk), .d(n_15774), .o(x_out_22_0) );
ms00f80 x_out_22_reg_10_ ( .ck(ispd_clk), .d(n_27684), .o(x_out_22_10) );
ms00f80 x_out_22_reg_11_ ( .ck(ispd_clk), .d(n_28295), .o(x_out_22_11) );
ms00f80 x_out_22_reg_12_ ( .ck(ispd_clk), .d(n_28669), .o(x_out_22_12) );
ms00f80 x_out_22_reg_13_ ( .ck(ispd_clk), .d(n_29021), .o(x_out_22_13) );
ms00f80 x_out_22_reg_14_ ( .ck(ispd_clk), .d(n_29396), .o(x_out_22_14) );
ms00f80 x_out_22_reg_15_ ( .ck(ispd_clk), .d(n_29587), .o(x_out_22_15) );
ms00f80 x_out_22_reg_18_ ( .ck(ispd_clk), .d(n_7251), .o(x_out_22_18) );
ms00f80 x_out_22_reg_19_ ( .ck(ispd_clk), .d(n_7223), .o(x_out_22_19) );
ms00f80 x_out_22_reg_1_ ( .ck(ispd_clk), .d(n_17914), .o(x_out_22_1) );
ms00f80 x_out_22_reg_20_ ( .ck(ispd_clk), .d(n_7277), .o(x_out_22_20) );
ms00f80 x_out_22_reg_21_ ( .ck(ispd_clk), .d(n_7328), .o(x_out_22_21) );
ms00f80 x_out_22_reg_22_ ( .ck(ispd_clk), .d(n_6485), .o(x_out_22_22) );
ms00f80 x_out_22_reg_23_ ( .ck(ispd_clk), .d(n_7288), .o(x_out_22_23) );
ms00f80 x_out_22_reg_24_ ( .ck(ispd_clk), .d(n_7290), .o(x_out_22_24) );
ms00f80 x_out_22_reg_25_ ( .ck(ispd_clk), .d(n_7418), .o(x_out_22_25) );
ms00f80 x_out_22_reg_26_ ( .ck(ispd_clk), .d(n_7342), .o(x_out_22_26) );
ms00f80 x_out_22_reg_27_ ( .ck(ispd_clk), .d(n_7403), .o(x_out_22_27) );
ms00f80 x_out_22_reg_28_ ( .ck(ispd_clk), .d(n_7230), .o(x_out_22_28) );
ms00f80 x_out_22_reg_29_ ( .ck(ispd_clk), .d(n_7367), .o(x_out_22_29) );
ms00f80 x_out_22_reg_2_ ( .ck(ispd_clk), .d(n_18792), .o(x_out_22_2) );
ms00f80 x_out_22_reg_30_ ( .ck(ispd_clk), .d(n_6431), .o(x_out_22_30) );
ms00f80 x_out_22_reg_31_ ( .ck(ispd_clk), .d(n_7260), .o(x_out_22_31) );
ms00f80 x_out_22_reg_32_ ( .ck(ispd_clk), .d(n_8018), .o(x_out_22_32) );
ms00f80 x_out_22_reg_33_ ( .ck(ispd_clk), .d(n_7350), .o(x_out_22_33) );
ms00f80 x_out_22_reg_3_ ( .ck(ispd_clk), .d(n_20178), .o(x_out_22_3) );
ms00f80 x_out_22_reg_4_ ( .ck(ispd_clk), .d(n_20957), .o(x_out_22_4) );
ms00f80 x_out_22_reg_5_ ( .ck(ispd_clk), .d(n_22051), .o(x_out_22_5) );
ms00f80 x_out_22_reg_6_ ( .ck(ispd_clk), .d(n_23290), .o(x_out_22_6) );
ms00f80 x_out_22_reg_7_ ( .ck(ispd_clk), .d(n_24595), .o(x_out_22_7) );
ms00f80 x_out_22_reg_8_ ( .ck(ispd_clk), .d(n_25879), .o(x_out_22_8) );
ms00f80 x_out_22_reg_9_ ( .ck(ispd_clk), .d(n_27011), .o(x_out_22_9) );
ms00f80 x_out_23_reg_0_ ( .ck(ispd_clk), .d(n_16083), .o(x_out_23_0) );
ms00f80 x_out_23_reg_10_ ( .ck(ispd_clk), .d(n_27546), .o(x_out_23_10) );
ms00f80 x_out_23_reg_11_ ( .ck(ispd_clk), .d(n_28206), .o(x_out_23_11) );
ms00f80 x_out_23_reg_12_ ( .ck(ispd_clk), .d(n_28595), .o(x_out_23_12) );
ms00f80 x_out_23_reg_13_ ( .ck(ispd_clk), .d(n_28931), .o(x_out_23_13) );
ms00f80 x_out_23_reg_14_ ( .ck(ispd_clk), .d(n_29270), .o(x_out_23_14) );
ms00f80 x_out_23_reg_15_ ( .ck(ispd_clk), .d(n_29540), .o(x_out_23_15) );
ms00f80 x_out_23_reg_18_ ( .ck(ispd_clk), .d(n_13100), .o(x_out_23_18) );
ms00f80 x_out_23_reg_19_ ( .ck(ispd_clk), .d(n_13849), .o(x_out_23_19) );
ms00f80 x_out_23_reg_1_ ( .ck(ispd_clk), .d(n_17929), .o(x_out_23_1) );
ms00f80 x_out_23_reg_20_ ( .ck(ispd_clk), .d(n_14971), .o(x_out_23_20) );
ms00f80 x_out_23_reg_21_ ( .ck(ispd_clk), .d(n_16294), .o(x_out_23_21) );
ms00f80 x_out_23_reg_22_ ( .ck(ispd_clk), .d(n_17423), .o(x_out_23_22) );
ms00f80 x_out_23_reg_23_ ( .ck(ispd_clk), .d(n_18042), .o(x_out_23_23) );
ms00f80 x_out_23_reg_24_ ( .ck(ispd_clk), .d(n_19317), .o(x_out_23_24) );
ms00f80 x_out_23_reg_25_ ( .ck(ispd_clk), .d(n_20028), .o(x_out_23_25) );
ms00f80 x_out_23_reg_26_ ( .ck(ispd_clk), .d(n_21114), .o(x_out_23_26) );
ms00f80 x_out_23_reg_27_ ( .ck(ispd_clk), .d(n_21930), .o(x_out_23_27) );
ms00f80 x_out_23_reg_28_ ( .ck(ispd_clk), .d(n_23164), .o(x_out_23_28) );
ms00f80 x_out_23_reg_29_ ( .ck(ispd_clk), .d(n_23841), .o(x_out_23_29) );
ms00f80 x_out_23_reg_2_ ( .ck(ispd_clk), .d(n_18802), .o(x_out_23_2) );
ms00f80 x_out_23_reg_30_ ( .ck(ispd_clk), .d(n_25144), .o(x_out_23_30) );
ms00f80 x_out_23_reg_31_ ( .ck(ispd_clk), .d(n_7357), .o(x_out_23_31) );
ms00f80 x_out_23_reg_32_ ( .ck(ispd_clk), .d(n_7240), .o(x_out_23_32) );
ms00f80 x_out_23_reg_33_ ( .ck(ispd_clk), .d(n_6480), .o(x_out_23_33) );
ms00f80 x_out_23_reg_3_ ( .ck(ispd_clk), .d(n_19840), .o(x_out_23_3) );
ms00f80 x_out_23_reg_4_ ( .ck(ispd_clk), .d(n_20665), .o(x_out_23_4) );
ms00f80 x_out_23_reg_5_ ( .ck(ispd_clk), .d(n_21774), .o(x_out_23_5) );
ms00f80 x_out_23_reg_6_ ( .ck(ispd_clk), .d(n_23056), .o(x_out_23_6) );
ms00f80 x_out_23_reg_7_ ( .ck(ispd_clk), .d(n_24310), .o(x_out_23_7) );
ms00f80 x_out_23_reg_8_ ( .ck(ispd_clk), .d(n_25684), .o(x_out_23_8) );
ms00f80 x_out_23_reg_9_ ( .ck(ispd_clk), .d(n_26539), .o(x_out_23_9) );
ms00f80 x_out_24_reg_0_ ( .ck(ispd_clk), .d(n_17001), .o(x_out_24_0) );
ms00f80 x_out_24_reg_10_ ( .ck(ispd_clk), .d(n_28088), .o(x_out_24_10) );
ms00f80 x_out_24_reg_11_ ( .ck(ispd_clk), .d(n_28485), .o(x_out_24_11) );
ms00f80 x_out_24_reg_12_ ( .ck(ispd_clk), .d(n_28841), .o(x_out_24_12) );
ms00f80 x_out_24_reg_13_ ( .ck(ispd_clk), .d(n_29178), .o(x_out_24_13) );
ms00f80 x_out_24_reg_14_ ( .ck(ispd_clk), .d(n_29470), .o(x_out_24_14) );
ms00f80 x_out_24_reg_15_ ( .ck(ispd_clk), .d(n_29651), .o(x_out_24_15) );
ms00f80 x_out_24_reg_18_ ( .ck(ispd_clk), .d(n_6738), .o(x_out_24_18) );
ms00f80 x_out_24_reg_19_ ( .ck(ispd_clk), .d(n_7329), .o(x_out_24_19) );
ms00f80 x_out_24_reg_1_ ( .ck(ispd_clk), .d(n_19161), .o(x_out_24_1) );
ms00f80 x_out_24_reg_20_ ( .ck(ispd_clk), .d(n_7281), .o(x_out_24_20) );
ms00f80 x_out_24_reg_21_ ( .ck(ispd_clk), .d(n_7310), .o(x_out_24_21) );
ms00f80 x_out_24_reg_22_ ( .ck(ispd_clk), .d(n_7301), .o(x_out_24_22) );
ms00f80 x_out_24_reg_23_ ( .ck(ispd_clk), .d(n_6495), .o(x_out_24_23) );
ms00f80 x_out_24_reg_24_ ( .ck(ispd_clk), .d(n_7305), .o(x_out_24_24) );
ms00f80 x_out_24_reg_25_ ( .ck(ispd_clk), .d(n_7321), .o(x_out_24_25) );
ms00f80 x_out_24_reg_26_ ( .ck(ispd_clk), .d(n_8166), .o(x_out_24_26) );
ms00f80 x_out_24_reg_27_ ( .ck(ispd_clk), .d(n_7337), .o(x_out_24_27) );
ms00f80 x_out_24_reg_28_ ( .ck(ispd_clk), .d(n_7341), .o(x_out_24_28) );
ms00f80 x_out_24_reg_29_ ( .ck(ispd_clk), .d(n_7286), .o(x_out_24_29) );
ms00f80 x_out_24_reg_2_ ( .ck(ispd_clk), .d(n_19839), .o(x_out_24_2) );
ms00f80 x_out_24_reg_30_ ( .ck(ispd_clk), .d(n_7358), .o(x_out_24_30) );
ms00f80 x_out_24_reg_31_ ( .ck(ispd_clk), .d(n_7262), .o(x_out_24_31) );
ms00f80 x_out_24_reg_32_ ( .ck(ispd_clk), .d(n_7256), .o(x_out_24_32) );
ms00f80 x_out_24_reg_33_ ( .ck(ispd_clk), .d(n_5952), .o(x_out_24_33) );
ms00f80 x_out_24_reg_3_ ( .ck(ispd_clk), .d(n_20958), .o(x_out_24_3) );
ms00f80 x_out_24_reg_4_ ( .ck(ispd_clk), .d(n_22068), .o(x_out_24_4) );
ms00f80 x_out_24_reg_5_ ( .ck(ispd_clk), .d(n_23321), .o(x_out_24_5) );
ms00f80 x_out_24_reg_6_ ( .ck(ispd_clk), .d(n_24618), .o(x_out_24_6) );
ms00f80 x_out_24_reg_7_ ( .ck(ispd_clk), .d(n_25898), .o(x_out_24_7) );
ms00f80 x_out_24_reg_8_ ( .ck(ispd_clk), .d(n_26536), .o(x_out_24_8) );
ms00f80 x_out_24_reg_9_ ( .ck(ispd_clk), .d(n_27353), .o(x_out_24_9) );
ms00f80 x_out_25_reg_0_ ( .ck(ispd_clk), .d(n_8685), .o(x_out_25_0) );
ms00f80 x_out_25_reg_10_ ( .ck(ispd_clk), .d(n_26681), .o(x_out_25_10) );
ms00f80 x_out_25_reg_11_ ( .ck(ispd_clk), .d(n_27462), .o(x_out_25_11) );
ms00f80 x_out_25_reg_12_ ( .ck(ispd_clk), .d(n_28127), .o(x_out_25_12) );
ms00f80 x_out_25_reg_13_ ( .ck(ispd_clk), .d(n_28529), .o(x_out_25_13) );
ms00f80 x_out_25_reg_14_ ( .ck(ispd_clk), .d(n_28948), .o(x_out_25_14) );
ms00f80 x_out_25_reg_15_ ( .ck(ispd_clk), .d(n_29306), .o(x_out_25_15) );
ms00f80 x_out_25_reg_18_ ( .ck(ispd_clk), .d(n_7344), .o(x_out_25_18) );
ms00f80 x_out_25_reg_19_ ( .ck(ispd_clk), .d(n_7346), .o(x_out_25_19) );
ms00f80 x_out_25_reg_1_ ( .ck(ispd_clk), .d(n_13770), .o(x_out_25_1) );
ms00f80 x_out_25_reg_20_ ( .ck(ispd_clk), .d(n_7319), .o(x_out_25_20) );
ms00f80 x_out_25_reg_21_ ( .ck(ispd_clk), .d(n_7354), .o(x_out_25_21) );
ms00f80 x_out_25_reg_22_ ( .ck(ispd_clk), .d(n_6501), .o(x_out_25_22) );
ms00f80 x_out_25_reg_23_ ( .ck(ispd_clk), .d(n_7326), .o(x_out_25_23) );
ms00f80 x_out_25_reg_24_ ( .ck(ispd_clk), .d(n_8134), .o(x_out_25_24) );
ms00f80 x_out_25_reg_25_ ( .ck(ispd_clk), .d(n_5775), .o(x_out_25_25) );
ms00f80 x_out_25_reg_26_ ( .ck(ispd_clk), .d(n_7265), .o(x_out_25_26) );
ms00f80 x_out_25_reg_27_ ( .ck(ispd_clk), .d(n_7318), .o(x_out_25_27) );
ms00f80 x_out_25_reg_28_ ( .ck(ispd_clk), .d(n_7371), .o(x_out_25_28) );
ms00f80 x_out_25_reg_29_ ( .ck(ispd_clk), .d(n_7214), .o(x_out_25_29) );
ms00f80 x_out_25_reg_2_ ( .ck(ispd_clk), .d(n_16037), .o(x_out_25_2) );
ms00f80 x_out_25_reg_30_ ( .ck(ispd_clk), .d(n_7425), .o(x_out_25_30) );
ms00f80 x_out_25_reg_31_ ( .ck(ispd_clk), .d(n_7356), .o(x_out_25_31) );
ms00f80 x_out_25_reg_32_ ( .ck(ispd_clk), .d(n_7233), .o(x_out_25_32) );
ms00f80 x_out_25_reg_33_ ( .ck(ispd_clk), .d(n_7238), .o(x_out_25_33) );
ms00f80 x_out_25_reg_3_ ( .ck(ispd_clk), .d(n_19110), .o(x_out_25_3) );
ms00f80 x_out_25_reg_4_ ( .ck(ispd_clk), .d(n_19159), .o(x_out_25_4) );
ms00f80 x_out_25_reg_5_ ( .ck(ispd_clk), .d(n_20538), .o(x_out_25_5) );
ms00f80 x_out_25_reg_6_ ( .ck(ispd_clk), .d(n_22021), .o(x_out_25_6) );
ms00f80 x_out_25_reg_7_ ( .ck(ispd_clk), .d(n_22961), .o(x_out_25_7) );
ms00f80 x_out_25_reg_8_ ( .ck(ispd_clk), .d(n_24207), .o(x_out_25_8) );
ms00f80 x_out_25_reg_9_ ( .ck(ispd_clk), .d(n_25548), .o(x_out_25_9) );
ms00f80 x_out_26_reg_0_ ( .ck(ispd_clk), .d(n_13992), .o(x_out_26_0) );
ms00f80 x_out_26_reg_10_ ( .ck(ispd_clk), .d(n_27704), .o(x_out_26_10) );
ms00f80 x_out_26_reg_11_ ( .ck(ispd_clk), .d(n_28316), .o(x_out_26_11) );
ms00f80 x_out_26_reg_12_ ( .ck(ispd_clk), .d(n_28683), .o(x_out_26_12) );
ms00f80 x_out_26_reg_13_ ( .ck(ispd_clk), .d(n_29038), .o(x_out_26_13) );
ms00f80 x_out_26_reg_14_ ( .ck(ispd_clk), .d(n_29341), .o(x_out_26_14) );
ms00f80 x_out_26_reg_15_ ( .ck(ispd_clk), .d(n_29618), .o(x_out_26_15) );
ms00f80 x_out_26_reg_18_ ( .ck(ispd_clk), .d(n_7345), .o(x_out_26_18) );
ms00f80 x_out_26_reg_19_ ( .ck(ispd_clk), .d(n_6498), .o(x_out_26_19) );
ms00f80 x_out_26_reg_1_ ( .ck(ispd_clk), .d(n_17915), .o(x_out_26_1) );
ms00f80 x_out_26_reg_20_ ( .ck(ispd_clk), .d(n_7276), .o(x_out_26_20) );
ms00f80 x_out_26_reg_21_ ( .ck(ispd_clk), .d(n_7401), .o(x_out_26_21) );
ms00f80 x_out_26_reg_22_ ( .ck(ispd_clk), .d(n_7302), .o(x_out_26_22) );
ms00f80 x_out_26_reg_23_ ( .ck(ispd_clk), .d(n_7374), .o(x_out_26_23) );
ms00f80 x_out_26_reg_24_ ( .ck(ispd_clk), .d(n_7271), .o(x_out_26_24) );
ms00f80 x_out_26_reg_25_ ( .ck(ispd_clk), .d(n_7368), .o(x_out_26_25) );
ms00f80 x_out_26_reg_26_ ( .ck(ispd_clk), .d(n_6456), .o(x_out_26_26) );
ms00f80 x_out_26_reg_27_ ( .ck(ispd_clk), .d(n_7297), .o(x_out_26_27) );
ms00f80 x_out_26_reg_28_ ( .ck(ispd_clk), .d(n_7324), .o(x_out_26_28) );
ms00f80 x_out_26_reg_29_ ( .ck(ispd_clk), .d(n_6489), .o(x_out_26_29) );
ms00f80 x_out_26_reg_2_ ( .ck(ispd_clk), .d(n_18528), .o(x_out_26_2) );
ms00f80 x_out_26_reg_30_ ( .ck(ispd_clk), .d(n_7293), .o(x_out_26_30) );
ms00f80 x_out_26_reg_31_ ( .ck(ispd_clk), .d(n_8205), .o(x_out_26_31) );
ms00f80 x_out_26_reg_32_ ( .ck(ispd_clk), .d(n_7259), .o(x_out_26_32) );
ms00f80 x_out_26_reg_33_ ( .ck(ispd_clk), .d(n_7252), .o(x_out_26_33) );
ms00f80 x_out_26_reg_3_ ( .ck(ispd_clk), .d(n_20890), .o(x_out_26_3) );
ms00f80 x_out_26_reg_4_ ( .ck(ispd_clk), .d(n_20972), .o(x_out_26_4) );
ms00f80 x_out_26_reg_5_ ( .ck(ispd_clk), .d(n_22065), .o(x_out_26_5) );
ms00f80 x_out_26_reg_6_ ( .ck(ispd_clk), .d(n_23316), .o(x_out_26_6) );
ms00f80 x_out_26_reg_7_ ( .ck(ispd_clk), .d(n_24614), .o(x_out_26_7) );
ms00f80 x_out_26_reg_8_ ( .ck(ispd_clk), .d(n_25894), .o(x_out_26_8) );
ms00f80 x_out_26_reg_9_ ( .ck(ispd_clk), .d(n_26803), .o(x_out_26_9) );
ms00f80 x_out_27_reg_0_ ( .ck(ispd_clk), .d(n_13877), .o(x_out_27_0) );
ms00f80 x_out_27_reg_10_ ( .ck(ispd_clk), .d(n_27701), .o(x_out_27_10) );
ms00f80 x_out_27_reg_11_ ( .ck(ispd_clk), .d(n_28312), .o(x_out_27_11) );
ms00f80 x_out_27_reg_12_ ( .ck(ispd_clk), .d(n_28681), .o(x_out_27_12) );
ms00f80 x_out_27_reg_13_ ( .ck(ispd_clk), .d(n_29035), .o(x_out_27_13) );
ms00f80 x_out_27_reg_14_ ( .ck(ispd_clk), .d(n_29338), .o(x_out_27_14) );
ms00f80 x_out_27_reg_15_ ( .ck(ispd_clk), .d(n_29616), .o(x_out_27_15) );
ms00f80 x_out_27_reg_18_ ( .ck(ispd_clk), .d(n_7365), .o(x_out_27_18) );
ms00f80 x_out_27_reg_19_ ( .ck(ispd_clk), .d(n_6486), .o(x_out_27_19) );
ms00f80 x_out_27_reg_1_ ( .ck(ispd_clk), .d(n_17927), .o(x_out_27_1) );
ms00f80 x_out_27_reg_20_ ( .ck(ispd_clk), .d(n_7327), .o(x_out_27_20) );
ms00f80 x_out_27_reg_21_ ( .ck(ispd_clk), .d(n_8038), .o(x_out_27_21) );
ms00f80 x_out_27_reg_22_ ( .ck(ispd_clk), .d(n_7280), .o(x_out_27_22) );
ms00f80 x_out_27_reg_23_ ( .ck(ispd_clk), .d(n_7376), .o(x_out_27_23) );
ms00f80 x_out_27_reg_24_ ( .ck(ispd_clk), .d(n_7316), .o(x_out_27_24) );
ms00f80 x_out_27_reg_25_ ( .ck(ispd_clk), .d(n_7363), .o(x_out_27_25) );
ms00f80 x_out_27_reg_26_ ( .ck(ispd_clk), .d(n_7282), .o(x_out_27_26) );
ms00f80 x_out_27_reg_27_ ( .ck(ispd_clk), .d(n_7333), .o(x_out_27_27) );
ms00f80 x_out_27_reg_28_ ( .ck(ispd_clk), .d(n_7279), .o(x_out_27_28) );
ms00f80 x_out_27_reg_29_ ( .ck(ispd_clk), .d(n_7232), .o(x_out_27_29) );
ms00f80 x_out_27_reg_2_ ( .ck(ispd_clk), .d(n_18527), .o(x_out_27_2) );
ms00f80 x_out_27_reg_30_ ( .ck(ispd_clk), .d(n_8002), .o(x_out_27_30) );
ms00f80 x_out_27_reg_31_ ( .ck(ispd_clk), .d(n_7362), .o(x_out_27_31) );
ms00f80 x_out_27_reg_32_ ( .ck(ispd_clk), .d(n_5776), .o(x_out_27_32) );
ms00f80 x_out_27_reg_33_ ( .ck(ispd_clk), .d(n_7249), .o(x_out_27_33) );
ms00f80 x_out_27_reg_3_ ( .ck(ispd_clk), .d(n_20889), .o(x_out_27_3) );
ms00f80 x_out_27_reg_4_ ( .ck(ispd_clk), .d(n_20971), .o(x_out_27_4) );
ms00f80 x_out_27_reg_5_ ( .ck(ispd_clk), .d(n_22059), .o(x_out_27_5) );
ms00f80 x_out_27_reg_6_ ( .ck(ispd_clk), .d(n_23310), .o(x_out_27_6) );
ms00f80 x_out_27_reg_7_ ( .ck(ispd_clk), .d(n_24613), .o(x_out_27_7) );
ms00f80 x_out_27_reg_8_ ( .ck(ispd_clk), .d(n_25904), .o(x_out_27_8) );
ms00f80 x_out_27_reg_9_ ( .ck(ispd_clk), .d(n_26799), .o(x_out_27_9) );
ms00f80 x_out_28_reg_0_ ( .ck(ispd_clk), .d(n_13989), .o(x_out_28_0) );
ms00f80 x_out_28_reg_10_ ( .ck(ispd_clk), .d(n_27351), .o(x_out_28_10) );
ms00f80 x_out_28_reg_11_ ( .ck(ispd_clk), .d(n_28087), .o(x_out_28_11) );
ms00f80 x_out_28_reg_12_ ( .ck(ispd_clk), .d(n_28484), .o(x_out_28_12) );
ms00f80 x_out_28_reg_13_ ( .ck(ispd_clk), .d(n_28827), .o(x_out_28_13) );
ms00f80 x_out_28_reg_14_ ( .ck(ispd_clk), .d(n_29175), .o(x_out_28_14) );
ms00f80 x_out_28_reg_15_ ( .ck(ispd_clk), .d(n_29498), .o(x_out_28_15) );
ms00f80 x_out_28_reg_18_ ( .ck(ispd_clk), .d(n_7378), .o(x_out_28_18) );
ms00f80 x_out_28_reg_19_ ( .ck(ispd_clk), .d(n_7314), .o(x_out_28_19) );
ms00f80 x_out_28_reg_1_ ( .ck(ispd_clk), .d(n_17926), .o(x_out_28_1) );
ms00f80 x_out_28_reg_20_ ( .ck(ispd_clk), .d(n_6499), .o(x_out_28_20) );
ms00f80 x_out_28_reg_21_ ( .ck(ispd_clk), .d(n_5785), .o(x_out_28_21) );
ms00f80 x_out_28_reg_22_ ( .ck(ispd_clk), .d(n_7370), .o(x_out_28_22) );
ms00f80 x_out_28_reg_23_ ( .ck(ispd_clk), .d(n_7375), .o(x_out_28_23) );
ms00f80 x_out_28_reg_24_ ( .ck(ispd_clk), .d(n_6493), .o(x_out_28_24) );
ms00f80 x_out_28_reg_25_ ( .ck(ispd_clk), .d(n_7355), .o(x_out_28_25) );
ms00f80 x_out_28_reg_26_ ( .ck(ispd_clk), .d(n_7294), .o(x_out_28_26) );
ms00f80 x_out_28_reg_27_ ( .ck(ispd_clk), .d(n_7335), .o(x_out_28_27) );
ms00f80 x_out_28_reg_28_ ( .ck(ispd_clk), .d(n_7339), .o(x_out_28_28) );
ms00f80 x_out_28_reg_29_ ( .ck(ispd_clk), .d(n_8005), .o(x_out_28_29) );
ms00f80 x_out_28_reg_2_ ( .ck(ispd_clk), .d(n_18524), .o(x_out_28_2) );
ms00f80 x_out_28_reg_30_ ( .ck(ispd_clk), .d(n_7372), .o(x_out_28_30) );
ms00f80 x_out_28_reg_31_ ( .ck(ispd_clk), .d(n_6430), .o(x_out_28_31) );
ms00f80 x_out_28_reg_32_ ( .ck(ispd_clk), .d(n_8057), .o(x_out_28_32) );
ms00f80 x_out_28_reg_33_ ( .ck(ispd_clk), .d(n_5787), .o(x_out_28_33) );
ms00f80 x_out_28_reg_3_ ( .ck(ispd_clk), .d(n_20888), .o(x_out_28_3) );
ms00f80 x_out_28_reg_4_ ( .ck(ispd_clk), .d(n_20968), .o(x_out_28_4) );
ms00f80 x_out_28_reg_5_ ( .ck(ispd_clk), .d(n_22063), .o(x_out_28_5) );
ms00f80 x_out_28_reg_6_ ( .ck(ispd_clk), .d(n_23307), .o(x_out_28_6) );
ms00f80 x_out_28_reg_7_ ( .ck(ispd_clk), .d(n_24610), .o(x_out_28_7) );
ms00f80 x_out_28_reg_8_ ( .ck(ispd_clk), .d(n_25668), .o(x_out_28_8) );
ms00f80 x_out_28_reg_9_ ( .ck(ispd_clk), .d(n_26237), .o(x_out_28_9) );
ms00f80 x_out_29_reg_0_ ( .ck(ispd_clk), .d(n_14748), .o(x_out_29_0) );
ms00f80 x_out_29_reg_10_ ( .ck(ispd_clk), .d(n_27699), .o(x_out_29_10) );
ms00f80 x_out_29_reg_11_ ( .ck(ispd_clk), .d(n_28308), .o(x_out_29_11) );
ms00f80 x_out_29_reg_12_ ( .ck(ispd_clk), .d(n_28680), .o(x_out_29_12) );
ms00f80 x_out_29_reg_13_ ( .ck(ispd_clk), .d(n_29034), .o(x_out_29_13) );
ms00f80 x_out_29_reg_14_ ( .ck(ispd_clk), .d(n_29408), .o(x_out_29_14) );
ms00f80 x_out_29_reg_15_ ( .ck(ispd_clk), .d(n_29611), .o(x_out_29_15) );
ms00f80 x_out_29_reg_18_ ( .ck(ispd_clk), .d(n_7255), .o(x_out_29_18) );
ms00f80 x_out_29_reg_19_ ( .ck(ispd_clk), .d(n_7234), .o(x_out_29_19) );
ms00f80 x_out_29_reg_1_ ( .ck(ispd_clk), .d(n_17925), .o(x_out_29_1) );
ms00f80 x_out_29_reg_20_ ( .ck(ispd_clk), .d(n_7235), .o(x_out_29_20) );
ms00f80 x_out_29_reg_21_ ( .ck(ispd_clk), .d(n_7377), .o(x_out_29_21) );
ms00f80 x_out_29_reg_22_ ( .ck(ispd_clk), .d(n_7236), .o(x_out_29_22) );
ms00f80 x_out_29_reg_23_ ( .ck(ispd_clk), .d(n_7379), .o(x_out_29_23) );
ms00f80 x_out_29_reg_24_ ( .ck(ispd_clk), .d(n_7242), .o(x_out_29_24) );
ms00f80 x_out_29_reg_25_ ( .ck(ispd_clk), .d(n_7388), .o(x_out_29_25) );
ms00f80 x_out_29_reg_26_ ( .ck(ispd_clk), .d(n_7244), .o(x_out_29_26) );
ms00f80 x_out_29_reg_27_ ( .ck(ispd_clk), .d(n_7246), .o(x_out_29_27) );
ms00f80 x_out_29_reg_28_ ( .ck(ispd_clk), .d(n_7248), .o(x_out_29_28) );
ms00f80 x_out_29_reg_29_ ( .ck(ispd_clk), .d(n_7392), .o(x_out_29_29) );
ms00f80 x_out_29_reg_2_ ( .ck(ispd_clk), .d(n_18800), .o(x_out_29_2) );
ms00f80 x_out_29_reg_30_ ( .ck(ispd_clk), .d(n_6490), .o(x_out_29_30) );
ms00f80 x_out_29_reg_31_ ( .ck(ispd_clk), .d(n_6094), .o(x_out_29_31) );
ms00f80 x_out_29_reg_32_ ( .ck(ispd_clk), .d(n_7393), .o(x_out_29_32) );
ms00f80 x_out_29_reg_33_ ( .ck(ispd_clk), .d(n_7407), .o(x_out_29_33) );
ms00f80 x_out_29_reg_3_ ( .ck(ispd_clk), .d(n_20887), .o(x_out_29_3) );
ms00f80 x_out_29_reg_4_ ( .ck(ispd_clk), .d(n_20967), .o(x_out_29_4) );
ms00f80 x_out_29_reg_5_ ( .ck(ispd_clk), .d(n_22062), .o(x_out_29_5) );
ms00f80 x_out_29_reg_6_ ( .ck(ispd_clk), .d(n_23306), .o(x_out_29_6) );
ms00f80 x_out_29_reg_7_ ( .ck(ispd_clk), .d(n_24609), .o(x_out_29_7) );
ms00f80 x_out_29_reg_8_ ( .ck(ispd_clk), .d(n_25889), .o(x_out_29_8) );
ms00f80 x_out_29_reg_9_ ( .ck(ispd_clk), .d(n_26790), .o(x_out_29_9) );
ms00f80 x_out_2_reg_0_ ( .ck(ispd_clk), .d(n_15542), .o(x_out_2_0) );
ms00f80 x_out_2_reg_10_ ( .ck(ispd_clk), .d(n_27549), .o(x_out_2_10) );
ms00f80 x_out_2_reg_11_ ( .ck(ispd_clk), .d(n_28209), .o(x_out_2_11) );
ms00f80 x_out_2_reg_12_ ( .ck(ispd_clk), .d(n_28602), .o(x_out_2_12) );
ms00f80 x_out_2_reg_13_ ( .ck(ispd_clk), .d(n_28913), .o(x_out_2_13) );
ms00f80 x_out_2_reg_14_ ( .ck(ispd_clk), .d(n_29337), .o(x_out_2_14) );
ms00f80 x_out_2_reg_15_ ( .ck(ispd_clk), .d(n_29561), .o(x_out_2_15) );
ms00f80 x_out_2_reg_18_ ( .ck(ispd_clk), .d(n_11416), .o(x_out_2_18) );
ms00f80 x_out_2_reg_19_ ( .ck(ispd_clk), .d(n_16371), .o(x_out_2_19) );
ms00f80 x_out_2_reg_1_ ( .ck(ispd_clk), .d(n_17701), .o(x_out_2_1) );
ms00f80 x_out_2_reg_20_ ( .ck(ispd_clk), .d(n_16009), .o(x_out_2_20) );
ms00f80 x_out_2_reg_21_ ( .ck(ispd_clk), .d(n_16433), .o(x_out_2_21) );
ms00f80 x_out_2_reg_22_ ( .ck(ispd_clk), .d(n_16754), .o(x_out_2_22) );
ms00f80 x_out_2_reg_23_ ( .ck(ispd_clk), .d(n_17924), .o(x_out_2_23) );
ms00f80 x_out_2_reg_24_ ( .ck(ispd_clk), .d(n_18576), .o(x_out_2_24) );
ms00f80 x_out_2_reg_25_ ( .ck(ispd_clk), .d(n_19892), .o(x_out_2_25) );
ms00f80 x_out_2_reg_26_ ( .ck(ispd_clk), .d(n_20703), .o(x_out_2_26) );
ms00f80 x_out_2_reg_27_ ( .ck(ispd_clk), .d(n_21811), .o(x_out_2_27) );
ms00f80 x_out_2_reg_28_ ( .ck(ispd_clk), .d(n_22467), .o(x_out_2_28) );
ms00f80 x_out_2_reg_29_ ( .ck(ispd_clk), .d(n_23716), .o(x_out_2_29) );
ms00f80 x_out_2_reg_2_ ( .ck(ispd_clk), .d(n_18798), .o(x_out_2_2) );
ms00f80 x_out_2_reg_30_ ( .ck(ispd_clk), .d(n_24402), .o(x_out_2_30) );
ms00f80 x_out_2_reg_31_ ( .ck(ispd_clk), .d(n_25427), .o(x_out_2_31) );
ms00f80 x_out_2_reg_32_ ( .ck(ispd_clk), .d(n_26331), .o(x_out_2_32) );
ms00f80 x_out_2_reg_33_ ( .ck(ispd_clk), .d(n_26330), .o(x_out_2_33) );
ms00f80 x_out_2_reg_3_ ( .ck(ispd_clk), .d(n_20182), .o(x_out_2_3) );
ms00f80 x_out_2_reg_4_ ( .ck(ispd_clk), .d(n_20966), .o(x_out_2_4) );
ms00f80 x_out_2_reg_5_ ( .ck(ispd_clk), .d(n_21767), .o(x_out_2_5) );
ms00f80 x_out_2_reg_6_ ( .ck(ispd_clk), .d(n_23050), .o(x_out_2_6) );
ms00f80 x_out_2_reg_7_ ( .ck(ispd_clk), .d(n_24297), .o(x_out_2_7) );
ms00f80 x_out_2_reg_8_ ( .ck(ispd_clk), .d(n_25666), .o(x_out_2_8) );
ms00f80 x_out_2_reg_9_ ( .ck(ispd_clk), .d(n_26523), .o(x_out_2_9) );
ms00f80 x_out_30_reg_0_ ( .ck(ispd_clk), .d(n_14721), .o(x_out_30_0) );
ms00f80 x_out_30_reg_10_ ( .ck(ispd_clk), .d(n_27698), .o(x_out_30_10) );
ms00f80 x_out_30_reg_11_ ( .ck(ispd_clk), .d(n_28306), .o(x_out_30_11) );
ms00f80 x_out_30_reg_12_ ( .ck(ispd_clk), .d(n_28679), .o(x_out_30_12) );
ms00f80 x_out_30_reg_13_ ( .ck(ispd_clk), .d(n_29031), .o(x_out_30_13) );
ms00f80 x_out_30_reg_14_ ( .ck(ispd_clk), .d(n_29406), .o(x_out_30_14) );
ms00f80 x_out_30_reg_15_ ( .ck(ispd_clk), .d(n_29608), .o(x_out_30_15) );
ms00f80 x_out_30_reg_18_ ( .ck(ispd_clk), .d(n_7447), .o(x_out_30_18) );
ms00f80 x_out_30_reg_19_ ( .ck(ispd_clk), .d(n_8202), .o(x_out_30_19) );
ms00f80 x_out_30_reg_1_ ( .ck(ispd_clk), .d(n_17923), .o(x_out_30_1) );
ms00f80 x_out_30_reg_20_ ( .ck(ispd_clk), .d(n_7300), .o(x_out_30_20) );
ms00f80 x_out_30_reg_21_ ( .ck(ispd_clk), .d(n_7352), .o(x_out_30_21) );
ms00f80 x_out_30_reg_22_ ( .ck(ispd_clk), .d(n_6484), .o(x_out_30_22) );
ms00f80 x_out_30_reg_23_ ( .ck(ispd_clk), .d(n_6401), .o(x_out_30_23) );
ms00f80 x_out_30_reg_24_ ( .ck(ispd_clk), .d(n_8201), .o(x_out_30_24) );
ms00f80 x_out_30_reg_25_ ( .ck(ispd_clk), .d(n_8009), .o(x_out_30_25) );
ms00f80 x_out_30_reg_26_ ( .ck(ispd_clk), .d(n_7313), .o(x_out_30_26) );
ms00f80 x_out_30_reg_27_ ( .ck(ispd_clk), .d(n_7299), .o(x_out_30_27) );
ms00f80 x_out_30_reg_28_ ( .ck(ispd_clk), .d(n_6487), .o(x_out_30_28) );
ms00f80 x_out_30_reg_29_ ( .ck(ispd_clk), .d(n_7292), .o(x_out_30_29) );
ms00f80 x_out_30_reg_2_ ( .ck(ispd_clk), .d(n_19109), .o(x_out_30_2) );
ms00f80 x_out_30_reg_30_ ( .ck(ispd_clk), .d(n_7353), .o(x_out_30_30) );
ms00f80 x_out_30_reg_31_ ( .ck(ispd_clk), .d(n_6408), .o(x_out_30_31) );
ms00f80 x_out_30_reg_32_ ( .ck(ispd_clk), .d(n_7576), .o(x_out_30_32) );
ms00f80 x_out_30_reg_33_ ( .ck(ispd_clk), .d(n_7574), .o(x_out_30_33) );
ms00f80 x_out_30_reg_3_ ( .ck(ispd_clk), .d(n_20886), .o(x_out_30_3) );
ms00f80 x_out_30_reg_4_ ( .ck(ispd_clk), .d(n_20965), .o(x_out_30_4) );
ms00f80 x_out_30_reg_5_ ( .ck(ispd_clk), .d(n_22061), .o(x_out_30_5) );
ms00f80 x_out_30_reg_6_ ( .ck(ispd_clk), .d(n_23305), .o(x_out_30_6) );
ms00f80 x_out_30_reg_7_ ( .ck(ispd_clk), .d(n_24608), .o(x_out_30_7) );
ms00f80 x_out_30_reg_8_ ( .ck(ispd_clk), .d(n_25888), .o(x_out_30_8) );
ms00f80 x_out_30_reg_9_ ( .ck(ispd_clk), .d(n_26785), .o(x_out_30_9) );
ms00f80 x_out_31_reg_0_ ( .ck(ispd_clk), .d(n_14695), .o(x_out_31_0) );
ms00f80 x_out_31_reg_10_ ( .ck(ispd_clk), .d(n_27696), .o(x_out_31_10) );
ms00f80 x_out_31_reg_11_ ( .ck(ispd_clk), .d(n_28304), .o(x_out_31_11) );
ms00f80 x_out_31_reg_12_ ( .ck(ispd_clk), .d(n_28678), .o(x_out_31_12) );
ms00f80 x_out_31_reg_13_ ( .ck(ispd_clk), .d(n_29030), .o(x_out_31_13) );
ms00f80 x_out_31_reg_14_ ( .ck(ispd_clk), .d(n_29404), .o(x_out_31_14) );
ms00f80 x_out_31_reg_15_ ( .ck(ispd_clk), .d(n_29606), .o(x_out_31_15) );
ms00f80 x_out_31_reg_18_ ( .ck(ispd_clk), .d(n_7394), .o(x_out_31_18) );
ms00f80 x_out_31_reg_19_ ( .ck(ispd_clk), .d(n_7322), .o(x_out_31_19) );
ms00f80 x_out_31_reg_1_ ( .ck(ispd_clk), .d(n_17922), .o(x_out_31_1) );
ms00f80 x_out_31_reg_20_ ( .ck(ispd_clk), .d(n_6479), .o(x_out_31_20) );
ms00f80 x_out_31_reg_21_ ( .ck(ispd_clk), .d(n_7258), .o(x_out_31_21) );
ms00f80 x_out_31_reg_22_ ( .ck(ispd_clk), .d(n_7267), .o(x_out_31_22) );
ms00f80 x_out_31_reg_23_ ( .ck(ispd_clk), .d(n_8203), .o(x_out_31_23) );
ms00f80 x_out_31_reg_24_ ( .ck(ispd_clk), .d(n_7273), .o(x_out_31_24) );
ms00f80 x_out_31_reg_25_ ( .ck(ispd_clk), .d(n_7351), .o(x_out_31_25) );
ms00f80 x_out_31_reg_26_ ( .ck(ispd_clk), .d(n_7295), .o(x_out_31_26) );
ms00f80 x_out_31_reg_27_ ( .ck(ispd_clk), .d(n_7309), .o(x_out_31_27) );
ms00f80 x_out_31_reg_28_ ( .ck(ispd_clk), .d(n_8207), .o(x_out_31_28) );
ms00f80 x_out_31_reg_29_ ( .ck(ispd_clk), .d(n_8007), .o(x_out_31_29) );
ms00f80 x_out_31_reg_2_ ( .ck(ispd_clk), .d(n_18522), .o(x_out_31_2) );
ms00f80 x_out_31_reg_30_ ( .ck(ispd_clk), .d(n_7343), .o(x_out_31_30) );
ms00f80 x_out_31_reg_31_ ( .ck(ispd_clk), .d(n_8199), .o(x_out_31_31) );
ms00f80 x_out_31_reg_32_ ( .ck(ispd_clk), .d(n_7306), .o(x_out_31_32) );
ms00f80 x_out_31_reg_33_ ( .ck(ispd_clk), .d(n_5971), .o(x_out_31_33) );
ms00f80 x_out_31_reg_3_ ( .ck(ispd_clk), .d(n_20885), .o(x_out_31_3) );
ms00f80 x_out_31_reg_4_ ( .ck(ispd_clk), .d(n_20964), .o(x_out_31_4) );
ms00f80 x_out_31_reg_5_ ( .ck(ispd_clk), .d(n_22060), .o(x_out_31_5) );
ms00f80 x_out_31_reg_6_ ( .ck(ispd_clk), .d(n_23302), .o(x_out_31_6) );
ms00f80 x_out_31_reg_7_ ( .ck(ispd_clk), .d(n_24606), .o(x_out_31_7) );
ms00f80 x_out_31_reg_8_ ( .ck(ispd_clk), .d(n_25887), .o(x_out_31_8) );
ms00f80 x_out_31_reg_9_ ( .ck(ispd_clk), .d(n_26783), .o(x_out_31_9) );
ms00f80 x_out_32_reg_0_ ( .ck(ispd_clk), .d(n_7412), .o(x_out_32_0) );
ms00f80 x_out_32_reg_10_ ( .ck(ispd_clk), .d(n_22377), .o(x_out_32_10) );
ms00f80 x_out_32_reg_11_ ( .ck(ispd_clk), .d(n_23655), .o(x_out_32_11) );
ms00f80 x_out_32_reg_12_ ( .ck(ispd_clk), .d(n_24985), .o(x_out_32_12) );
ms00f80 x_out_32_reg_13_ ( .ck(ispd_clk), .d(n_26183), .o(x_out_32_13) );
ms00f80 x_out_32_reg_14_ ( .ck(ispd_clk), .d(n_27076), .o(x_out_32_14) );
ms00f80 x_out_32_reg_15_ ( .ck(ispd_clk), .d(n_27891), .o(x_out_32_15) );
ms00f80 x_out_32_reg_1_ ( .ck(ispd_clk), .d(n_11024), .o(x_out_32_1) );
ms00f80 x_out_32_reg_2_ ( .ck(ispd_clk), .d(n_12571), .o(x_out_32_2) );
ms00f80 x_out_32_reg_3_ ( .ck(ispd_clk), .d(n_14130), .o(x_out_32_3) );
ms00f80 x_out_32_reg_4_ ( .ck(ispd_clk), .d(n_14591), .o(x_out_32_4) );
ms00f80 x_out_32_reg_5_ ( .ck(ispd_clk), .d(n_16292), .o(x_out_32_5) );
ms00f80 x_out_32_reg_6_ ( .ck(ispd_clk), .d(n_17421), .o(x_out_32_6) );
ms00f80 x_out_32_reg_7_ ( .ck(ispd_clk), .d(n_18574), .o(x_out_32_7) );
ms00f80 x_out_32_reg_8_ ( .ck(ispd_clk), .d(n_19890), .o(x_out_32_8) );
ms00f80 x_out_32_reg_9_ ( .ck(ispd_clk), .d(n_21325), .o(x_out_32_9) );
ms00f80 x_out_33_reg_0_ ( .ck(ispd_clk), .d(n_16794), .o(x_out_33_0) );
ms00f80 x_out_33_reg_10_ ( .ck(ispd_clk), .d(n_28263), .o(x_out_33_10) );
ms00f80 x_out_33_reg_11_ ( .ck(ispd_clk), .d(n_28652), .o(x_out_33_11) );
ms00f80 x_out_33_reg_12_ ( .ck(ispd_clk), .d(n_29100), .o(x_out_33_12) );
ms00f80 x_out_33_reg_13_ ( .ck(ispd_clk), .d(n_29353), .o(x_out_33_13) );
ms00f80 x_out_33_reg_14_ ( .ck(ispd_clk), .d(n_29584), .o(x_out_33_14) );
ms00f80 x_out_33_reg_15_ ( .ck(ispd_clk), .d(n_29662), .o(x_out_33_15) );
ms00f80 x_out_33_reg_18_ ( .ck(ispd_clk), .d(n_14209), .o(x_out_33_18) );
ms00f80 x_out_33_reg_19_ ( .ck(ispd_clk), .d(n_17224), .o(x_out_33_19) );
ms00f80 x_out_33_reg_1_ ( .ck(ispd_clk), .d(n_19833), .o(x_out_33_1) );
ms00f80 x_out_33_reg_20_ ( .ck(ispd_clk), .d(n_17373), .o(x_out_33_20) );
ms00f80 x_out_33_reg_21_ ( .ck(ispd_clk), .d(n_18013), .o(x_out_33_21) );
ms00f80 x_out_33_reg_22_ ( .ck(ispd_clk), .d(n_18987), .o(x_out_33_22) );
ms00f80 x_out_33_reg_23_ ( .ck(ispd_clk), .d(n_19993), .o(x_out_33_23) );
ms00f80 x_out_33_reg_24_ ( .ck(ispd_clk), .d(n_20440), .o(x_out_33_24) );
ms00f80 x_out_33_reg_25_ ( .ck(ispd_clk), .d(n_21903), .o(x_out_33_25) );
ms00f80 x_out_33_reg_26_ ( .ck(ispd_clk), .d(n_22552), .o(x_out_33_26) );
ms00f80 x_out_33_reg_27_ ( .ck(ispd_clk), .d(n_23810), .o(x_out_33_27) );
ms00f80 x_out_33_reg_28_ ( .ck(ispd_clk), .d(n_24178), .o(x_out_33_28) );
ms00f80 x_out_33_reg_29_ ( .ck(ispd_clk), .d(n_25522), .o(x_out_33_29) );
ms00f80 x_out_33_reg_2_ ( .ck(ispd_clk), .d(n_21265), .o(x_out_33_2) );
ms00f80 x_out_33_reg_30_ ( .ck(ispd_clk), .d(n_26051), .o(x_out_33_30) );
ms00f80 x_out_33_reg_31_ ( .ck(ispd_clk), .d(n_26566), .o(x_out_33_31) );
ms00f80 x_out_33_reg_32_ ( .ck(ispd_clk), .d(n_26562), .o(x_out_33_32) );
ms00f80 x_out_33_reg_33_ ( .ck(ispd_clk), .d(n_26564), .o(x_out_33_33) );
ms00f80 x_out_33_reg_3_ ( .ck(ispd_clk), .d(n_22610), .o(x_out_33_3) );
ms00f80 x_out_33_reg_4_ ( .ck(ispd_clk), .d(n_23611), .o(x_out_33_4) );
ms00f80 x_out_33_reg_5_ ( .ck(ispd_clk), .d(n_24605), .o(x_out_33_5) );
ms00f80 x_out_33_reg_6_ ( .ck(ispd_clk), .d(n_25355), .o(x_out_33_6) );
ms00f80 x_out_33_reg_7_ ( .ck(ispd_clk), .d(n_26233), .o(x_out_33_7) );
ms00f80 x_out_33_reg_8_ ( .ck(ispd_clk), .d(n_27152), .o(x_out_33_8) );
ms00f80 x_out_33_reg_9_ ( .ck(ispd_clk), .d(n_27791), .o(x_out_33_9) );
ms00f80 x_out_34_reg_0_ ( .ck(ispd_clk), .d(n_15535), .o(x_out_34_0) );
ms00f80 x_out_34_reg_10_ ( .ck(ispd_clk), .d(n_28085), .o(x_out_34_10) );
ms00f80 x_out_34_reg_11_ ( .ck(ispd_clk), .d(n_28480), .o(x_out_34_11) );
ms00f80 x_out_34_reg_12_ ( .ck(ispd_clk), .d(n_28821), .o(x_out_34_12) );
ms00f80 x_out_34_reg_13_ ( .ck(ispd_clk), .d(n_29251), .o(x_out_34_13) );
ms00f80 x_out_34_reg_14_ ( .ck(ispd_clk), .d(n_29465), .o(x_out_34_14) );
ms00f80 x_out_34_reg_15_ ( .ck(ispd_clk), .d(n_29660), .o(x_out_34_15) );
ms00f80 x_out_34_reg_18_ ( .ck(ispd_clk), .d(n_11414), .o(x_out_34_18) );
ms00f80 x_out_34_reg_19_ ( .ck(ispd_clk), .d(n_17515), .o(x_out_34_19) );
ms00f80 x_out_34_reg_1_ ( .ck(ispd_clk), .d(n_19152), .o(x_out_34_1) );
ms00f80 x_out_34_reg_20_ ( .ck(ispd_clk), .d(n_17844), .o(x_out_34_20) );
ms00f80 x_out_34_reg_21_ ( .ck(ispd_clk), .d(n_18410), .o(x_out_34_21) );
ms00f80 x_out_34_reg_22_ ( .ck(ispd_clk), .d(n_19108), .o(x_out_34_22) );
ms00f80 x_out_34_reg_23_ ( .ck(ispd_clk), .d(n_19748), .o(x_out_34_23) );
ms00f80 x_out_34_reg_24_ ( .ck(ispd_clk), .d(n_20536), .o(x_out_34_24) );
ms00f80 x_out_34_reg_25_ ( .ck(ispd_clk), .d(n_21324), .o(x_out_34_25) );
ms00f80 x_out_34_reg_26_ ( .ck(ispd_clk), .d(n_22106), .o(x_out_34_26) );
ms00f80 x_out_34_reg_27_ ( .ck(ispd_clk), .d(n_23078), .o(x_out_34_27) );
ms00f80 x_out_34_reg_28_ ( .ck(ispd_clk), .d(n_24037), .o(x_out_34_28) );
ms00f80 x_out_34_reg_29_ ( .ck(ispd_clk), .d(n_25036), .o(x_out_34_29) );
ms00f80 x_out_34_reg_2_ ( .ck(ispd_clk), .d(n_20181), .o(x_out_34_2) );
ms00f80 x_out_34_reg_30_ ( .ck(ispd_clk), .d(n_25741), .o(x_out_34_30) );
ms00f80 x_out_34_reg_31_ ( .ck(ispd_clk), .d(n_26311), .o(x_out_34_31) );
ms00f80 x_out_34_reg_32_ ( .ck(ispd_clk), .d(n_26635), .o(x_out_34_32) );
ms00f80 x_out_34_reg_33_ ( .ck(ispd_clk), .d(n_26634), .o(x_out_34_33) );
ms00f80 x_out_34_reg_3_ ( .ck(ispd_clk), .d(n_21602), .o(x_out_34_3) );
ms00f80 x_out_34_reg_4_ ( .ck(ispd_clk), .d(n_22309), .o(x_out_34_4) );
ms00f80 x_out_34_reg_5_ ( .ck(ispd_clk), .d(n_23301), .o(x_out_34_5) );
ms00f80 x_out_34_reg_6_ ( .ck(ispd_clk), .d(n_24295), .o(x_out_34_6) );
ms00f80 x_out_34_reg_7_ ( .ck(ispd_clk), .d(n_25353), .o(x_out_34_7) );
ms00f80 x_out_34_reg_8_ ( .ck(ispd_clk), .d(n_26231), .o(x_out_34_8) );
ms00f80 x_out_34_reg_9_ ( .ck(ispd_clk), .d(n_27349), .o(x_out_34_9) );
ms00f80 x_out_35_reg_0_ ( .ck(ispd_clk), .d(n_16980), .o(x_out_35_0) );
ms00f80 x_out_35_reg_10_ ( .ck(ispd_clk), .d(n_28478), .o(x_out_35_10) );
ms00f80 x_out_35_reg_11_ ( .ck(ispd_clk), .d(n_28819), .o(x_out_35_11) );
ms00f80 x_out_35_reg_12_ ( .ck(ispd_clk), .d(n_29250), .o(x_out_35_12) );
ms00f80 x_out_35_reg_13_ ( .ck(ispd_clk), .d(n_29464), .o(x_out_35_13) );
ms00f80 x_out_35_reg_14_ ( .ck(ispd_clk), .d(n_29644), .o(x_out_35_14) );
ms00f80 x_out_35_reg_15_ ( .ck(ispd_clk), .d(n_29695), .o(x_out_35_15) );
ms00f80 x_out_35_reg_18_ ( .ck(ispd_clk), .d(n_10720), .o(x_out_35_18) );
ms00f80 x_out_35_reg_19_ ( .ck(ispd_clk), .d(n_16775), .o(x_out_35_19) );
ms00f80 x_out_35_reg_1_ ( .ck(ispd_clk), .d(n_19832), .o(x_out_35_1) );
ms00f80 x_out_35_reg_20_ ( .ck(ispd_clk), .d(n_17372), .o(x_out_35_20) );
ms00f80 x_out_35_reg_21_ ( .ck(ispd_clk), .d(n_17920), .o(x_out_35_21) );
ms00f80 x_out_35_reg_22_ ( .ck(ispd_clk), .d(n_18796), .o(x_out_35_22) );
ms00f80 x_out_35_reg_23_ ( .ck(ispd_clk), .d(n_19281), .o(x_out_35_23) );
ms00f80 x_out_35_reg_24_ ( .ck(ispd_clk), .d(n_20319), .o(x_out_35_24) );
ms00f80 x_out_35_reg_25_ ( .ck(ispd_clk), .d(n_21080), .o(x_out_35_25) );
ms00f80 x_out_35_reg_26_ ( .ck(ispd_clk), .d(n_21902), .o(x_out_35_26) );
ms00f80 x_out_35_reg_27_ ( .ck(ispd_clk), .d(n_23133), .o(x_out_35_27) );
ms00f80 x_out_35_reg_28_ ( .ck(ispd_clk), .d(n_23809), .o(x_out_35_28) );
ms00f80 x_out_35_reg_29_ ( .ck(ispd_clk), .d(n_24819), .o(x_out_35_29) );
ms00f80 x_out_35_reg_2_ ( .ck(ispd_clk), .d(n_21643), .o(x_out_35_2) );
ms00f80 x_out_35_reg_30_ ( .ck(ispd_clk), .d(n_25520), .o(x_out_35_30) );
ms00f80 x_out_35_reg_31_ ( .ck(ispd_clk), .d(n_26679), .o(x_out_35_31) );
ms00f80 x_out_35_reg_32_ ( .ck(ispd_clk), .d(n_27048), .o(x_out_35_32) );
ms00f80 x_out_35_reg_33_ ( .ck(ispd_clk), .d(n_27045), .o(x_out_35_33) );
ms00f80 x_out_35_reg_3_ ( .ck(ispd_clk), .d(n_22376), .o(x_out_35_3) );
ms00f80 x_out_35_reg_4_ ( .ck(ispd_clk), .d(n_23299), .o(x_out_35_4) );
ms00f80 x_out_35_reg_5_ ( .ck(ispd_clk), .d(n_24294), .o(x_out_35_5) );
ms00f80 x_out_35_reg_6_ ( .ck(ispd_clk), .d(n_25351), .o(x_out_35_6) );
ms00f80 x_out_35_reg_7_ ( .ck(ispd_clk), .d(n_26228), .o(x_out_35_7) );
ms00f80 x_out_35_reg_8_ ( .ck(ispd_clk), .d(n_27348), .o(x_out_35_8) );
ms00f80 x_out_35_reg_9_ ( .ck(ispd_clk), .d(n_28083), .o(x_out_35_9) );
ms00f80 x_out_36_reg_0_ ( .ck(ispd_clk), .d(n_11146), .o(x_out_36_0) );
ms00f80 x_out_36_reg_10_ ( .ck(ispd_clk), .d(n_27014), .o(x_out_36_10) );
ms00f80 x_out_36_reg_11_ ( .ck(ispd_clk), .d(n_27859), .o(x_out_36_11) );
ms00f80 x_out_36_reg_12_ ( .ck(ispd_clk), .d(n_28398), .o(x_out_36_12) );
ms00f80 x_out_36_reg_13_ ( .ck(ispd_clk), .d(n_28772), .o(x_out_36_13) );
ms00f80 x_out_36_reg_14_ ( .ck(ispd_clk), .d(n_29109), .o(x_out_36_14) );
ms00f80 x_out_36_reg_15_ ( .ck(ispd_clk), .d(n_29463), .o(x_out_36_15) );
ms00f80 x_out_36_reg_18_ ( .ck(ispd_clk), .d(n_11074), .o(x_out_36_18) );
ms00f80 x_out_36_reg_19_ ( .ck(ispd_clk), .d(n_16968), .o(x_out_36_19) );
ms00f80 x_out_36_reg_1_ ( .ck(ispd_clk), .d(n_16752), .o(x_out_36_1) );
ms00f80 x_out_36_reg_20_ ( .ck(ispd_clk), .d(n_17371), .o(x_out_36_20) );
ms00f80 x_out_36_reg_21_ ( .ck(ispd_clk), .d(n_17919), .o(x_out_36_21) );
ms00f80 x_out_36_reg_22_ ( .ck(ispd_clk), .d(n_18519), .o(x_out_36_22) );
ms00f80 x_out_36_reg_23_ ( .ck(ispd_clk), .d(n_19439), .o(x_out_36_23) );
ms00f80 x_out_36_reg_24_ ( .ck(ispd_clk), .d(n_20534), .o(x_out_36_24) );
ms00f80 x_out_36_reg_25_ ( .ck(ispd_clk), .d(n_21641), .o(x_out_36_25) );
ms00f80 x_out_36_reg_26_ ( .ck(ispd_clk), .d(n_22375), .o(x_out_36_26) );
ms00f80 x_out_36_reg_27_ ( .ck(ispd_clk), .d(n_23369), .o(x_out_36_27) );
ms00f80 x_out_36_reg_28_ ( .ck(ispd_clk), .d(n_24324), .o(x_out_36_28) );
ms00f80 x_out_36_reg_29_ ( .ck(ispd_clk), .d(n_25374), .o(x_out_36_29) );
ms00f80 x_out_36_reg_2_ ( .ck(ispd_clk), .d(n_18409), .o(x_out_36_2) );
ms00f80 x_out_36_reg_30_ ( .ck(ispd_clk), .d(n_25727), .o(x_out_36_30) );
ms00f80 x_out_36_reg_31_ ( .ck(ispd_clk), .d(n_26580), .o(x_out_36_31) );
ms00f80 x_out_36_reg_32_ ( .ck(ispd_clk), .d(n_26608), .o(x_out_36_32) );
ms00f80 x_out_36_reg_33_ ( .ck(ispd_clk), .d(n_26607), .o(x_out_36_33) );
ms00f80 x_out_36_reg_3_ ( .ck(ispd_clk), .d(n_19747), .o(x_out_36_3) );
ms00f80 x_out_36_reg_4_ ( .ck(ispd_clk), .d(n_20882), .o(x_out_36_4) );
ms00f80 x_out_36_reg_5_ ( .ck(ispd_clk), .d(n_21601), .o(x_out_36_5) );
ms00f80 x_out_36_reg_6_ ( .ck(ispd_clk), .d(n_22308), .o(x_out_36_6) );
ms00f80 x_out_36_reg_7_ ( .ck(ispd_clk), .d(n_23610), .o(x_out_36_7) );
ms00f80 x_out_36_reg_8_ ( .ck(ispd_clk), .d(n_24920), .o(x_out_36_8) );
ms00f80 x_out_36_reg_9_ ( .ck(ispd_clk), .d(n_26127), .o(x_out_36_9) );
ms00f80 x_out_37_reg_0_ ( .ck(ispd_clk), .d(n_16979), .o(x_out_37_0) );
ms00f80 x_out_37_reg_10_ ( .ck(ispd_clk), .d(n_28365), .o(x_out_37_10) );
ms00f80 x_out_37_reg_11_ ( .ck(ispd_clk), .d(n_28741), .o(x_out_37_11) );
ms00f80 x_out_37_reg_12_ ( .ck(ispd_clk), .d(n_29174), .o(x_out_37_12) );
ms00f80 x_out_37_reg_13_ ( .ck(ispd_clk), .d(n_29410), .o(x_out_37_13) );
ms00f80 x_out_37_reg_14_ ( .ck(ispd_clk), .d(n_29647), .o(x_out_37_14) );
ms00f80 x_out_37_reg_15_ ( .ck(ispd_clk), .d(n_29705), .o(x_out_37_15) );
ms00f80 x_out_37_reg_18_ ( .ck(ispd_clk), .d(n_7410), .o(x_out_37_18) );
ms00f80 x_out_37_reg_19_ ( .ck(ispd_clk), .d(n_10608), .o(x_out_37_19) );
ms00f80 x_out_37_reg_1_ ( .ck(ispd_clk), .d(n_20180), .o(x_out_37_1) );
ms00f80 x_out_37_reg_20_ ( .ck(ispd_clk), .d(n_11674), .o(x_out_37_20) );
ms00f80 x_out_37_reg_21_ ( .ck(ispd_clk), .d(n_14129), .o(x_out_37_21) );
ms00f80 x_out_37_reg_22_ ( .ck(ispd_clk), .d(n_15664), .o(x_out_37_22) );
ms00f80 x_out_37_reg_23_ ( .ck(ispd_clk), .d(n_16291), .o(x_out_37_23) );
ms00f80 x_out_37_reg_24_ ( .ck(ispd_clk), .d(n_16875), .o(x_out_37_24) );
ms00f80 x_out_37_reg_25_ ( .ck(ispd_clk), .d(n_18041), .o(x_out_37_25) );
ms00f80 x_out_37_reg_26_ ( .ck(ispd_clk), .d(n_19366), .o(x_out_37_26) );
ms00f80 x_out_37_reg_27_ ( .ck(ispd_clk), .d(n_20352), .o(x_out_37_27) );
ms00f80 x_out_37_reg_28_ ( .ck(ispd_clk), .d(n_21452), .o(x_out_37_28) );
ms00f80 x_out_37_reg_29_ ( .ck(ispd_clk), .d(n_22751), .o(x_out_37_29) );
ms00f80 x_out_37_reg_2_ ( .ck(ispd_clk), .d(n_21264), .o(x_out_37_2) );
ms00f80 x_out_37_reg_30_ ( .ck(ispd_clk), .d(n_23714), .o(x_out_37_30) );
ms00f80 x_out_37_reg_31_ ( .ck(ispd_clk), .d(n_24711), .o(x_out_37_31) );
ms00f80 x_out_37_reg_32_ ( .ck(ispd_clk), .d(n_25099), .o(x_out_37_32) );
ms00f80 x_out_37_reg_33_ ( .ck(ispd_clk), .d(n_24850), .o(x_out_37_33) );
ms00f80 x_out_37_reg_3_ ( .ck(ispd_clk), .d(n_22056), .o(x_out_37_3) );
ms00f80 x_out_37_reg_4_ ( .ck(ispd_clk), .d(n_23048), .o(x_out_37_4) );
ms00f80 x_out_37_reg_5_ ( .ck(ispd_clk), .d(n_24293), .o(x_out_37_5) );
ms00f80 x_out_37_reg_6_ ( .ck(ispd_clk), .d(n_25024), .o(x_out_37_6) );
ms00f80 x_out_37_reg_7_ ( .ck(ispd_clk), .d(n_25971), .o(x_out_37_7) );
ms00f80 x_out_37_reg_8_ ( .ck(ispd_clk), .d(n_27150), .o(x_out_37_8) );
ms00f80 x_out_37_reg_9_ ( .ck(ispd_clk), .d(n_27928), .o(x_out_37_9) );
ms00f80 x_out_38_reg_0_ ( .ck(ispd_clk), .d(n_14286), .o(x_out_38_0) );
ms00f80 x_out_38_reg_10_ ( .ck(ispd_clk), .d(n_26843), .o(x_out_38_10) );
ms00f80 x_out_38_reg_11_ ( .ck(ispd_clk), .d(n_27747), .o(x_out_38_11) );
ms00f80 x_out_38_reg_12_ ( .ck(ispd_clk), .d(n_28235), .o(x_out_38_12) );
ms00f80 x_out_38_reg_13_ ( .ck(ispd_clk), .d(n_28712), .o(x_out_38_13) );
ms00f80 x_out_38_reg_14_ ( .ck(ispd_clk), .d(n_29069), .o(x_out_38_14) );
ms00f80 x_out_38_reg_15_ ( .ck(ispd_clk), .d(n_29300), .o(x_out_38_15) );
ms00f80 x_out_38_reg_18_ ( .ck(ispd_clk), .d(n_17221), .o(x_out_38_18) );
ms00f80 x_out_38_reg_19_ ( .ck(ispd_clk), .d(n_17936), .o(x_out_38_19) );
ms00f80 x_out_38_reg_1_ ( .ck(ispd_clk), .d(n_17370), .o(x_out_38_1) );
ms00f80 x_out_38_reg_20_ ( .ck(ispd_clk), .d(n_20224), .o(x_out_38_20) );
ms00f80 x_out_38_reg_21_ ( .ck(ispd_clk), .d(n_21323), .o(x_out_38_21) );
ms00f80 x_out_38_reg_22_ ( .ck(ispd_clk), .d(n_21809), .o(x_out_38_22) );
ms00f80 x_out_38_reg_23_ ( .ck(ispd_clk), .d(n_23077), .o(x_out_38_23) );
ms00f80 x_out_38_reg_24_ ( .ck(ispd_clk), .d(n_23713), .o(x_out_38_24) );
ms00f80 x_out_38_reg_25_ ( .ck(ispd_clk), .d(n_25035), .o(x_out_38_25) );
ms00f80 x_out_38_reg_26_ ( .ck(ispd_clk), .d(n_25422), .o(x_out_38_26) );
ms00f80 x_out_38_reg_27_ ( .ck(ispd_clk), .d(n_26620), .o(x_out_38_27) );
ms00f80 x_out_38_reg_28_ ( .ck(ispd_clk), .d(n_27029), .o(x_out_38_28) );
ms00f80 x_out_38_reg_29_ ( .ck(ispd_clk), .d(n_27913), .o(x_out_38_29) );
ms00f80 x_out_38_reg_2_ ( .ck(ispd_clk), .d(n_18280), .o(x_out_38_2) );
ms00f80 x_out_38_reg_30_ ( .ck(ispd_clk), .d(n_28124), .o(x_out_38_30) );
ms00f80 x_out_38_reg_31_ ( .ck(ispd_clk), .d(n_28635), .o(x_out_38_31) );
ms00f80 x_out_38_reg_32_ ( .ck(ispd_clk), .d(n_28708), .o(x_out_38_32) );
ms00f80 x_out_38_reg_33_ ( .ck(ispd_clk), .d(n_28716), .o(x_out_38_33) );
ms00f80 x_out_38_reg_3_ ( .ck(ispd_clk), .d(n_19438), .o(x_out_38_3) );
ms00f80 x_out_38_reg_4_ ( .ck(ispd_clk), .d(n_20533), .o(x_out_38_4) );
ms00f80 x_out_38_reg_5_ ( .ck(ispd_clk), .d(n_21322), .o(x_out_38_5) );
ms00f80 x_out_38_reg_6_ ( .ck(ispd_clk), .d(n_22105), .o(x_out_38_6) );
ms00f80 x_out_38_reg_7_ ( .ck(ispd_clk), .d(n_23367), .o(x_out_38_7) );
ms00f80 x_out_38_reg_8_ ( .ck(ispd_clk), .d(n_24665), .o(x_out_38_8) );
ms00f80 x_out_38_reg_9_ ( .ck(ispd_clk), .d(n_25933), .o(x_out_38_9) );
ms00f80 x_out_39_reg_0_ ( .ck(ispd_clk), .d(n_13925), .o(x_out_39_0) );
ms00f80 x_out_39_reg_10_ ( .ck(ispd_clk), .d(n_27690), .o(x_out_39_10) );
ms00f80 x_out_39_reg_11_ ( .ck(ispd_clk), .d(n_28301), .o(x_out_39_11) );
ms00f80 x_out_39_reg_12_ ( .ck(ispd_clk), .d(n_28673), .o(x_out_39_12) );
ms00f80 x_out_39_reg_13_ ( .ck(ispd_clk), .d(n_29027), .o(x_out_39_13) );
ms00f80 x_out_39_reg_14_ ( .ck(ispd_clk), .d(n_29401), .o(x_out_39_14) );
ms00f80 x_out_39_reg_15_ ( .ck(ispd_clk), .d(n_29592), .o(x_out_39_15) );
ms00f80 x_out_39_reg_18_ ( .ck(ispd_clk), .d(n_14627), .o(x_out_39_18) );
ms00f80 x_out_39_reg_19_ ( .ck(ispd_clk), .d(n_17219), .o(x_out_39_19) );
ms00f80 x_out_39_reg_1_ ( .ck(ispd_clk), .d(n_17917), .o(x_out_39_1) );
ms00f80 x_out_39_reg_20_ ( .ck(ispd_clk), .d(n_17368), .o(x_out_39_20) );
ms00f80 x_out_39_reg_21_ ( .ck(ispd_clk), .d(n_18279), .o(x_out_39_21) );
ms00f80 x_out_39_reg_22_ ( .ck(ispd_clk), .d(n_18986), .o(x_out_39_22) );
ms00f80 x_out_39_reg_23_ ( .ck(ispd_clk), .d(n_20318), .o(x_out_39_23) );
ms00f80 x_out_39_reg_24_ ( .ck(ispd_clk), .d(n_20800), .o(x_out_39_24) );
ms00f80 x_out_39_reg_25_ ( .ck(ispd_clk), .d(n_22158), .o(x_out_39_25) );
ms00f80 x_out_39_reg_26_ ( .ck(ispd_clk), .d(n_22849), .o(x_out_39_26) );
ms00f80 x_out_39_reg_27_ ( .ck(ispd_clk), .d(n_24089), .o(x_out_39_27) );
ms00f80 x_out_39_reg_28_ ( .ck(ispd_clk), .d(n_24492), .o(x_out_39_28) );
ms00f80 x_out_39_reg_29_ ( .ck(ispd_clk), .d(n_25796), .o(x_out_39_29) );
ms00f80 x_out_39_reg_2_ ( .ck(ispd_clk), .d(n_19437), .o(x_out_39_2) );
ms00f80 x_out_39_reg_30_ ( .ck(ispd_clk), .d(n_26437), .o(x_out_39_30) );
ms00f80 x_out_39_reg_31_ ( .ck(ispd_clk), .d(n_27346), .o(x_out_39_31) );
ms00f80 x_out_39_reg_32_ ( .ck(ispd_clk), .d(n_27788), .o(x_out_39_32) );
ms00f80 x_out_39_reg_33_ ( .ck(ispd_clk), .d(n_27687), .o(x_out_39_33) );
ms00f80 x_out_39_reg_3_ ( .ck(ispd_clk), .d(n_20179), .o(x_out_39_3) );
ms00f80 x_out_39_reg_4_ ( .ck(ispd_clk), .d(n_20961), .o(x_out_39_4) );
ms00f80 x_out_39_reg_5_ ( .ck(ispd_clk), .d(n_22055), .o(x_out_39_5) );
ms00f80 x_out_39_reg_6_ ( .ck(ispd_clk), .d(n_23297), .o(x_out_39_6) );
ms00f80 x_out_39_reg_7_ ( .ck(ispd_clk), .d(n_24601), .o(x_out_39_7) );
ms00f80 x_out_39_reg_8_ ( .ck(ispd_clk), .d(n_25884), .o(x_out_39_8) );
ms00f80 x_out_39_reg_9_ ( .ck(ispd_clk), .d(n_26771), .o(x_out_39_9) );
ms00f80 x_out_3_reg_0_ ( .ck(ispd_clk), .d(n_16974), .o(x_out_3_0) );
ms00f80 x_out_3_reg_10_ ( .ck(ispd_clk), .d(n_28298), .o(x_out_3_10) );
ms00f80 x_out_3_reg_11_ ( .ck(ispd_clk), .d(n_28672), .o(x_out_3_11) );
ms00f80 x_out_3_reg_12_ ( .ck(ispd_clk), .d(n_29024), .o(x_out_3_12) );
ms00f80 x_out_3_reg_13_ ( .ck(ispd_clk), .d(n_29399), .o(x_out_3_13) );
ms00f80 x_out_3_reg_14_ ( .ck(ispd_clk), .d(n_29524), .o(x_out_3_14) );
ms00f80 x_out_3_reg_15_ ( .ck(ispd_clk), .d(n_29656), .o(x_out_3_15) );
ms00f80 x_out_3_reg_18_ ( .ck(ispd_clk), .d(n_10661), .o(x_out_3_18) );
ms00f80 x_out_3_reg_19_ ( .ck(ispd_clk), .d(n_16076), .o(x_out_3_19) );
ms00f80 x_out_3_reg_1_ ( .ck(ispd_clk), .d(n_18278), .o(x_out_3_1) );
ms00f80 x_out_3_reg_20_ ( .ck(ispd_clk), .d(n_14665), .o(x_out_3_20) );
ms00f80 x_out_3_reg_21_ ( .ck(ispd_clk), .d(n_15931), .o(x_out_3_21) );
ms00f80 x_out_3_reg_22_ ( .ck(ispd_clk), .d(n_17078), .o(x_out_3_22) );
ms00f80 x_out_3_reg_23_ ( .ck(ispd_clk), .d(n_17774), .o(x_out_3_23) );
ms00f80 x_out_3_reg_24_ ( .ck(ispd_clk), .d(n_18985), .o(x_out_3_24) );
ms00f80 x_out_3_reg_25_ ( .ck(ispd_clk), .d(n_19651), .o(x_out_3_25) );
ms00f80 x_out_3_reg_26_ ( .ck(ispd_clk), .d(n_20799), .o(x_out_3_26) );
ms00f80 x_out_3_reg_27_ ( .ck(ispd_clk), .d(n_21538), .o(x_out_3_27) );
ms00f80 x_out_3_reg_28_ ( .ck(ispd_clk), .d(n_22848), .o(x_out_3_28) );
ms00f80 x_out_3_reg_29_ ( .ck(ispd_clk), .d(n_23545), .o(x_out_3_29) );
ms00f80 x_out_3_reg_2_ ( .ck(ispd_clk), .d(n_20223), .o(x_out_3_2) );
ms00f80 x_out_3_reg_30_ ( .ck(ispd_clk), .d(n_24491), .o(x_out_3_30) );
ms00f80 x_out_3_reg_31_ ( .ck(ispd_clk), .d(n_25233), .o(x_out_3_31) );
ms00f80 x_out_3_reg_32_ ( .ck(ispd_clk), .d(n_27074), .o(x_out_3_32) );
ms00f80 x_out_3_reg_33_ ( .ck(ispd_clk), .d(n_27072), .o(x_out_3_33) );
ms00f80 x_out_3_reg_3_ ( .ck(ispd_clk), .d(n_21640), .o(x_out_3_3) );
ms00f80 x_out_3_reg_4_ ( .ck(ispd_clk), .d(n_22053), .o(x_out_3_4) );
ms00f80 x_out_3_reg_5_ ( .ck(ispd_clk), .d(n_23295), .o(x_out_3_5) );
ms00f80 x_out_3_reg_6_ ( .ck(ispd_clk), .d(n_24598), .o(x_out_3_6) );
ms00f80 x_out_3_reg_7_ ( .ck(ispd_clk), .d(n_25881), .o(x_out_3_7) );
ms00f80 x_out_3_reg_8_ ( .ck(ispd_clk), .d(n_26766), .o(x_out_3_8) );
ms00f80 x_out_3_reg_9_ ( .ck(ispd_clk), .d(n_27685), .o(x_out_3_9) );
ms00f80 x_out_40_reg_0_ ( .ck(ispd_clk), .d(n_6071), .o(x_out_40_0) );
ms00f80 x_out_40_reg_10_ ( .ck(ispd_clk), .d(n_22371), .o(x_out_40_10) );
ms00f80 x_out_40_reg_11_ ( .ck(ispd_clk), .d(n_23652), .o(x_out_40_11) );
ms00f80 x_out_40_reg_12_ ( .ck(ispd_clk), .d(n_24663), .o(x_out_40_12) );
ms00f80 x_out_40_reg_13_ ( .ck(ispd_clk), .d(n_25969), .o(x_out_40_13) );
ms00f80 x_out_40_reg_14_ ( .ck(ispd_clk), .d(n_25970), .o(x_out_40_14) );
ms00f80 x_out_40_reg_15_ ( .ck(ispd_clk), .d(n_26924), .o(x_out_40_15) );
ms00f80 x_out_40_reg_18_ ( .ck(ispd_clk), .d(n_14626), .o(x_out_40_18) );
ms00f80 x_out_40_reg_19_ ( .ck(ispd_clk), .d(n_16566), .o(x_out_40_19) );
ms00f80 x_out_40_reg_1_ ( .ck(ispd_clk), .d(n_11022), .o(x_out_40_1) );
ms00f80 x_out_40_reg_20_ ( .ck(ispd_clk), .d(n_17077), .o(x_out_40_20) );
ms00f80 x_out_40_reg_21_ ( .ck(ispd_clk), .d(n_18010), .o(x_out_40_21) );
ms00f80 x_out_40_reg_22_ ( .ck(ispd_clk), .d(n_18984), .o(x_out_40_22) );
ms00f80 x_out_40_reg_23_ ( .ck(ispd_clk), .d(n_19991), .o(x_out_40_23) );
ms00f80 x_out_40_reg_24_ ( .ck(ispd_clk), .d(n_20798), .o(x_out_40_24) );
ms00f80 x_out_40_reg_25_ ( .ck(ispd_clk), .d(n_21899), .o(x_out_40_25) );
ms00f80 x_out_40_reg_26_ ( .ck(ispd_clk), .d(n_22847), .o(x_out_40_26) );
ms00f80 x_out_40_reg_27_ ( .ck(ispd_clk), .d(n_23807), .o(x_out_40_27) );
ms00f80 x_out_40_reg_28_ ( .ck(ispd_clk), .d(n_24490), .o(x_out_40_28) );
ms00f80 x_out_40_reg_29_ ( .ck(ispd_clk), .d(n_25518), .o(x_out_40_29) );
ms00f80 x_out_40_reg_2_ ( .ck(ispd_clk), .d(n_12570), .o(x_out_40_2) );
ms00f80 x_out_40_reg_30_ ( .ck(ispd_clk), .d(n_26436), .o(x_out_40_30) );
ms00f80 x_out_40_reg_31_ ( .ck(ispd_clk), .d(n_27148), .o(x_out_40_31) );
ms00f80 x_out_40_reg_32_ ( .ck(ispd_clk), .d(n_27611), .o(x_out_40_32) );
ms00f80 x_out_40_reg_33_ ( .ck(ispd_clk), .d(n_27485), .o(x_out_40_33) );
ms00f80 x_out_40_reg_3_ ( .ck(ispd_clk), .d(n_13768), .o(x_out_40_3) );
ms00f80 x_out_40_reg_4_ ( .ck(ispd_clk), .d(n_14993), .o(x_out_40_4) );
ms00f80 x_out_40_reg_5_ ( .ck(ispd_clk), .d(n_16290), .o(x_out_40_5) );
ms00f80 x_out_40_reg_6_ ( .ck(ispd_clk), .d(n_17420), .o(x_out_40_6) );
ms00f80 x_out_40_reg_7_ ( .ck(ispd_clk), .d(n_18573), .o(x_out_40_7) );
ms00f80 x_out_40_reg_8_ ( .ck(ispd_clk), .d(n_19889), .o(x_out_40_8) );
ms00f80 x_out_40_reg_9_ ( .ck(ispd_clk), .d(n_21321), .o(x_out_40_9) );
ms00f80 x_out_41_reg_0_ ( .ck(ispd_clk), .d(n_16972), .o(x_out_41_0) );
ms00f80 x_out_41_reg_10_ ( .ck(ispd_clk), .d(n_28598), .o(x_out_41_10) );
ms00f80 x_out_41_reg_11_ ( .ck(ispd_clk), .d(n_28910), .o(x_out_41_11) );
ms00f80 x_out_41_reg_12_ ( .ck(ispd_clk), .d(n_29302), .o(x_out_41_12) );
ms00f80 x_out_41_reg_13_ ( .ck(ispd_clk), .d(n_29629), .o(x_out_41_13) );
ms00f80 x_out_41_reg_14_ ( .ck(ispd_clk), .d(n_29688), .o(x_out_41_14) );
ms00f80 x_out_41_reg_15_ ( .ck(ispd_clk), .d(n_29709), .o(x_out_41_15) );
ms00f80 x_out_41_reg_18_ ( .ck(ispd_clk), .d(n_14623), .o(x_out_41_18) );
ms00f80 x_out_41_reg_19_ ( .ck(ispd_clk), .d(n_16570), .o(x_out_41_19) );
ms00f80 x_out_41_reg_1_ ( .ck(ispd_clk), .d(n_21572), .o(x_out_41_1) );
ms00f80 x_out_41_reg_20_ ( .ck(ispd_clk), .d(n_17365), .o(x_out_41_20) );
ms00f80 x_out_41_reg_21_ ( .ck(ispd_clk), .d(n_18277), .o(x_out_41_21) );
ms00f80 x_out_41_reg_22_ ( .ck(ispd_clk), .d(n_19277), .o(x_out_41_22) );
ms00f80 x_out_41_reg_23_ ( .ck(ispd_clk), .d(n_20317), .o(x_out_41_23) );
ms00f80 x_out_41_reg_24_ ( .ck(ispd_clk), .d(n_21075), .o(x_out_41_24) );
ms00f80 x_out_41_reg_25_ ( .ck(ispd_clk), .d(n_22157), .o(x_out_41_25) );
ms00f80 x_out_41_reg_26_ ( .ck(ispd_clk), .d(n_23129), .o(x_out_41_26) );
ms00f80 x_out_41_reg_27_ ( .ck(ispd_clk), .d(n_24088), .o(x_out_41_27) );
ms00f80 x_out_41_reg_28_ ( .ck(ispd_clk), .d(n_24816), .o(x_out_41_28) );
ms00f80 x_out_41_reg_29_ ( .ck(ispd_clk), .d(n_25795), .o(x_out_41_29) );
ms00f80 x_out_41_reg_2_ ( .ck(ispd_clk), .d(n_22276), .o(x_out_41_2) );
ms00f80 x_out_41_reg_30_ ( .ck(ispd_clk), .d(n_26675), .o(x_out_41_30) );
ms00f80 x_out_41_reg_31_ ( .ck(ispd_clk), .d(n_27344), .o(x_out_41_31) );
ms00f80 x_out_41_reg_32_ ( .ck(ispd_clk), .d(n_27615), .o(x_out_41_32) );
ms00f80 x_out_41_reg_33_ ( .ck(ispd_clk), .d(n_27610), .o(x_out_41_33) );
ms00f80 x_out_41_reg_3_ ( .ck(ispd_clk), .d(n_22949), .o(x_out_41_3) );
ms00f80 x_out_41_reg_4_ ( .ck(ispd_clk), .d(n_23920), .o(x_out_41_4) );
ms00f80 x_out_41_reg_5_ ( .ck(ispd_clk), .d(n_24919), .o(x_out_41_5) );
ms00f80 x_out_41_reg_6_ ( .ck(ispd_clk), .d(n_26122), .o(x_out_41_6) );
ms00f80 x_out_41_reg_7_ ( .ck(ispd_clk), .d(n_27243), .o(x_out_41_7) );
ms00f80 x_out_41_reg_8_ ( .ck(ispd_clk), .d(n_27682), .o(x_out_41_8) );
ms00f80 x_out_41_reg_9_ ( .ck(ispd_clk), .d(n_28207), .o(x_out_41_9) );
ms00f80 x_out_42_reg_0_ ( .ck(ispd_clk), .d(n_17237), .o(x_out_42_0) );
ms00f80 x_out_42_reg_10_ ( .ck(ispd_clk), .d(n_28769), .o(x_out_42_10) );
ms00f80 x_out_42_reg_11_ ( .ck(ispd_clk), .d(n_29105), .o(x_out_42_11) );
ms00f80 x_out_42_reg_12_ ( .ck(ispd_clk), .d(n_29462), .o(x_out_42_12) );
ms00f80 x_out_42_reg_13_ ( .ck(ispd_clk), .d(n_29638), .o(x_out_42_13) );
ms00f80 x_out_42_reg_14_ ( .ck(ispd_clk), .d(n_29708), .o(x_out_42_14) );
ms00f80 x_out_42_reg_15_ ( .ck(ispd_clk), .d(n_29710), .o(x_out_42_15) );
ms00f80 x_out_42_reg_18_ ( .ck(ispd_clk), .d(n_14622), .o(x_out_42_18) );
ms00f80 x_out_42_reg_19_ ( .ck(ispd_clk), .d(n_16569), .o(x_out_42_19) );
ms00f80 x_out_42_reg_1_ ( .ck(ispd_clk), .d(n_21197), .o(x_out_42_1) );
ms00f80 x_out_42_reg_20_ ( .ck(ispd_clk), .d(n_17364), .o(x_out_42_20) );
ms00f80 x_out_42_reg_21_ ( .ck(ispd_clk), .d(n_18276), .o(x_out_42_21) );
ms00f80 x_out_42_reg_22_ ( .ck(ispd_clk), .d(n_19276), .o(x_out_42_22) );
ms00f80 x_out_42_reg_23_ ( .ck(ispd_clk), .d(n_20316), .o(x_out_42_23) );
ms00f80 x_out_42_reg_24_ ( .ck(ispd_clk), .d(n_21074), .o(x_out_42_24) );
ms00f80 x_out_42_reg_25_ ( .ck(ispd_clk), .d(n_22156), .o(x_out_42_25) );
ms00f80 x_out_42_reg_26_ ( .ck(ispd_clk), .d(n_23128), .o(x_out_42_26) );
ms00f80 x_out_42_reg_27_ ( .ck(ispd_clk), .d(n_24087), .o(x_out_42_27) );
ms00f80 x_out_42_reg_28_ ( .ck(ispd_clk), .d(n_25091), .o(x_out_42_28) );
ms00f80 x_out_42_reg_29_ ( .ck(ispd_clk), .d(n_25794), .o(x_out_42_29) );
ms00f80 x_out_42_reg_2_ ( .ck(ispd_clk), .d(n_22589), .o(x_out_42_2) );
ms00f80 x_out_42_reg_30_ ( .ck(ispd_clk), .d(n_26672), .o(x_out_42_30) );
ms00f80 x_out_42_reg_31_ ( .ck(ispd_clk), .d(n_27343), .o(x_out_42_31) );
ms00f80 x_out_42_reg_32_ ( .ck(ispd_clk), .d(n_27860), .o(x_out_42_32) );
ms00f80 x_out_42_reg_33_ ( .ck(ispd_clk), .d(n_28019), .o(x_out_42_33) );
ms00f80 x_out_42_reg_3_ ( .ck(ispd_clk), .d(n_23246), .o(x_out_42_3) );
ms00f80 x_out_42_reg_4_ ( .ck(ispd_clk), .d(n_23609), .o(x_out_42_4) );
ms00f80 x_out_42_reg_5_ ( .ck(ispd_clk), .d(n_24918), .o(x_out_42_5) );
ms00f80 x_out_42_reg_6_ ( .ck(ispd_clk), .d(n_26121), .o(x_out_42_6) );
ms00f80 x_out_42_reg_7_ ( .ck(ispd_clk), .d(n_27242), .o(x_out_42_7) );
ms00f80 x_out_42_reg_8_ ( .ck(ispd_clk), .d(n_27858), .o(x_out_42_8) );
ms00f80 x_out_42_reg_9_ ( .ck(ispd_clk), .d(n_28396), .o(x_out_42_9) );
ms00f80 x_out_43_reg_0_ ( .ck(ispd_clk), .d(n_16780), .o(x_out_43_0) );
ms00f80 x_out_43_reg_10_ ( .ck(ispd_clk), .d(n_28107), .o(x_out_43_10) );
ms00f80 x_out_43_reg_11_ ( .ck(ispd_clk), .d(n_28527), .o(x_out_43_11) );
ms00f80 x_out_43_reg_12_ ( .ck(ispd_clk), .d(n_28981), .o(x_out_43_12) );
ms00f80 x_out_43_reg_13_ ( .ck(ispd_clk), .d(n_29256), .o(x_out_43_13) );
ms00f80 x_out_43_reg_14_ ( .ck(ispd_clk), .d(n_29497), .o(x_out_43_14) );
ms00f80 x_out_43_reg_15_ ( .ck(ispd_clk), .d(n_29685), .o(x_out_43_15) );
ms00f80 x_out_43_reg_18_ ( .ck(ispd_clk), .d(n_17218), .o(x_out_43_18) );
ms00f80 x_out_43_reg_19_ ( .ck(ispd_clk), .d(n_17935), .o(x_out_43_19) );
ms00f80 x_out_43_reg_1_ ( .ck(ispd_clk), .d(n_19826), .o(x_out_43_1) );
ms00f80 x_out_43_reg_20_ ( .ck(ispd_clk), .d(n_19275), .o(x_out_43_20) );
ms00f80 x_out_43_reg_21_ ( .ck(ispd_clk), .d(n_20315), .o(x_out_43_21) );
ms00f80 x_out_43_reg_22_ ( .ck(ispd_clk), .d(n_20797), .o(x_out_43_22) );
ms00f80 x_out_43_reg_23_ ( .ck(ispd_clk), .d(n_22155), .o(x_out_43_23) );
ms00f80 x_out_43_reg_24_ ( .ck(ispd_clk), .d(n_22846), .o(x_out_43_24) );
ms00f80 x_out_43_reg_25_ ( .ck(ispd_clk), .d(n_24086), .o(x_out_43_25) );
ms00f80 x_out_43_reg_26_ ( .ck(ispd_clk), .d(n_24815), .o(x_out_43_26) );
ms00f80 x_out_43_reg_27_ ( .ck(ispd_clk), .d(n_25793), .o(x_out_43_27) );
ms00f80 x_out_43_reg_28_ ( .ck(ispd_clk), .d(n_26434), .o(x_out_43_28) );
ms00f80 x_out_43_reg_29_ ( .ck(ispd_clk), .d(n_27341), .o(x_out_43_29) );
ms00f80 x_out_43_reg_2_ ( .ck(ispd_clk), .d(n_21263), .o(x_out_43_2) );
ms00f80 x_out_43_reg_30_ ( .ck(ispd_clk), .d(n_27647), .o(x_out_43_30) );
ms00f80 x_out_43_reg_31_ ( .ck(ispd_clk), .d(n_28324), .o(x_out_43_31) );
ms00f80 x_out_43_reg_32_ ( .ck(ispd_clk), .d(n_28511), .o(x_out_43_32) );
ms00f80 x_out_43_reg_33_ ( .ck(ispd_clk), .d(n_28645), .o(x_out_43_33) );
ms00f80 x_out_43_reg_3_ ( .ck(ispd_clk), .d(n_22307), .o(x_out_43_3) );
ms00f80 x_out_43_reg_4_ ( .ck(ispd_clk), .d(n_23292), .o(x_out_43_4) );
ms00f80 x_out_43_reg_5_ ( .ck(ispd_clk), .d(n_24291), .o(x_out_43_5) );
ms00f80 x_out_43_reg_6_ ( .ck(ispd_clk), .d(n_25022), .o(x_out_43_6) );
ms00f80 x_out_43_reg_7_ ( .ck(ispd_clk), .d(n_26220), .o(x_out_43_7) );
ms00f80 x_out_43_reg_8_ ( .ck(ispd_clk), .d(n_26923), .o(x_out_43_8) );
ms00f80 x_out_43_reg_9_ ( .ck(ispd_clk), .d(n_27614), .o(x_out_43_9) );
ms00f80 x_out_44_reg_0_ ( .ck(ispd_clk), .d(n_14225), .o(x_out_44_0) );
ms00f80 x_out_44_reg_10_ ( .ck(ispd_clk), .d(n_27927), .o(x_out_44_10) );
ms00f80 x_out_44_reg_11_ ( .ck(ispd_clk), .d(n_28359), .o(x_out_44_11) );
ms00f80 x_out_44_reg_12_ ( .ck(ispd_clk), .d(n_28736), .o(x_out_44_12) );
ms00f80 x_out_44_reg_13_ ( .ck(ispd_clk), .d(n_29167), .o(x_out_44_13) );
ms00f80 x_out_44_reg_14_ ( .ck(ispd_clk), .d(n_29437), .o(x_out_44_14) );
ms00f80 x_out_44_reg_15_ ( .ck(ispd_clk), .d(n_29646), .o(x_out_44_15) );
ms00f80 x_out_44_reg_18_ ( .ck(ispd_clk), .d(n_7226), .o(x_out_44_18) );
ms00f80 x_out_44_reg_19_ ( .ck(ispd_clk), .d(n_9802), .o(x_out_44_19) );
ms00f80 x_out_44_reg_1_ ( .ck(ispd_clk), .d(n_19150), .o(x_out_44_1) );
ms00f80 x_out_44_reg_20_ ( .ck(ispd_clk), .d(n_12869), .o(x_out_44_20) );
ms00f80 x_out_44_reg_21_ ( .ck(ispd_clk), .d(n_13767), .o(x_out_44_21) );
ms00f80 x_out_44_reg_22_ ( .ck(ispd_clk), .d(n_14520), .o(x_out_44_22) );
ms00f80 x_out_44_reg_23_ ( .ck(ispd_clk), .d(n_15276), .o(x_out_44_23) );
ms00f80 x_out_44_reg_24_ ( .ck(ispd_clk), .d(n_15977), .o(x_out_44_24) );
ms00f80 x_out_44_reg_25_ ( .ck(ispd_clk), .d(n_16874), .o(x_out_44_25) );
ms00f80 x_out_44_reg_26_ ( .ck(ispd_clk), .d(n_17797), .o(x_out_44_26) );
ms00f80 x_out_44_reg_27_ ( .ck(ispd_clk), .d(n_18673), .o(x_out_44_27) );
ms00f80 x_out_44_reg_28_ ( .ck(ispd_clk), .d(n_19675), .o(x_out_44_28) );
ms00f80 x_out_44_reg_29_ ( .ck(ispd_clk), .d(n_20463), .o(x_out_44_29) );
ms00f80 x_out_44_reg_2_ ( .ck(ispd_clk), .d(n_20493), .o(x_out_44_2) );
ms00f80 x_out_44_reg_30_ ( .ck(ispd_clk), .d(n_21561), .o(x_out_44_30) );
ms00f80 x_out_44_reg_31_ ( .ck(ispd_clk), .d(n_22576), .o(x_out_44_31) );
ms00f80 x_out_44_reg_32_ ( .ck(ispd_clk), .d(n_23228), .o(x_out_44_32) );
ms00f80 x_out_44_reg_33_ ( .ck(ispd_clk), .d(n_23571), .o(x_out_44_33) );
ms00f80 x_out_44_reg_3_ ( .ck(ispd_clk), .d(n_21987), .o(x_out_44_3) );
ms00f80 x_out_44_reg_4_ ( .ck(ispd_clk), .d(n_22609), .o(x_out_44_4) );
ms00f80 x_out_44_reg_5_ ( .ck(ispd_clk), .d(n_23289), .o(x_out_44_5) );
ms00f80 x_out_44_reg_6_ ( .ck(ispd_clk), .d(n_24290), .o(x_out_44_6) );
ms00f80 x_out_44_reg_7_ ( .ck(ispd_clk), .d(n_25656), .o(x_out_44_7) );
ms00f80 x_out_44_reg_8_ ( .ck(ispd_clk), .d(n_26516), .o(x_out_44_8) );
ms00f80 x_out_44_reg_9_ ( .ck(ispd_clk), .d(n_27147), .o(x_out_44_9) );
ms00f80 x_out_45_reg_0_ ( .ck(ispd_clk), .d(n_14639), .o(x_out_45_0) );
ms00f80 x_out_45_reg_10_ ( .ck(ispd_clk), .d(n_28011), .o(x_out_45_10) );
ms00f80 x_out_45_reg_11_ ( .ck(ispd_clk), .d(n_28424), .o(x_out_45_11) );
ms00f80 x_out_45_reg_12_ ( .ck(ispd_clk), .d(n_28867), .o(x_out_45_12) );
ms00f80 x_out_45_reg_13_ ( .ck(ispd_clk), .d(n_29206), .o(x_out_45_13) );
ms00f80 x_out_45_reg_14_ ( .ck(ispd_clk), .d(n_29493), .o(x_out_45_14) );
ms00f80 x_out_45_reg_15_ ( .ck(ispd_clk), .d(n_29657), .o(x_out_45_15) );
ms00f80 x_out_45_reg_18_ ( .ck(ispd_clk), .d(n_11771), .o(x_out_45_18) );
ms00f80 x_out_45_reg_19_ ( .ck(ispd_clk), .d(n_16751), .o(x_out_45_19) );
ms00f80 x_out_45_reg_1_ ( .ck(ispd_clk), .d(n_19149), .o(x_out_45_1) );
ms00f80 x_out_45_reg_20_ ( .ck(ispd_clk), .d(n_17601), .o(x_out_45_20) );
ms00f80 x_out_45_reg_21_ ( .ck(ispd_clk), .d(n_18275), .o(x_out_45_21) );
ms00f80 x_out_45_reg_22_ ( .ck(ispd_clk), .d(n_19436), .o(x_out_45_22) );
ms00f80 x_out_45_reg_23_ ( .ck(ispd_clk), .d(n_20532), .o(x_out_45_23) );
ms00f80 x_out_45_reg_24_ ( .ck(ispd_clk), .d(n_21599), .o(x_out_45_24) );
ms00f80 x_out_45_reg_25_ ( .ck(ispd_clk), .d(n_22050), .o(x_out_45_25) );
ms00f80 x_out_45_reg_26_ ( .ck(ispd_clk), .d(n_22958), .o(x_out_45_26) );
ms00f80 x_out_45_reg_27_ ( .ck(ispd_clk), .d(n_23937), .o(x_out_45_27) );
ms00f80 x_out_45_reg_28_ ( .ck(ispd_clk), .d(n_24983), .o(x_out_45_28) );
ms00f80 x_out_45_reg_29_ ( .ck(ispd_clk), .d(n_25878), .o(x_out_45_29) );
ms00f80 x_out_45_reg_2_ ( .ck(ispd_clk), .d(n_20177), .o(x_out_45_2) );
ms00f80 x_out_45_reg_30_ ( .ck(ispd_clk), .d(n_26760), .o(x_out_45_30) );
ms00f80 x_out_45_reg_31_ ( .ck(ispd_clk), .d(n_27146), .o(x_out_45_31) );
ms00f80 x_out_45_reg_32_ ( .ck(ispd_clk), .d(n_27640), .o(x_out_45_32) );
ms00f80 x_out_45_reg_33_ ( .ck(ispd_clk), .d(n_27641), .o(x_out_45_33) );
ms00f80 x_out_45_reg_3_ ( .ck(ispd_clk), .d(n_20956), .o(x_out_45_3) );
ms00f80 x_out_45_reg_4_ ( .ck(ispd_clk), .d(n_22284), .o(x_out_45_4) );
ms00f80 x_out_45_reg_5_ ( .ck(ispd_clk), .d(n_22957), .o(x_out_45_5) );
ms00f80 x_out_45_reg_6_ ( .ck(ispd_clk), .d(n_23936), .o(x_out_45_6) );
ms00f80 x_out_45_reg_7_ ( .ck(ispd_clk), .d(n_25282), .o(x_out_45_7) );
ms00f80 x_out_45_reg_8_ ( .ck(ispd_clk), .d(n_26450), .o(x_out_45_8) );
ms00f80 x_out_45_reg_9_ ( .ck(ispd_clk), .d(n_27260), .o(x_out_45_9) );
ms00f80 x_out_46_reg_0_ ( .ck(ispd_clk), .d(n_8617), .o(x_out_46_0) );
ms00f80 x_out_46_reg_10_ ( .ck(ispd_clk), .d(n_27261), .o(x_out_46_10) );
ms00f80 x_out_46_reg_11_ ( .ck(ispd_clk), .d(n_28010), .o(x_out_46_11) );
ms00f80 x_out_46_reg_12_ ( .ck(ispd_clk), .d(n_28422), .o(x_out_46_12) );
ms00f80 x_out_46_reg_13_ ( .ck(ispd_clk), .d(n_28866), .o(x_out_46_13) );
ms00f80 x_out_46_reg_14_ ( .ck(ispd_clk), .d(n_29205), .o(x_out_46_14) );
ms00f80 x_out_46_reg_15_ ( .ck(ispd_clk), .d(n_29492), .o(x_out_46_15) );
ms00f80 x_out_46_reg_18_ ( .ck(ispd_clk), .d(n_11417), .o(x_out_46_18) );
ms00f80 x_out_46_reg_19_ ( .ck(ispd_clk), .d(n_16969), .o(x_out_46_19) );
ms00f80 x_out_46_reg_1_ ( .ck(ispd_clk), .d(n_15448), .o(x_out_46_1) );
ms00f80 x_out_46_reg_20_ ( .ck(ispd_clk), .d(n_17600), .o(x_out_46_20) );
ms00f80 x_out_46_reg_21_ ( .ck(ispd_clk), .d(n_18144), .o(x_out_46_21) );
ms00f80 x_out_46_reg_22_ ( .ck(ispd_clk), .d(n_18791), .o(x_out_46_22) );
ms00f80 x_out_46_reg_23_ ( .ck(ispd_clk), .d(n_19512), .o(x_out_46_23) );
ms00f80 x_out_46_reg_24_ ( .ck(ispd_clk), .d(n_20659), .o(x_out_46_24) );
ms00f80 x_out_46_reg_25_ ( .ck(ispd_clk), .d(n_21405), .o(x_out_46_25) );
ms00f80 x_out_46_reg_26_ ( .ck(ispd_clk), .d(n_22428), .o(x_out_46_26) );
ms00f80 x_out_46_reg_27_ ( .ck(ispd_clk), .d(n_23408), .o(x_out_46_27) );
ms00f80 x_out_46_reg_28_ ( .ck(ispd_clk), .d(n_24361), .o(x_out_46_28) );
ms00f80 x_out_46_reg_29_ ( .ck(ispd_clk), .d(n_25400), .o(x_out_46_29) );
ms00f80 x_out_46_reg_2_ ( .ck(ispd_clk), .d(n_16432), .o(x_out_46_2) );
ms00f80 x_out_46_reg_30_ ( .ck(ispd_clk), .d(n_26306), .o(x_out_46_30) );
ms00f80 x_out_46_reg_31_ ( .ck(ispd_clk), .d(n_26621), .o(x_out_46_31) );
ms00f80 x_out_46_reg_32_ ( .ck(ispd_clk), .d(n_27001), .o(x_out_46_32) );
ms00f80 x_out_46_reg_33_ ( .ck(ispd_clk), .d(n_27000), .o(x_out_46_33) );
ms00f80 x_out_46_reg_3_ ( .ck(ispd_clk), .d(n_20176), .o(x_out_46_3) );
ms00f80 x_out_46_reg_4_ ( .ck(ispd_clk), .d(n_21196), .o(x_out_46_4) );
ms00f80 x_out_46_reg_5_ ( .ck(ispd_clk), .d(n_22017), .o(x_out_46_5) );
ms00f80 x_out_46_reg_6_ ( .ck(ispd_clk), .d(n_22642), .o(x_out_46_6) );
ms00f80 x_out_46_reg_7_ ( .ck(ispd_clk), .d(n_23934), .o(x_out_46_7) );
ms00f80 x_out_46_reg_8_ ( .ck(ispd_clk), .d(n_25280), .o(x_out_46_8) );
ms00f80 x_out_46_reg_9_ ( .ck(ispd_clk), .d(n_26449), .o(x_out_46_9) );
ms00f80 x_out_47_reg_0_ ( .ck(ispd_clk), .d(n_17519), .o(x_out_47_0) );
ms00f80 x_out_47_reg_10_ ( .ck(ispd_clk), .d(n_28668), .o(x_out_47_10) );
ms00f80 x_out_47_reg_11_ ( .ck(ispd_clk), .d(n_29020), .o(x_out_47_11) );
ms00f80 x_out_47_reg_12_ ( .ck(ispd_clk), .d(n_29394), .o(x_out_47_12) );
ms00f80 x_out_47_reg_13_ ( .ck(ispd_clk), .d(n_29585), .o(x_out_47_13) );
ms00f80 x_out_47_reg_14_ ( .ck(ispd_clk), .d(n_29672), .o(x_out_47_14) );
ms00f80 x_out_47_reg_15_ ( .ck(ispd_clk), .d(n_29706), .o(x_out_47_15) );
ms00f80 x_out_47_reg_18_ ( .ck(ispd_clk), .d(n_15758), .o(x_out_47_18) );
ms00f80 x_out_47_reg_19_ ( .ck(ispd_clk), .d(n_17863), .o(x_out_47_19) );
ms00f80 x_out_47_reg_1_ ( .ck(ispd_clk), .d(n_20909), .o(x_out_47_1) );
ms00f80 x_out_47_reg_20_ ( .ck(ispd_clk), .d(n_19112), .o(x_out_47_20) );
ms00f80 x_out_47_reg_21_ ( .ck(ispd_clk), .d(n_19841), .o(x_out_47_21) );
ms00f80 x_out_47_reg_22_ ( .ck(ispd_clk), .d(n_20666), .o(x_out_47_22) );
ms00f80 x_out_47_reg_23_ ( .ck(ispd_clk), .d(n_21083), .o(x_out_47_23) );
ms00f80 x_out_47_reg_24_ ( .ck(ispd_clk), .d(n_22431), .o(x_out_47_24) );
ms00f80 x_out_47_reg_25_ ( .ck(ispd_clk), .d(n_23136), .o(x_out_47_25) );
ms00f80 x_out_47_reg_26_ ( .ck(ispd_clk), .d(n_24364), .o(x_out_47_26) );
ms00f80 x_out_47_reg_27_ ( .ck(ispd_clk), .d(n_24822), .o(x_out_47_27) );
ms00f80 x_out_47_reg_28_ ( .ck(ispd_clk), .d(n_26014), .o(x_out_47_28) );
ms00f80 x_out_47_reg_29_ ( .ck(ispd_clk), .d(n_26688), .o(x_out_47_29) );
ms00f80 x_out_47_reg_2_ ( .ck(ispd_clk), .d(n_22278), .o(x_out_47_2) );
ms00f80 x_out_47_reg_30_ ( .ck(ispd_clk), .d(n_27566), .o(x_out_47_30) );
ms00f80 x_out_47_reg_31_ ( .ck(ispd_clk), .d(n_27935), .o(x_out_47_31) );
ms00f80 x_out_47_reg_32_ ( .ck(ispd_clk), .d(n_27990), .o(x_out_47_32) );
ms00f80 x_out_47_reg_33_ ( .ck(ispd_clk), .d(n_27987), .o(x_out_47_33) );
ms00f80 x_out_47_reg_3_ ( .ck(ispd_clk), .d(n_22950), .o(x_out_47_3) );
ms00f80 x_out_47_reg_4_ ( .ck(ispd_clk), .d(n_23326), .o(x_out_47_4) );
ms00f80 x_out_47_reg_5_ ( .ck(ispd_clk), .d(n_24624), .o(x_out_47_5) );
ms00f80 x_out_47_reg_6_ ( .ck(ispd_clk), .d(n_25908), .o(x_out_47_6) );
ms00f80 x_out_47_reg_7_ ( .ck(ispd_clk), .d(n_26814), .o(x_out_47_7) );
ms00f80 x_out_47_reg_8_ ( .ck(ispd_clk), .d(n_27720), .o(x_out_47_8) );
ms00f80 x_out_47_reg_9_ ( .ck(ispd_clk), .d(n_28321), .o(x_out_47_9) );
ms00f80 x_out_48_reg_0_ ( .ck(ispd_clk), .d(n_15570), .o(x_out_48_0) );
ms00f80 x_out_48_reg_10_ ( .ck(ispd_clk), .d(n_28320), .o(x_out_48_10) );
ms00f80 x_out_48_reg_11_ ( .ck(ispd_clk), .d(n_28691), .o(x_out_48_11) );
ms00f80 x_out_48_reg_12_ ( .ck(ispd_clk), .d(n_29049), .o(x_out_48_12) );
ms00f80 x_out_48_reg_13_ ( .ck(ispd_clk), .d(n_29349), .o(x_out_48_13) );
ms00f80 x_out_48_reg_14_ ( .ck(ispd_clk), .d(n_29601), .o(x_out_48_14) );
ms00f80 x_out_48_reg_15_ ( .ck(ispd_clk), .d(n_29693), .o(x_out_48_15) );
ms00f80 x_out_48_reg_18_ ( .ck(ispd_clk), .d(n_11472), .o(x_out_48_18) );
ms00f80 x_out_48_reg_19_ ( .ck(ispd_clk), .d(n_16777), .o(x_out_48_19) );
ms00f80 x_out_48_reg_1_ ( .ck(ispd_clk), .d(n_19751), .o(x_out_48_1) );
ms00f80 x_out_48_reg_20_ ( .ck(ispd_clk), .d(n_17376), .o(x_out_48_20) );
ms00f80 x_out_48_reg_21_ ( .ck(ispd_clk), .d(n_17928), .o(x_out_48_21) );
ms00f80 x_out_48_reg_22_ ( .ck(ispd_clk), .d(n_18532), .o(x_out_48_22) );
ms00f80 x_out_48_reg_23_ ( .ck(ispd_clk), .d(n_19164), .o(x_out_48_23) );
ms00f80 x_out_48_reg_24_ ( .ck(ispd_clk), .d(n_20228), .o(x_out_48_24) );
ms00f80 x_out_48_reg_25_ ( .ck(ispd_clk), .d(n_21326), .o(x_out_48_25) );
ms00f80 x_out_48_reg_26_ ( .ck(ispd_clk), .d(n_22112), .o(x_out_48_26) );
ms00f80 x_out_48_reg_27_ ( .ck(ispd_clk), .d(n_23079), .o(x_out_48_27) );
ms00f80 x_out_48_reg_28_ ( .ck(ispd_clk), .d(n_24040), .o(x_out_48_28) );
ms00f80 x_out_48_reg_29_ ( .ck(ispd_clk), .d(n_25038), .o(x_out_48_29) );
ms00f80 x_out_48_reg_2_ ( .ck(ispd_clk), .d(n_20504), .o(x_out_48_2) );
ms00f80 x_out_48_reg_30_ ( .ck(ispd_clk), .d(n_25743), .o(x_out_48_30) );
ms00f80 x_out_48_reg_31_ ( .ck(ispd_clk), .d(n_26023), .o(x_out_48_31) );
ms00f80 x_out_48_reg_32_ ( .ck(ispd_clk), .d(n_26626), .o(x_out_48_32) );
ms00f80 x_out_48_reg_33_ ( .ck(ispd_clk), .d(n_26625), .o(x_out_48_33) );
ms00f80 x_out_48_reg_3_ ( .ck(ispd_clk), .d(n_21611), .o(x_out_48_3) );
ms00f80 x_out_48_reg_4_ ( .ck(ispd_clk), .d(n_22314), .o(x_out_48_4) );
ms00f80 x_out_48_reg_5_ ( .ck(ispd_clk), .d(n_23325), .o(x_out_48_5) );
ms00f80 x_out_48_reg_6_ ( .ck(ispd_clk), .d(n_24623), .o(x_out_48_6) );
ms00f80 x_out_48_reg_7_ ( .ck(ispd_clk), .d(n_25907), .o(x_out_48_7) );
ms00f80 x_out_48_reg_8_ ( .ck(ispd_clk), .d(n_26812), .o(x_out_48_8) );
ms00f80 x_out_48_reg_9_ ( .ck(ispd_clk), .d(n_27719), .o(x_out_48_9) );
ms00f80 x_out_49_reg_0_ ( .ck(ispd_clk), .d(n_16373), .o(x_out_49_0) );
ms00f80 x_out_49_reg_10_ ( .ck(ispd_clk), .d(n_28319), .o(x_out_49_10) );
ms00f80 x_out_49_reg_11_ ( .ck(ispd_clk), .d(n_28690), .o(x_out_49_11) );
ms00f80 x_out_49_reg_12_ ( .ck(ispd_clk), .d(n_29045), .o(x_out_49_12) );
ms00f80 x_out_49_reg_13_ ( .ck(ispd_clk), .d(n_29346), .o(x_out_49_13) );
ms00f80 x_out_49_reg_14_ ( .ck(ispd_clk), .d(n_29600), .o(x_out_49_14) );
ms00f80 x_out_49_reg_15_ ( .ck(ispd_clk), .d(n_29692), .o(x_out_49_15) );
ms00f80 x_out_49_reg_18_ ( .ck(ispd_clk), .d(n_16647), .o(x_out_49_18) );
ms00f80 x_out_49_reg_19_ ( .ck(ispd_clk), .d(n_17624), .o(x_out_49_19) );
ms00f80 x_out_49_reg_1_ ( .ck(ispd_clk), .d(n_19750), .o(x_out_49_1) );
ms00f80 x_out_49_reg_20_ ( .ck(ispd_clk), .d(n_19111), .o(x_out_49_20) );
ms00f80 x_out_49_reg_21_ ( .ck(ispd_clk), .d(n_20189), .o(x_out_49_21) );
ms00f80 x_out_49_reg_22_ ( .ck(ispd_clk), .d(n_21268), .o(x_out_49_22) );
ms00f80 x_out_49_reg_23_ ( .ck(ispd_clk), .d(n_22073), .o(x_out_49_23) );
ms00f80 x_out_49_reg_24_ ( .ck(ispd_clk), .d(n_23057), .o(x_out_49_24) );
ms00f80 x_out_49_reg_25_ ( .ck(ispd_clk), .d(n_24022), .o(x_out_49_25) );
ms00f80 x_out_49_reg_26_ ( .ck(ispd_clk), .d(n_25025), .o(x_out_49_26) );
ms00f80 x_out_49_reg_27_ ( .ck(ispd_clk), .d(n_25731), .o(x_out_49_27) );
ms00f80 x_out_49_reg_28_ ( .ck(ispd_clk), .d(n_26603), .o(x_out_49_28) );
ms00f80 x_out_49_reg_29_ ( .ck(ispd_clk), .d(n_27399), .o(x_out_49_29) );
ms00f80 x_out_49_reg_2_ ( .ck(ispd_clk), .d(n_20503), .o(x_out_49_2) );
ms00f80 x_out_49_reg_30_ ( .ck(ispd_clk), .d(n_27650), .o(x_out_49_30) );
ms00f80 x_out_49_reg_31_ ( .ck(ispd_clk), .d(n_27751), .o(x_out_49_31) );
ms00f80 x_out_49_reg_32_ ( .ck(ispd_clk), .d(n_27752), .o(x_out_49_32) );
ms00f80 x_out_49_reg_33_ ( .ck(ispd_clk), .d(n_27749), .o(x_out_49_33) );
ms00f80 x_out_49_reg_3_ ( .ck(ispd_clk), .d(n_21610), .o(x_out_49_3) );
ms00f80 x_out_49_reg_4_ ( .ck(ispd_clk), .d(n_22312), .o(x_out_49_4) );
ms00f80 x_out_49_reg_5_ ( .ck(ispd_clk), .d(n_23324), .o(x_out_49_5) );
ms00f80 x_out_49_reg_6_ ( .ck(ispd_clk), .d(n_24621), .o(x_out_49_6) );
ms00f80 x_out_49_reg_7_ ( .ck(ispd_clk), .d(n_25902), .o(x_out_49_7) );
ms00f80 x_out_49_reg_8_ ( .ck(ispd_clk), .d(n_26811), .o(x_out_49_8) );
ms00f80 x_out_49_reg_9_ ( .ck(ispd_clk), .d(n_27716), .o(x_out_49_9) );
ms00f80 x_out_4_reg_0_ ( .ck(ispd_clk), .d(n_11174), .o(x_out_4_0) );
ms00f80 x_out_4_reg_10_ ( .ck(ispd_clk), .d(n_26415), .o(x_out_4_10) );
ms00f80 x_out_4_reg_11_ ( .ck(ispd_clk), .d(n_27252), .o(x_out_4_11) );
ms00f80 x_out_4_reg_12_ ( .ck(ispd_clk), .d(n_27998), .o(x_out_4_12) );
ms00f80 x_out_4_reg_13_ ( .ck(ispd_clk), .d(n_28515), .o(x_out_4_13) );
ms00f80 x_out_4_reg_14_ ( .ck(ispd_clk), .d(n_28853), .o(x_out_4_14) );
ms00f80 x_out_4_reg_15_ ( .ck(ispd_clk), .d(n_29180), .o(x_out_4_15) );
ms00f80 x_out_4_reg_18_ ( .ck(ispd_clk), .d(n_11076), .o(x_out_4_18) );
ms00f80 x_out_4_reg_19_ ( .ck(ispd_clk), .d(n_15757), .o(x_out_4_19) );
ms00f80 x_out_4_reg_1_ ( .ck(ispd_clk), .d(n_15455), .o(x_out_4_1) );
ms00f80 x_out_4_reg_20_ ( .ck(ispd_clk), .d(n_15716), .o(x_out_4_20) );
ms00f80 x_out_4_reg_21_ ( .ck(ispd_clk), .d(n_16228), .o(x_out_4_21) );
ms00f80 x_out_4_reg_22_ ( .ck(ispd_clk), .d(n_16930), .o(x_out_4_22) );
ms00f80 x_out_4_reg_23_ ( .ck(ispd_clk), .d(n_18152), .o(x_out_4_23) );
ms00f80 x_out_4_reg_24_ ( .ck(ispd_clk), .d(n_18853), .o(x_out_4_24) );
ms00f80 x_out_4_reg_25_ ( .ck(ispd_clk), .d(n_20227), .o(x_out_4_25) );
ms00f80 x_out_4_reg_26_ ( .ck(ispd_clk), .d(n_21011), .o(x_out_4_26) );
ms00f80 x_out_4_reg_27_ ( .ck(ispd_clk), .d(n_22110), .o(x_out_4_27) );
ms00f80 x_out_4_reg_28_ ( .ck(ispd_clk), .d(n_22755), .o(x_out_4_28) );
ms00f80 x_out_4_reg_29_ ( .ck(ispd_clk), .d(n_24039), .o(x_out_4_29) );
ms00f80 x_out_4_reg_2_ ( .ck(ispd_clk), .d(n_17192), .o(x_out_4_2) );
ms00f80 x_out_4_reg_30_ ( .ck(ispd_clk), .d(n_24325), .o(x_out_4_30) );
ms00f80 x_out_4_reg_31_ ( .ck(ispd_clk), .d(n_25707), .o(x_out_4_31) );
ms00f80 x_out_4_reg_32_ ( .ck(ispd_clk), .d(n_26931), .o(x_out_4_32) );
ms00f80 x_out_4_reg_33_ ( .ck(ispd_clk), .d(n_26930), .o(x_out_4_33) );
ms00f80 x_out_4_reg_3_ ( .ck(ispd_clk), .d(n_18686), .o(x_out_4_3) );
ms00f80 x_out_4_reg_4_ ( .ck(ispd_clk), .d(n_18801), .o(x_out_4_4) );
ms00f80 x_out_4_reg_5_ ( .ck(ispd_clk), .d(n_20188), .o(x_out_4_5) );
ms00f80 x_out_4_reg_6_ ( .ck(ispd_clk), .d(n_21609), .o(x_out_4_6) );
ms00f80 x_out_4_reg_7_ ( .ck(ispd_clk), .d(n_22621), .o(x_out_4_7) );
ms00f80 x_out_4_reg_8_ ( .ck(ispd_clk), .d(n_23922), .o(x_out_4_8) );
ms00f80 x_out_4_reg_9_ ( .ck(ispd_clk), .d(n_25257), .o(x_out_4_9) );
ms00f80 x_out_50_reg_0_ ( .ck(ispd_clk), .d(n_15221), .o(x_out_50_0) );
ms00f80 x_out_50_reg_10_ ( .ck(ispd_clk), .d(n_28318), .o(x_out_50_10) );
ms00f80 x_out_50_reg_11_ ( .ck(ispd_clk), .d(n_28689), .o(x_out_50_11) );
ms00f80 x_out_50_reg_12_ ( .ck(ispd_clk), .d(n_29043), .o(x_out_50_12) );
ms00f80 x_out_50_reg_13_ ( .ck(ispd_clk), .d(n_29344), .o(x_out_50_13) );
ms00f80 x_out_50_reg_14_ ( .ck(ispd_clk), .d(n_29598), .o(x_out_50_14) );
ms00f80 x_out_50_reg_15_ ( .ck(ispd_clk), .d(n_29689), .o(x_out_50_15) );
ms00f80 x_out_50_reg_18_ ( .ck(ispd_clk), .d(n_13854), .o(x_out_50_18) );
ms00f80 x_out_50_reg_19_ ( .ck(ispd_clk), .d(n_17516), .o(x_out_50_19) );
ms00f80 x_out_50_reg_1_ ( .ck(ispd_clk), .d(n_19443), .o(x_out_50_1) );
ms00f80 x_out_50_reg_20_ ( .ck(ispd_clk), .d(n_17847), .o(x_out_50_20) );
ms00f80 x_out_50_reg_21_ ( .ck(ispd_clk), .d(n_18531), .o(x_out_50_21) );
ms00f80 x_out_50_reg_22_ ( .ck(ispd_clk), .d(n_19515), .o(x_out_50_22) );
ms00f80 x_out_50_reg_23_ ( .ck(ispd_clk), .d(n_20664), .o(x_out_50_23) );
ms00f80 x_out_50_reg_24_ ( .ck(ispd_clk), .d(n_21407), .o(x_out_50_24) );
ms00f80 x_out_50_reg_25_ ( .ck(ispd_clk), .d(n_22430), .o(x_out_50_25) );
ms00f80 x_out_50_reg_26_ ( .ck(ispd_clk), .d(n_23410), .o(x_out_50_26) );
ms00f80 x_out_50_reg_27_ ( .ck(ispd_clk), .d(n_24363), .o(x_out_50_27) );
ms00f80 x_out_50_reg_28_ ( .ck(ispd_clk), .d(n_25096), .o(x_out_50_28) );
ms00f80 x_out_50_reg_29_ ( .ck(ispd_clk), .d(n_26013), .o(x_out_50_29) );
ms00f80 x_out_50_reg_2_ ( .ck(ispd_clk), .d(n_20892), .o(x_out_50_2) );
ms00f80 x_out_50_reg_30_ ( .ck(ispd_clk), .d(n_26349), .o(x_out_50_30) );
ms00f80 x_out_50_reg_31_ ( .ck(ispd_clk), .d(n_27453), .o(x_out_50_31) );
ms00f80 x_out_50_reg_32_ ( .ck(ispd_clk), .d(n_27451), .o(x_out_50_32) );
ms00f80 x_out_50_reg_33_ ( .ck(ispd_clk), .d(n_27448), .o(x_out_50_33) );
ms00f80 x_out_50_reg_3_ ( .ck(ispd_clk), .d(n_21998), .o(x_out_50_3) );
ms00f80 x_out_50_reg_4_ ( .ck(ispd_clk), .d(n_22072), .o(x_out_50_4) );
ms00f80 x_out_50_reg_5_ ( .ck(ispd_clk), .d(n_23323), .o(x_out_50_5) );
ms00f80 x_out_50_reg_6_ ( .ck(ispd_clk), .d(n_24620), .o(x_out_50_6) );
ms00f80 x_out_50_reg_7_ ( .ck(ispd_clk), .d(n_25900), .o(x_out_50_7) );
ms00f80 x_out_50_reg_8_ ( .ck(ispd_clk), .d(n_26810), .o(x_out_50_8) );
ms00f80 x_out_50_reg_9_ ( .ck(ispd_clk), .d(n_27713), .o(x_out_50_9) );
ms00f80 x_out_51_reg_0_ ( .ck(ispd_clk), .d(n_15855), .o(x_out_51_0) );
ms00f80 x_out_51_reg_10_ ( .ck(ispd_clk), .d(n_28317), .o(x_out_51_10) );
ms00f80 x_out_51_reg_11_ ( .ck(ispd_clk), .d(n_28687), .o(x_out_51_11) );
ms00f80 x_out_51_reg_12_ ( .ck(ispd_clk), .d(n_29042), .o(x_out_51_12) );
ms00f80 x_out_51_reg_13_ ( .ck(ispd_clk), .d(n_29343), .o(x_out_51_13) );
ms00f80 x_out_51_reg_14_ ( .ck(ispd_clk), .d(n_29596), .o(x_out_51_14) );
ms00f80 x_out_51_reg_15_ ( .ck(ispd_clk), .d(n_29686), .o(x_out_51_15) );
ms00f80 x_out_51_reg_18_ ( .ck(ispd_clk), .d(n_17229), .o(x_out_51_18) );
ms00f80 x_out_51_reg_19_ ( .ck(ispd_clk), .d(n_18422), .o(x_out_51_19) );
ms00f80 x_out_51_reg_1_ ( .ck(ispd_clk), .d(n_19442), .o(x_out_51_1) );
ms00f80 x_out_51_reg_20_ ( .ck(ispd_clk), .d(n_19284), .o(x_out_51_20) );
ms00f80 x_out_51_reg_21_ ( .ck(ispd_clk), .d(n_20321), .o(x_out_51_21) );
ms00f80 x_out_51_reg_22_ ( .ck(ispd_clk), .d(n_21406), .o(x_out_51_22) );
ms00f80 x_out_51_reg_23_ ( .ck(ispd_clk), .d(n_22160), .o(x_out_51_23) );
ms00f80 x_out_51_reg_24_ ( .ck(ispd_clk), .d(n_23409), .o(x_out_51_24) );
ms00f80 x_out_51_reg_25_ ( .ck(ispd_clk), .d(n_24091), .o(x_out_51_25) );
ms00f80 x_out_51_reg_26_ ( .ck(ispd_clk), .d(n_25095), .o(x_out_51_26) );
ms00f80 x_out_51_reg_27_ ( .ck(ispd_clk), .d(n_25800), .o(x_out_51_27) );
ms00f80 x_out_51_reg_28_ ( .ck(ispd_clk), .d(n_27209), .o(x_out_51_28) );
ms00f80 x_out_51_reg_29_ ( .ck(ispd_clk), .d(n_27447), .o(x_out_51_29) );
ms00f80 x_out_51_reg_2_ ( .ck(ispd_clk), .d(n_20891), .o(x_out_51_2) );
ms00f80 x_out_51_reg_30_ ( .ck(ispd_clk), .d(n_27895), .o(x_out_51_30) );
ms00f80 x_out_51_reg_31_ ( .ck(ispd_clk), .d(n_27897), .o(x_out_51_31) );
ms00f80 x_out_51_reg_32_ ( .ck(ispd_clk), .d(n_27893), .o(x_out_51_32) );
ms00f80 x_out_51_reg_33_ ( .ck(ispd_clk), .d(n_27892), .o(x_out_51_33) );
ms00f80 x_out_51_reg_3_ ( .ck(ispd_clk), .d(n_21997), .o(x_out_51_3) );
ms00f80 x_out_51_reg_4_ ( .ck(ispd_clk), .d(n_22070), .o(x_out_51_4) );
ms00f80 x_out_51_reg_5_ ( .ck(ispd_clk), .d(n_23322), .o(x_out_51_5) );
ms00f80 x_out_51_reg_6_ ( .ck(ispd_clk), .d(n_24619), .o(x_out_51_6) );
ms00f80 x_out_51_reg_7_ ( .ck(ispd_clk), .d(n_25899), .o(x_out_51_7) );
ms00f80 x_out_51_reg_8_ ( .ck(ispd_clk), .d(n_26809), .o(x_out_51_8) );
ms00f80 x_out_51_reg_9_ ( .ck(ispd_clk), .d(n_27711), .o(x_out_51_9) );
ms00f80 x_out_52_reg_0_ ( .ck(ispd_clk), .d(n_15852), .o(x_out_52_0) );
ms00f80 x_out_52_reg_10_ ( .ck(ispd_clk), .d(n_28220), .o(x_out_52_10) );
ms00f80 x_out_52_reg_11_ ( .ck(ispd_clk), .d(n_28622), .o(x_out_52_11) );
ms00f80 x_out_52_reg_12_ ( .ck(ispd_clk), .d(n_28929), .o(x_out_52_12) );
ms00f80 x_out_52_reg_13_ ( .ck(ispd_clk), .d(n_29268), .o(x_out_52_13) );
ms00f80 x_out_52_reg_14_ ( .ck(ispd_clk), .d(n_29532), .o(x_out_52_14) );
ms00f80 x_out_52_reg_15_ ( .ck(ispd_clk), .d(n_29670), .o(x_out_52_15) );
ms00f80 x_out_52_reg_1_ ( .ck(ispd_clk), .d(n_19163), .o(x_out_52_1) );
ms00f80 x_out_52_reg_2_ ( .ck(ispd_clk), .d(n_20502), .o(x_out_52_2) );
ms00f80 x_out_52_reg_3_ ( .ck(ispd_clk), .d(n_21607), .o(x_out_52_3) );
ms00f80 x_out_52_reg_4_ ( .ck(ispd_clk), .d(n_21773), .o(x_out_52_4) );
ms00f80 x_out_52_reg_5_ ( .ck(ispd_clk), .d(n_23055), .o(x_out_52_5) );
ms00f80 x_out_52_reg_6_ ( .ck(ispd_clk), .d(n_24309), .o(x_out_52_6) );
ms00f80 x_out_52_reg_7_ ( .ck(ispd_clk), .d(n_25682), .o(x_out_52_7) );
ms00f80 x_out_52_reg_8_ ( .ck(ispd_clk), .d(n_26538), .o(x_out_52_8) );
ms00f80 x_out_52_reg_9_ ( .ck(ispd_clk), .d(n_27561), .o(x_out_52_9) );
ms00f80 x_out_53_reg_0_ ( .ck(ispd_clk), .d(n_15860), .o(x_out_53_0) );
ms00f80 x_out_53_reg_10_ ( .ck(ispd_clk), .d(n_28219), .o(x_out_53_10) );
ms00f80 x_out_53_reg_11_ ( .ck(ispd_clk), .d(n_28619), .o(x_out_53_11) );
ms00f80 x_out_53_reg_12_ ( .ck(ispd_clk), .d(n_28926), .o(x_out_53_12) );
ms00f80 x_out_53_reg_13_ ( .ck(ispd_clk), .d(n_29265), .o(x_out_53_13) );
ms00f80 x_out_53_reg_14_ ( .ck(ispd_clk), .d(n_29530), .o(x_out_53_14) );
ms00f80 x_out_53_reg_15_ ( .ck(ispd_clk), .d(n_29667), .o(x_out_53_15) );
ms00f80 x_out_53_reg_18_ ( .ck(ispd_clk), .d(n_6482), .o(x_out_53_18) );
ms00f80 x_out_53_reg_19_ ( .ck(ispd_clk), .d(n_7224), .o(x_out_53_19) );
ms00f80 x_out_53_reg_1_ ( .ck(ispd_clk), .d(n_19162), .o(x_out_53_1) );
ms00f80 x_out_53_reg_20_ ( .ck(ispd_clk), .d(n_7416), .o(x_out_53_20) );
ms00f80 x_out_53_reg_21_ ( .ck(ispd_clk), .d(n_8004), .o(x_out_53_21) );
ms00f80 x_out_53_reg_22_ ( .ck(ispd_clk), .d(n_9210), .o(x_out_53_22) );
ms00f80 x_out_53_reg_23_ ( .ck(ispd_clk), .d(n_11026), .o(x_out_53_23) );
ms00f80 x_out_53_reg_24_ ( .ck(ispd_clk), .d(n_12145), .o(x_out_53_24) );
ms00f80 x_out_53_reg_25_ ( .ck(ispd_clk), .d(n_13359), .o(x_out_53_25) );
ms00f80 x_out_53_reg_26_ ( .ck(ispd_clk), .d(n_14522), .o(x_out_53_26) );
ms00f80 x_out_53_reg_27_ ( .ck(ispd_clk), .d(n_15191), .o(x_out_53_27) );
ms00f80 x_out_53_reg_28_ ( .ck(ispd_clk), .d(n_15927), .o(x_out_53_28) );
ms00f80 x_out_53_reg_29_ ( .ck(ispd_clk), .d(n_16283), .o(x_out_53_29) );
ms00f80 x_out_53_reg_2_ ( .ck(ispd_clk), .d(n_20501), .o(x_out_53_2) );
ms00f80 x_out_53_reg_30_ ( .ck(ispd_clk), .d(n_15964), .o(x_out_53_30) );
ms00f80 x_out_53_reg_31_ ( .ck(ispd_clk), .d(n_15968), .o(x_out_53_31) );
ms00f80 x_out_53_reg_32_ ( .ck(ispd_clk), .d(n_15966), .o(x_out_53_32) );
ms00f80 x_out_53_reg_33_ ( .ck(ispd_clk), .d(n_15965), .o(x_out_53_33) );
ms00f80 x_out_53_reg_3_ ( .ck(ispd_clk), .d(n_21606), .o(x_out_53_3) );
ms00f80 x_out_53_reg_4_ ( .ck(ispd_clk), .d(n_21772), .o(x_out_53_4) );
ms00f80 x_out_53_reg_5_ ( .ck(ispd_clk), .d(n_23054), .o(x_out_53_5) );
ms00f80 x_out_53_reg_6_ ( .ck(ispd_clk), .d(n_24308), .o(x_out_53_6) );
ms00f80 x_out_53_reg_7_ ( .ck(ispd_clk), .d(n_25681), .o(x_out_53_7) );
ms00f80 x_out_53_reg_8_ ( .ck(ispd_clk), .d(n_26537), .o(x_out_53_8) );
ms00f80 x_out_53_reg_9_ ( .ck(ispd_clk), .d(n_27560), .o(x_out_53_9) );
ms00f80 x_out_54_reg_0_ ( .ck(ispd_clk), .d(n_15848), .o(x_out_54_0) );
ms00f80 x_out_54_reg_10_ ( .ck(ispd_clk), .d(n_28218), .o(x_out_54_10) );
ms00f80 x_out_54_reg_11_ ( .ck(ispd_clk), .d(n_28617), .o(x_out_54_11) );
ms00f80 x_out_54_reg_12_ ( .ck(ispd_clk), .d(n_28925), .o(x_out_54_12) );
ms00f80 x_out_54_reg_13_ ( .ck(ispd_clk), .d(n_29263), .o(x_out_54_13) );
ms00f80 x_out_54_reg_14_ ( .ck(ispd_clk), .d(n_29528), .o(x_out_54_14) );
ms00f80 x_out_54_reg_15_ ( .ck(ispd_clk), .d(n_29684), .o(x_out_54_15) );
ms00f80 x_out_54_reg_18_ ( .ck(ispd_clk), .d(n_7257), .o(x_out_54_18) );
ms00f80 x_out_54_reg_19_ ( .ck(ispd_clk), .d(n_7411), .o(x_out_54_19) );
ms00f80 x_out_54_reg_1_ ( .ck(ispd_clk), .d(n_19440), .o(x_out_54_1) );
ms00f80 x_out_54_reg_20_ ( .ck(ispd_clk), .d(n_6691), .o(x_out_54_20) );
ms00f80 x_out_54_reg_21_ ( .ck(ispd_clk), .d(n_8003), .o(x_out_54_21) );
ms00f80 x_out_54_reg_22_ ( .ck(ispd_clk), .d(n_9212), .o(x_out_54_22) );
ms00f80 x_out_54_reg_23_ ( .ck(ispd_clk), .d(n_11025), .o(x_out_54_23) );
ms00f80 x_out_54_reg_24_ ( .ck(ispd_clk), .d(n_12144), .o(x_out_54_24) );
ms00f80 x_out_54_reg_25_ ( .ck(ispd_clk), .d(n_13358), .o(x_out_54_25) );
ms00f80 x_out_54_reg_26_ ( .ck(ispd_clk), .d(n_14521), .o(x_out_54_26) );
ms00f80 x_out_54_reg_27_ ( .ck(ispd_clk), .d(n_15190), .o(x_out_54_27) );
ms00f80 x_out_54_reg_28_ ( .ck(ispd_clk), .d(n_15943), .o(x_out_54_28) );
ms00f80 x_out_54_reg_29_ ( .ck(ispd_clk), .d(n_16278), .o(x_out_54_29) );
ms00f80 x_out_54_reg_2_ ( .ck(ispd_clk), .d(n_20186), .o(x_out_54_2) );
ms00f80 x_out_54_reg_30_ ( .ck(ispd_clk), .d(n_17067), .o(x_out_54_30) );
ms00f80 x_out_54_reg_31_ ( .ck(ispd_clk), .d(n_16799), .o(x_out_54_31) );
ms00f80 x_out_54_reg_32_ ( .ck(ispd_clk), .d(n_16778), .o(x_out_54_32) );
ms00f80 x_out_54_reg_33_ ( .ck(ispd_clk), .d(n_16797), .o(x_out_54_33) );
ms00f80 x_out_54_reg_3_ ( .ck(ispd_clk), .d(n_21605), .o(x_out_54_3) );
ms00f80 x_out_54_reg_4_ ( .ck(ispd_clk), .d(n_22311), .o(x_out_54_4) );
ms00f80 x_out_54_reg_5_ ( .ck(ispd_clk), .d(n_23320), .o(x_out_54_5) );
ms00f80 x_out_54_reg_6_ ( .ck(ispd_clk), .d(n_24307), .o(x_out_54_6) );
ms00f80 x_out_54_reg_7_ ( .ck(ispd_clk), .d(n_25679), .o(x_out_54_7) );
ms00f80 x_out_54_reg_8_ ( .ck(ispd_clk), .d(n_26535), .o(x_out_54_8) );
ms00f80 x_out_54_reg_9_ ( .ck(ispd_clk), .d(n_27559), .o(x_out_54_9) );
ms00f80 x_out_55_reg_0_ ( .ck(ispd_clk), .d(n_16110), .o(x_out_55_0) );
ms00f80 x_out_55_reg_10_ ( .ck(ispd_clk), .d(n_28217), .o(x_out_55_10) );
ms00f80 x_out_55_reg_11_ ( .ck(ispd_clk), .d(n_28616), .o(x_out_55_11) );
ms00f80 x_out_55_reg_12_ ( .ck(ispd_clk), .d(n_28923), .o(x_out_55_12) );
ms00f80 x_out_55_reg_13_ ( .ck(ispd_clk), .d(n_29260), .o(x_out_55_13) );
ms00f80 x_out_55_reg_14_ ( .ck(ispd_clk), .d(n_29525), .o(x_out_55_14) );
ms00f80 x_out_55_reg_15_ ( .ck(ispd_clk), .d(n_29681), .o(x_out_55_15) );
ms00f80 x_out_55_reg_18_ ( .ck(ispd_clk), .d(n_13098), .o(x_out_55_18) );
ms00f80 x_out_55_reg_19_ ( .ck(ispd_clk), .d(n_15478), .o(x_out_55_19) );
ms00f80 x_out_55_reg_1_ ( .ck(ispd_clk), .d(n_19160), .o(x_out_55_1) );
ms00f80 x_out_55_reg_20_ ( .ck(ispd_clk), .d(n_16558), .o(x_out_55_20) );
ms00f80 x_out_55_reg_21_ ( .ck(ispd_clk), .d(n_17422), .o(x_out_55_21) );
ms00f80 x_out_55_reg_22_ ( .ck(ispd_clk), .d(n_18324), .o(x_out_55_22) );
ms00f80 x_out_55_reg_23_ ( .ck(ispd_clk), .d(n_19561), .o(x_out_55_23) );
ms00f80 x_out_55_reg_24_ ( .ck(ispd_clk), .d(n_20353), .o(x_out_55_24) );
ms00f80 x_out_55_reg_25_ ( .ck(ispd_clk), .d(n_21455), .o(x_out_55_25) );
ms00f80 x_out_55_reg_26_ ( .ck(ispd_clk), .d(n_22192), .o(x_out_55_26) );
ms00f80 x_out_55_reg_27_ ( .ck(ispd_clk), .d(n_23456), .o(x_out_55_27) );
ms00f80 x_out_55_reg_28_ ( .ck(ispd_clk), .d(n_24122), .o(x_out_55_28) );
ms00f80 x_out_55_reg_29_ ( .ck(ispd_clk), .d(n_25136), .o(x_out_55_29) );
ms00f80 x_out_55_reg_2_ ( .ck(ispd_clk), .d(n_20505), .o(x_out_55_2) );
ms00f80 x_out_55_reg_30_ ( .ck(ispd_clk), .d(n_25809), .o(x_out_55_30) );
ms00f80 x_out_55_reg_31_ ( .ck(ispd_clk), .d(n_25812), .o(x_out_55_31) );
ms00f80 x_out_55_reg_32_ ( .ck(ispd_clk), .d(n_25811), .o(x_out_55_32) );
ms00f80 x_out_55_reg_33_ ( .ck(ispd_clk), .d(n_25808), .o(x_out_55_33) );
ms00f80 x_out_55_reg_3_ ( .ck(ispd_clk), .d(n_21604), .o(x_out_55_3) );
ms00f80 x_out_55_reg_4_ ( .ck(ispd_clk), .d(n_21771), .o(x_out_55_4) );
ms00f80 x_out_55_reg_5_ ( .ck(ispd_clk), .d(n_23053), .o(x_out_55_5) );
ms00f80 x_out_55_reg_6_ ( .ck(ispd_clk), .d(n_24306), .o(x_out_55_6) );
ms00f80 x_out_55_reg_7_ ( .ck(ispd_clk), .d(n_25678), .o(x_out_55_7) );
ms00f80 x_out_55_reg_8_ ( .ck(ispd_clk), .d(n_26534), .o(x_out_55_8) );
ms00f80 x_out_55_reg_9_ ( .ck(ispd_clk), .d(n_27557), .o(x_out_55_9) );
ms00f80 x_out_56_reg_0_ ( .ck(ispd_clk), .d(n_16992), .o(x_out_56_0) );
ms00f80 x_out_56_reg_10_ ( .ck(ispd_clk), .d(n_28368), .o(x_out_56_10) );
ms00f80 x_out_56_reg_11_ ( .ck(ispd_clk), .d(n_28758), .o(x_out_56_11) );
ms00f80 x_out_56_reg_12_ ( .ck(ispd_clk), .d(n_29108), .o(x_out_56_12) );
ms00f80 x_out_56_reg_13_ ( .ck(ispd_clk), .d(n_29416), .o(x_out_56_13) );
ms00f80 x_out_56_reg_14_ ( .ck(ispd_clk), .d(n_29649), .o(x_out_56_14) );
ms00f80 x_out_56_reg_15_ ( .ck(ispd_clk), .d(n_29699), .o(x_out_56_15) );
ms00f80 x_out_56_reg_18_ ( .ck(ispd_clk), .d(n_7628), .o(x_out_56_18) );
ms00f80 x_out_56_reg_19_ ( .ck(ispd_clk), .d(n_6535), .o(x_out_56_19) );
ms00f80 x_out_56_reg_1_ ( .ck(ispd_clk), .d(n_20539), .o(x_out_56_1) );
ms00f80 x_out_56_reg_20_ ( .ck(ispd_clk), .d(n_6692), .o(x_out_56_20) );
ms00f80 x_out_56_reg_21_ ( .ck(ispd_clk), .d(n_7999), .o(x_out_56_21) );
ms00f80 x_out_56_reg_22_ ( .ck(ispd_clk), .d(n_9211), .o(x_out_56_22) );
ms00f80 x_out_56_reg_23_ ( .ck(ispd_clk), .d(n_11023), .o(x_out_56_23) );
ms00f80 x_out_56_reg_24_ ( .ck(ispd_clk), .d(n_12143), .o(x_out_56_24) );
ms00f80 x_out_56_reg_25_ ( .ck(ispd_clk), .d(n_13357), .o(x_out_56_25) );
ms00f80 x_out_56_reg_26_ ( .ck(ispd_clk), .d(n_14519), .o(x_out_56_26) );
ms00f80 x_out_56_reg_27_ ( .ck(ispd_clk), .d(n_15189), .o(x_out_56_27) );
ms00f80 x_out_56_reg_28_ ( .ck(ispd_clk), .d(n_15942), .o(x_out_56_28) );
ms00f80 x_out_56_reg_29_ ( .ck(ispd_clk), .d(n_16557), .o(x_out_56_29) );
ms00f80 x_out_56_reg_2_ ( .ck(ispd_clk), .d(n_21996), .o(x_out_56_2) );
ms00f80 x_out_56_reg_30_ ( .ck(ispd_clk), .d(n_16821), .o(x_out_56_30) );
ms00f80 x_out_56_reg_31_ ( .ck(ispd_clk), .d(n_17406), .o(x_out_56_31) );
ms00f80 x_out_56_reg_32_ ( .ck(ispd_clk), .d(n_17100), .o(x_out_56_32) );
ms00f80 x_out_56_reg_33_ ( .ck(ispd_clk), .d(n_17098), .o(x_out_56_33) );
ms00f80 x_out_56_reg_3_ ( .ck(ispd_clk), .d(n_22620), .o(x_out_56_3) );
ms00f80 x_out_56_reg_4_ ( .ck(ispd_clk), .d(n_23052), .o(x_out_56_4) );
ms00f80 x_out_56_reg_5_ ( .ck(ispd_clk), .d(n_24305), .o(x_out_56_5) );
ms00f80 x_out_56_reg_6_ ( .ck(ispd_clk), .d(n_25676), .o(x_out_56_6) );
ms00f80 x_out_56_reg_7_ ( .ck(ispd_clk), .d(n_26533), .o(x_out_56_7) );
ms00f80 x_out_56_reg_8_ ( .ck(ispd_clk), .d(n_27352), .o(x_out_56_8) );
ms00f80 x_out_56_reg_9_ ( .ck(ispd_clk), .d(n_27932), .o(x_out_56_9) );
ms00f80 x_out_57_reg_0_ ( .ck(ispd_clk), .d(n_8681), .o(x_out_57_0) );
ms00f80 x_out_57_reg_10_ ( .ck(ispd_clk), .d(n_27267), .o(x_out_57_10) );
ms00f80 x_out_57_reg_11_ ( .ck(ispd_clk), .d(n_28015), .o(x_out_57_11) );
ms00f80 x_out_57_reg_12_ ( .ck(ispd_clk), .d(n_28429), .o(x_out_57_12) );
ms00f80 x_out_57_reg_13_ ( .ck(ispd_clk), .d(n_28871), .o(x_out_57_13) );
ms00f80 x_out_57_reg_14_ ( .ck(ispd_clk), .d(n_29211), .o(x_out_57_14) );
ms00f80 x_out_57_reg_15_ ( .ck(ispd_clk), .d(n_29500), .o(x_out_57_15) );
ms00f80 x_out_57_reg_18_ ( .ck(ispd_clk), .d(n_7331), .o(x_out_57_18) );
ms00f80 x_out_57_reg_19_ ( .ck(ispd_clk), .d(n_7386), .o(x_out_57_19) );
ms00f80 x_out_57_reg_1_ ( .ck(ispd_clk), .d(n_15454), .o(x_out_57_1) );
ms00f80 x_out_57_reg_20_ ( .ck(ispd_clk), .d(n_7439), .o(x_out_57_20) );
ms00f80 x_out_57_reg_21_ ( .ck(ispd_clk), .d(n_8373), .o(x_out_57_21) );
ms00f80 x_out_57_reg_22_ ( .ck(ispd_clk), .d(n_10561), .o(x_out_57_22) );
ms00f80 x_out_57_reg_23_ ( .ck(ispd_clk), .d(n_12309), .o(x_out_57_23) );
ms00f80 x_out_57_reg_24_ ( .ck(ispd_clk), .d(n_12961), .o(x_out_57_24) );
ms00f80 x_out_57_reg_25_ ( .ck(ispd_clk), .d(n_13700), .o(x_out_57_25) );
ms00f80 x_out_57_reg_26_ ( .ck(ispd_clk), .d(n_15078), .o(x_out_57_26) );
ms00f80 x_out_57_reg_27_ ( .ck(ispd_clk), .d(n_15722), .o(x_out_57_27) );
ms00f80 x_out_57_reg_28_ ( .ck(ispd_clk), .d(n_16467), .o(x_out_57_28) );
ms00f80 x_out_57_reg_29_ ( .ck(ispd_clk), .d(n_16755), .o(x_out_57_29) );
ms00f80 x_out_57_reg_2_ ( .ck(ispd_clk), .d(n_17190), .o(x_out_57_2) );
ms00f80 x_out_57_reg_30_ ( .ck(ispd_clk), .d(n_17023), .o(x_out_57_30) );
ms00f80 x_out_57_reg_31_ ( .ck(ispd_clk), .d(n_17682), .o(x_out_57_31) );
ms00f80 x_out_57_reg_32_ ( .ck(ispd_clk), .d(n_17638), .o(x_out_57_32) );
ms00f80 x_out_57_reg_33_ ( .ck(ispd_clk), .d(n_17636), .o(x_out_57_33) );
ms00f80 x_out_57_reg_3_ ( .ck(ispd_clk), .d(n_20185), .o(x_out_57_3) );
ms00f80 x_out_57_reg_4_ ( .ck(ispd_clk), .d(n_21198), .o(x_out_57_4) );
ms00f80 x_out_57_reg_5_ ( .ck(ispd_clk), .d(n_22020), .o(x_out_57_5) );
ms00f80 x_out_57_reg_6_ ( .ck(ispd_clk), .d(n_22645), .o(x_out_57_6) );
ms00f80 x_out_57_reg_7_ ( .ck(ispd_clk), .d(n_23940), .o(x_out_57_7) );
ms00f80 x_out_57_reg_8_ ( .ck(ispd_clk), .d(n_25286), .o(x_out_57_8) );
ms00f80 x_out_57_reg_9_ ( .ck(ispd_clk), .d(n_26455), .o(x_out_57_9) );
ms00f80 x_out_58_reg_0_ ( .ck(ispd_clk), .d(n_13991), .o(x_out_58_0) );
ms00f80 x_out_58_reg_10_ ( .ck(ispd_clk), .d(n_28216), .o(x_out_58_10) );
ms00f80 x_out_58_reg_11_ ( .ck(ispd_clk), .d(n_28614), .o(x_out_58_11) );
ms00f80 x_out_58_reg_12_ ( .ck(ispd_clk), .d(n_28921), .o(x_out_58_12) );
ms00f80 x_out_58_reg_13_ ( .ck(ispd_clk), .d(n_29258), .o(x_out_58_13) );
ms00f80 x_out_58_reg_14_ ( .ck(ispd_clk), .d(n_29573), .o(x_out_58_14) );
ms00f80 x_out_58_reg_15_ ( .ck(ispd_clk), .d(n_29668), .o(x_out_58_15) );
ms00f80 x_out_58_reg_18_ ( .ck(ispd_clk), .d(n_7284), .o(x_out_58_18) );
ms00f80 x_out_58_reg_19_ ( .ck(ispd_clk), .d(n_7397), .o(x_out_58_19) );
ms00f80 x_out_58_reg_1_ ( .ck(ispd_clk), .d(n_19158), .o(x_out_58_1) );
ms00f80 x_out_58_reg_20_ ( .ck(ispd_clk), .d(n_6752), .o(x_out_58_20) );
ms00f80 x_out_58_reg_21_ ( .ck(ispd_clk), .d(n_8380), .o(x_out_58_21) );
ms00f80 x_out_58_reg_22_ ( .ck(ispd_clk), .d(n_9277), .o(x_out_58_22) );
ms00f80 x_out_58_reg_23_ ( .ck(ispd_clk), .d(n_10928), .o(x_out_58_23) );
ms00f80 x_out_58_reg_24_ ( .ck(ispd_clk), .d(n_12195), .o(x_out_58_24) );
ms00f80 x_out_58_reg_25_ ( .ck(ispd_clk), .d(n_13272), .o(x_out_58_25) );
ms00f80 x_out_58_reg_26_ ( .ck(ispd_clk), .d(n_14544), .o(x_out_58_26) );
ms00f80 x_out_58_reg_27_ ( .ck(ispd_clk), .d(n_15453), .o(x_out_58_27) );
ms00f80 x_out_58_reg_28_ ( .ck(ispd_clk), .d(n_16439), .o(x_out_58_28) );
ms00f80 x_out_58_reg_29_ ( .ck(ispd_clk), .d(n_16927), .o(x_out_58_29) );
ms00f80 x_out_58_reg_2_ ( .ck(ispd_clk), .d(n_20500), .o(x_out_58_2) );
ms00f80 x_out_58_reg_30_ ( .ck(ispd_clk), .d(n_17316), .o(x_out_58_30) );
ms00f80 x_out_58_reg_31_ ( .ck(ispd_clk), .d(n_17886), .o(x_out_58_31) );
ms00f80 x_out_58_reg_32_ ( .ck(ispd_clk), .d(n_17627), .o(x_out_58_32) );
ms00f80 x_out_58_reg_33_ ( .ck(ispd_clk), .d(n_17629), .o(x_out_58_33) );
ms00f80 x_out_58_reg_3_ ( .ck(ispd_clk), .d(n_21995), .o(x_out_58_3) );
ms00f80 x_out_58_reg_4_ ( .ck(ispd_clk), .d(n_22619), .o(x_out_58_4) );
ms00f80 x_out_58_reg_5_ ( .ck(ispd_clk), .d(n_23318), .o(x_out_58_5) );
ms00f80 x_out_58_reg_6_ ( .ck(ispd_clk), .d(n_24304), .o(x_out_58_6) );
ms00f80 x_out_58_reg_7_ ( .ck(ispd_clk), .d(n_25675), .o(x_out_58_7) );
ms00f80 x_out_58_reg_8_ ( .ck(ispd_clk), .d(n_26532), .o(x_out_58_8) );
ms00f80 x_out_58_reg_9_ ( .ck(ispd_clk), .d(n_27556), .o(x_out_58_9) );
ms00f80 x_out_59_reg_0_ ( .ck(ispd_clk), .d(n_13942), .o(x_out_59_0) );
ms00f80 x_out_59_reg_10_ ( .ck(ispd_clk), .d(n_28215), .o(x_out_59_10) );
ms00f80 x_out_59_reg_11_ ( .ck(ispd_clk), .d(n_28613), .o(x_out_59_11) );
ms00f80 x_out_59_reg_12_ ( .ck(ispd_clk), .d(n_28920), .o(x_out_59_12) );
ms00f80 x_out_59_reg_13_ ( .ck(ispd_clk), .d(n_29257), .o(x_out_59_13) );
ms00f80 x_out_59_reg_14_ ( .ck(ispd_clk), .d(n_29572), .o(x_out_59_14) );
ms00f80 x_out_59_reg_15_ ( .ck(ispd_clk), .d(n_29665), .o(x_out_59_15) );
ms00f80 x_out_59_reg_18_ ( .ck(ispd_clk), .d(n_7588), .o(x_out_59_18) );
ms00f80 x_out_59_reg_19_ ( .ck(ispd_clk), .d(n_7387), .o(x_out_59_19) );
ms00f80 x_out_59_reg_1_ ( .ck(ispd_clk), .d(n_19157), .o(x_out_59_1) );
ms00f80 x_out_59_reg_20_ ( .ck(ispd_clk), .d(n_7536), .o(x_out_59_20) );
ms00f80 x_out_59_reg_21_ ( .ck(ispd_clk), .d(n_8381), .o(x_out_59_21) );
ms00f80 x_out_59_reg_22_ ( .ck(ispd_clk), .d(n_9243), .o(x_out_59_22) );
ms00f80 x_out_59_reg_23_ ( .ck(ispd_clk), .d(n_10925), .o(x_out_59_23) );
ms00f80 x_out_59_reg_24_ ( .ck(ispd_clk), .d(n_12193), .o(x_out_59_24) );
ms00f80 x_out_59_reg_25_ ( .ck(ispd_clk), .d(n_13267), .o(x_out_59_25) );
ms00f80 x_out_59_reg_26_ ( .ck(ispd_clk), .d(n_14523), .o(x_out_59_26) );
ms00f80 x_out_59_reg_27_ ( .ck(ispd_clk), .d(n_15669), .o(x_out_59_27) );
ms00f80 x_out_59_reg_28_ ( .ck(ispd_clk), .d(n_16431), .o(x_out_59_28) );
ms00f80 x_out_59_reg_29_ ( .ck(ispd_clk), .d(n_16924), .o(x_out_59_29) );
ms00f80 x_out_59_reg_2_ ( .ck(ispd_clk), .d(n_20499), .o(x_out_59_2) );
ms00f80 x_out_59_reg_30_ ( .ck(ispd_clk), .d(n_17314), .o(x_out_59_30) );
ms00f80 x_out_59_reg_31_ ( .ck(ispd_clk), .d(n_17885), .o(x_out_59_31) );
ms00f80 x_out_59_reg_32_ ( .ck(ispd_clk), .d(n_17635), .o(x_out_59_32) );
ms00f80 x_out_59_reg_33_ ( .ck(ispd_clk), .d(n_17633), .o(x_out_59_33) );
ms00f80 x_out_59_reg_3_ ( .ck(ispd_clk), .d(n_21994), .o(x_out_59_3) );
ms00f80 x_out_59_reg_4_ ( .ck(ispd_clk), .d(n_22618), .o(x_out_59_4) );
ms00f80 x_out_59_reg_5_ ( .ck(ispd_clk), .d(n_23317), .o(x_out_59_5) );
ms00f80 x_out_59_reg_6_ ( .ck(ispd_clk), .d(n_24303), .o(x_out_59_6) );
ms00f80 x_out_59_reg_7_ ( .ck(ispd_clk), .d(n_25673), .o(x_out_59_7) );
ms00f80 x_out_59_reg_8_ ( .ck(ispd_clk), .d(n_26530), .o(x_out_59_8) );
ms00f80 x_out_59_reg_9_ ( .ck(ispd_clk), .d(n_27554), .o(x_out_59_9) );
ms00f80 x_out_5_reg_0_ ( .ck(ispd_clk), .d(n_16989), .o(x_out_5_0) );
ms00f80 x_out_5_reg_10_ ( .ck(ispd_clk), .d(n_28315), .o(x_out_5_10) );
ms00f80 x_out_5_reg_11_ ( .ck(ispd_clk), .d(n_28684), .o(x_out_5_11) );
ms00f80 x_out_5_reg_12_ ( .ck(ispd_clk), .d(n_29039), .o(x_out_5_12) );
ms00f80 x_out_5_reg_13_ ( .ck(ispd_clk), .d(n_29342), .o(x_out_5_13) );
ms00f80 x_out_5_reg_14_ ( .ck(ispd_clk), .d(n_29620), .o(x_out_5_14) );
ms00f80 x_out_5_reg_15_ ( .ck(ispd_clk), .d(n_29696), .o(x_out_5_15) );
ms00f80 x_out_5_reg_18_ ( .ck(ispd_clk), .d(n_7408), .o(x_out_5_18) );
ms00f80 x_out_5_reg_19_ ( .ck(ispd_clk), .d(n_7438), .o(x_out_5_19) );
ms00f80 x_out_5_reg_1_ ( .ck(ispd_clk), .d(n_18530), .o(x_out_5_1) );
ms00f80 x_out_5_reg_20_ ( .ck(ispd_clk), .d(n_8001), .o(x_out_5_20) );
ms00f80 x_out_5_reg_21_ ( .ck(ispd_clk), .d(n_12311), .o(x_out_5_21) );
ms00f80 x_out_5_reg_22_ ( .ck(ispd_clk), .d(n_13356), .o(x_out_5_22) );
ms00f80 x_out_5_reg_23_ ( .ck(ispd_clk), .d(n_14579), .o(x_out_5_23) );
ms00f80 x_out_5_reg_24_ ( .ck(ispd_clk), .d(n_15980), .o(x_out_5_24) );
ms00f80 x_out_5_reg_25_ ( .ck(ispd_clk), .d(n_16634), .o(x_out_5_25) );
ms00f80 x_out_5_reg_26_ ( .ck(ispd_clk), .d(n_18088), .o(x_out_5_26) );
ms00f80 x_out_5_reg_27_ ( .ck(ispd_clk), .d(n_18674), .o(x_out_5_27) );
ms00f80 x_out_5_reg_28_ ( .ck(ispd_clk), .d(n_20355), .o(x_out_5_28) );
ms00f80 x_out_5_reg_29_ ( .ck(ispd_clk), .d(n_21113), .o(x_out_5_29) );
ms00f80 x_out_5_reg_2_ ( .ck(ispd_clk), .d(n_19828), .o(x_out_5_2) );
ms00f80 x_out_5_reg_30_ ( .ck(ispd_clk), .d(n_22469), .o(x_out_5_30) );
ms00f80 x_out_5_reg_31_ ( .ck(ispd_clk), .d(n_23163), .o(x_out_5_31) );
ms00f80 x_out_5_reg_32_ ( .ck(ispd_clk), .d(n_24721), .o(x_out_5_32) );
ms00f80 x_out_5_reg_33_ ( .ck(ispd_clk), .d(n_24489), .o(x_out_5_33) );
ms00f80 x_out_5_reg_3_ ( .ck(ispd_clk), .d(n_20973), .o(x_out_5_3) );
ms00f80 x_out_5_reg_4_ ( .ck(ispd_clk), .d(n_22066), .o(x_out_5_4) );
ms00f80 x_out_5_reg_5_ ( .ck(ispd_clk), .d(n_23293), .o(x_out_5_5) );
ms00f80 x_out_5_reg_6_ ( .ck(ispd_clk), .d(n_24616), .o(x_out_5_6) );
ms00f80 x_out_5_reg_7_ ( .ck(ispd_clk), .d(n_25896), .o(x_out_5_7) );
ms00f80 x_out_5_reg_8_ ( .ck(ispd_clk), .d(n_26806), .o(x_out_5_8) );
ms00f80 x_out_5_reg_9_ ( .ck(ispd_clk), .d(n_27702), .o(x_out_5_9) );
ms00f80 x_out_60_reg_0_ ( .ck(ispd_clk), .d(n_13986), .o(x_out_60_0) );
ms00f80 x_out_60_reg_10_ ( .ck(ispd_clk), .d(n_27931), .o(x_out_60_10) );
ms00f80 x_out_60_reg_11_ ( .ck(ispd_clk), .d(n_28367), .o(x_out_60_11) );
ms00f80 x_out_60_reg_12_ ( .ck(ispd_clk), .d(n_28752), .o(x_out_60_12) );
ms00f80 x_out_60_reg_13_ ( .ck(ispd_clk), .d(n_29103), .o(x_out_60_13) );
ms00f80 x_out_60_reg_14_ ( .ck(ispd_clk), .d(n_29446), .o(x_out_60_14) );
ms00f80 x_out_60_reg_15_ ( .ck(ispd_clk), .d(n_29650), .o(x_out_60_15) );
ms00f80 x_out_60_reg_18_ ( .ck(ispd_clk), .d(n_7360), .o(x_out_60_18) );
ms00f80 x_out_60_reg_19_ ( .ck(ispd_clk), .d(n_7228), .o(x_out_60_19) );
ms00f80 x_out_60_reg_1_ ( .ck(ispd_clk), .d(n_19156), .o(x_out_60_1) );
ms00f80 x_out_60_reg_20_ ( .ck(ispd_clk), .d(n_7485), .o(x_out_60_20) );
ms00f80 x_out_60_reg_21_ ( .ck(ispd_clk), .d(n_8208), .o(x_out_60_21) );
ms00f80 x_out_60_reg_22_ ( .ck(ispd_clk), .d(n_9274), .o(x_out_60_22) );
ms00f80 x_out_60_reg_23_ ( .ck(ispd_clk), .d(n_10929), .o(x_out_60_23) );
ms00f80 x_out_60_reg_24_ ( .ck(ispd_clk), .d(n_12192), .o(x_out_60_24) );
ms00f80 x_out_60_reg_25_ ( .ck(ispd_clk), .d(n_13271), .o(x_out_60_25) );
ms00f80 x_out_60_reg_26_ ( .ck(ispd_clk), .d(n_14543), .o(x_out_60_26) );
ms00f80 x_out_60_reg_27_ ( .ck(ispd_clk), .d(n_15452), .o(x_out_60_27) );
ms00f80 x_out_60_reg_28_ ( .ck(ispd_clk), .d(n_16437), .o(x_out_60_28) );
ms00f80 x_out_60_reg_29_ ( .ck(ispd_clk), .d(n_16716), .o(x_out_60_29) );
ms00f80 x_out_60_reg_2_ ( .ck(ispd_clk), .d(n_20498), .o(x_out_60_2) );
ms00f80 x_out_60_reg_30_ ( .ck(ispd_clk), .d(n_17604), .o(x_out_60_30) );
ms00f80 x_out_60_reg_31_ ( .ck(ispd_clk), .d(n_17541), .o(x_out_60_31) );
ms00f80 x_out_60_reg_32_ ( .ck(ispd_clk), .d(n_17232), .o(x_out_60_32) );
ms00f80 x_out_60_reg_33_ ( .ck(ispd_clk), .d(n_17234), .o(x_out_60_33) );
ms00f80 x_out_60_reg_3_ ( .ck(ispd_clk), .d(n_21993), .o(x_out_60_3) );
ms00f80 x_out_60_reg_4_ ( .ck(ispd_clk), .d(n_22617), .o(x_out_60_4) );
ms00f80 x_out_60_reg_5_ ( .ck(ispd_clk), .d(n_23314), .o(x_out_60_5) );
ms00f80 x_out_60_reg_6_ ( .ck(ispd_clk), .d(n_24302), .o(x_out_60_6) );
ms00f80 x_out_60_reg_7_ ( .ck(ispd_clk), .d(n_25672), .o(x_out_60_7) );
ms00f80 x_out_60_reg_8_ ( .ck(ispd_clk), .d(n_26238), .o(x_out_60_8) );
ms00f80 x_out_60_reg_9_ ( .ck(ispd_clk), .d(n_27155), .o(x_out_60_9) );
ms00f80 x_out_61_reg_0_ ( .ck(ispd_clk), .d(n_14664), .o(x_out_61_0) );
ms00f80 x_out_61_reg_10_ ( .ck(ispd_clk), .d(n_28214), .o(x_out_61_10) );
ms00f80 x_out_61_reg_11_ ( .ck(ispd_clk), .d(n_28612), .o(x_out_61_11) );
ms00f80 x_out_61_reg_12_ ( .ck(ispd_clk), .d(n_28919), .o(x_out_61_12) );
ms00f80 x_out_61_reg_13_ ( .ck(ispd_clk), .d(n_29254), .o(x_out_61_13) );
ms00f80 x_out_61_reg_14_ ( .ck(ispd_clk), .d(n_29570), .o(x_out_61_14) );
ms00f80 x_out_61_reg_15_ ( .ck(ispd_clk), .d(n_29682), .o(x_out_61_15) );
ms00f80 x_out_61_reg_18_ ( .ck(ispd_clk), .d(n_7366), .o(x_out_61_18) );
ms00f80 x_out_61_reg_19_ ( .ck(ispd_clk), .d(n_7395), .o(x_out_61_19) );
ms00f80 x_out_61_reg_1_ ( .ck(ispd_clk), .d(n_19155), .o(x_out_61_1) );
ms00f80 x_out_61_reg_20_ ( .ck(ispd_clk), .d(n_7465), .o(x_out_61_20) );
ms00f80 x_out_61_reg_21_ ( .ck(ispd_clk), .d(n_8383), .o(x_out_61_21) );
ms00f80 x_out_61_reg_22_ ( .ck(ispd_clk), .d(n_9273), .o(x_out_61_22) );
ms00f80 x_out_61_reg_23_ ( .ck(ispd_clk), .d(n_10927), .o(x_out_61_23) );
ms00f80 x_out_61_reg_24_ ( .ck(ispd_clk), .d(n_12189), .o(x_out_61_24) );
ms00f80 x_out_61_reg_25_ ( .ck(ispd_clk), .d(n_13270), .o(x_out_61_25) );
ms00f80 x_out_61_reg_26_ ( .ck(ispd_clk), .d(n_14542), .o(x_out_61_26) );
ms00f80 x_out_61_reg_27_ ( .ck(ispd_clk), .d(n_15451), .o(x_out_61_27) );
ms00f80 x_out_61_reg_28_ ( .ck(ispd_clk), .d(n_16436), .o(x_out_61_28) );
ms00f80 x_out_61_reg_29_ ( .ck(ispd_clk), .d(n_16718), .o(x_out_61_29) );
ms00f80 x_out_61_reg_2_ ( .ck(ispd_clk), .d(n_20497), .o(x_out_61_2) );
ms00f80 x_out_61_reg_30_ ( .ck(ispd_clk), .d(n_17603), .o(x_out_61_30) );
ms00f80 x_out_61_reg_31_ ( .ck(ispd_clk), .d(n_17539), .o(x_out_61_31) );
ms00f80 x_out_61_reg_32_ ( .ck(ispd_clk), .d(n_17262), .o(x_out_61_32) );
ms00f80 x_out_61_reg_33_ ( .ck(ispd_clk), .d(n_17260), .o(x_out_61_33) );
ms00f80 x_out_61_reg_3_ ( .ck(ispd_clk), .d(n_21992), .o(x_out_61_3) );
ms00f80 x_out_61_reg_4_ ( .ck(ispd_clk), .d(n_22616), .o(x_out_61_4) );
ms00f80 x_out_61_reg_5_ ( .ck(ispd_clk), .d(n_23313), .o(x_out_61_5) );
ms00f80 x_out_61_reg_6_ ( .ck(ispd_clk), .d(n_24301), .o(x_out_61_6) );
ms00f80 x_out_61_reg_7_ ( .ck(ispd_clk), .d(n_25671), .o(x_out_61_7) );
ms00f80 x_out_61_reg_8_ ( .ck(ispd_clk), .d(n_26528), .o(x_out_61_8) );
ms00f80 x_out_61_reg_9_ ( .ck(ispd_clk), .d(n_27553), .o(x_out_61_9) );
ms00f80 x_out_62_reg_0_ ( .ck(ispd_clk), .d(n_14790), .o(x_out_62_0) );
ms00f80 x_out_62_reg_10_ ( .ck(ispd_clk), .d(n_28213), .o(x_out_62_10) );
ms00f80 x_out_62_reg_11_ ( .ck(ispd_clk), .d(n_28611), .o(x_out_62_11) );
ms00f80 x_out_62_reg_12_ ( .ck(ispd_clk), .d(n_28917), .o(x_out_62_12) );
ms00f80 x_out_62_reg_13_ ( .ck(ispd_clk), .d(n_29253), .o(x_out_62_13) );
ms00f80 x_out_62_reg_14_ ( .ck(ispd_clk), .d(n_29569), .o(x_out_62_14) );
ms00f80 x_out_62_reg_15_ ( .ck(ispd_clk), .d(n_29680), .o(x_out_62_15) );
ms00f80 x_out_62_reg_18_ ( .ck(ispd_clk), .d(n_8028), .o(x_out_62_18) );
ms00f80 x_out_62_reg_19_ ( .ck(ispd_clk), .d(n_7398), .o(x_out_62_19) );
ms00f80 x_out_62_reg_1_ ( .ck(ispd_clk), .d(n_19154), .o(x_out_62_1) );
ms00f80 x_out_62_reg_20_ ( .ck(ispd_clk), .d(n_7493), .o(x_out_62_20) );
ms00f80 x_out_62_reg_21_ ( .ck(ispd_clk), .d(n_8382), .o(x_out_62_21) );
ms00f80 x_out_62_reg_22_ ( .ck(ispd_clk), .d(n_9268), .o(x_out_62_22) );
ms00f80 x_out_62_reg_23_ ( .ck(ispd_clk), .d(n_10926), .o(x_out_62_23) );
ms00f80 x_out_62_reg_24_ ( .ck(ispd_clk), .d(n_12188), .o(x_out_62_24) );
ms00f80 x_out_62_reg_25_ ( .ck(ispd_clk), .d(n_13269), .o(x_out_62_25) );
ms00f80 x_out_62_reg_26_ ( .ck(ispd_clk), .d(n_14541), .o(x_out_62_26) );
ms00f80 x_out_62_reg_27_ ( .ck(ispd_clk), .d(n_15450), .o(x_out_62_27) );
ms00f80 x_out_62_reg_28_ ( .ck(ispd_clk), .d(n_16435), .o(x_out_62_28) );
ms00f80 x_out_62_reg_29_ ( .ck(ispd_clk), .d(n_16926), .o(x_out_62_29) );
ms00f80 x_out_62_reg_2_ ( .ck(ispd_clk), .d(n_20496), .o(x_out_62_2) );
ms00f80 x_out_62_reg_30_ ( .ck(ispd_clk), .d(n_17315), .o(x_out_62_30) );
ms00f80 x_out_62_reg_31_ ( .ck(ispd_clk), .d(n_17887), .o(x_out_62_31) );
ms00f80 x_out_62_reg_32_ ( .ck(ispd_clk), .d(n_17632), .o(x_out_62_32) );
ms00f80 x_out_62_reg_33_ ( .ck(ispd_clk), .d(n_17630), .o(x_out_62_33) );
ms00f80 x_out_62_reg_3_ ( .ck(ispd_clk), .d(n_21991), .o(x_out_62_3) );
ms00f80 x_out_62_reg_4_ ( .ck(ispd_clk), .d(n_22614), .o(x_out_62_4) );
ms00f80 x_out_62_reg_5_ ( .ck(ispd_clk), .d(n_23312), .o(x_out_62_5) );
ms00f80 x_out_62_reg_6_ ( .ck(ispd_clk), .d(n_24300), .o(x_out_62_6) );
ms00f80 x_out_62_reg_7_ ( .ck(ispd_clk), .d(n_25670), .o(x_out_62_7) );
ms00f80 x_out_62_reg_8_ ( .ck(ispd_clk), .d(n_26526), .o(x_out_62_8) );
ms00f80 x_out_62_reg_9_ ( .ck(ispd_clk), .d(n_27552), .o(x_out_62_9) );
ms00f80 x_out_63_reg_0_ ( .ck(ispd_clk), .d(n_14758), .o(x_out_63_0) );
ms00f80 x_out_63_reg_10_ ( .ck(ispd_clk), .d(n_28212), .o(x_out_63_10) );
ms00f80 x_out_63_reg_11_ ( .ck(ispd_clk), .d(n_28609), .o(x_out_63_11) );
ms00f80 x_out_63_reg_12_ ( .ck(ispd_clk), .d(n_28915), .o(x_out_63_12) );
ms00f80 x_out_63_reg_13_ ( .ck(ispd_clk), .d(n_29252), .o(x_out_63_13) );
ms00f80 x_out_63_reg_14_ ( .ck(ispd_clk), .d(n_29566), .o(x_out_63_14) );
ms00f80 x_out_63_reg_15_ ( .ck(ispd_clk), .d(n_29678), .o(x_out_63_15) );
ms00f80 x_out_63_reg_18_ ( .ck(ispd_clk), .d(n_7348), .o(x_out_63_18) );
ms00f80 x_out_63_reg_19_ ( .ck(ispd_clk), .d(n_7227), .o(x_out_63_19) );
ms00f80 x_out_63_reg_1_ ( .ck(ispd_clk), .d(n_19153), .o(x_out_63_1) );
ms00f80 x_out_63_reg_20_ ( .ck(ispd_clk), .d(n_7444), .o(x_out_63_20) );
ms00f80 x_out_63_reg_21_ ( .ck(ispd_clk), .d(n_7373), .o(x_out_63_21) );
ms00f80 x_out_63_reg_22_ ( .ck(ispd_clk), .d(n_9236), .o(x_out_63_22) );
ms00f80 x_out_63_reg_23_ ( .ck(ispd_clk), .d(n_10924), .o(x_out_63_23) );
ms00f80 x_out_63_reg_24_ ( .ck(ispd_clk), .d(n_12181), .o(x_out_63_24) );
ms00f80 x_out_63_reg_25_ ( .ck(ispd_clk), .d(n_13268), .o(x_out_63_25) );
ms00f80 x_out_63_reg_26_ ( .ck(ispd_clk), .d(n_14540), .o(x_out_63_26) );
ms00f80 x_out_63_reg_27_ ( .ck(ispd_clk), .d(n_15449), .o(x_out_63_27) );
ms00f80 x_out_63_reg_28_ ( .ck(ispd_clk), .d(n_16434), .o(x_out_63_28) );
ms00f80 x_out_63_reg_29_ ( .ck(ispd_clk), .d(n_16717), .o(x_out_63_29) );
ms00f80 x_out_63_reg_2_ ( .ck(ispd_clk), .d(n_20495), .o(x_out_63_2) );
ms00f80 x_out_63_reg_30_ ( .ck(ispd_clk), .d(n_17602), .o(x_out_63_30) );
ms00f80 x_out_63_reg_31_ ( .ck(ispd_clk), .d(n_17540), .o(x_out_63_31) );
ms00f80 x_out_63_reg_32_ ( .ck(ispd_clk), .d(n_17259), .o(x_out_63_32) );
ms00f80 x_out_63_reg_33_ ( .ck(ispd_clk), .d(n_17257), .o(x_out_63_33) );
ms00f80 x_out_63_reg_3_ ( .ck(ispd_clk), .d(n_21990), .o(x_out_63_3) );
ms00f80 x_out_63_reg_4_ ( .ck(ispd_clk), .d(n_22613), .o(x_out_63_4) );
ms00f80 x_out_63_reg_5_ ( .ck(ispd_clk), .d(n_23311), .o(x_out_63_5) );
ms00f80 x_out_63_reg_6_ ( .ck(ispd_clk), .d(n_24299), .o(x_out_63_6) );
ms00f80 x_out_63_reg_7_ ( .ck(ispd_clk), .d(n_25669), .o(x_out_63_7) );
ms00f80 x_out_63_reg_8_ ( .ck(ispd_clk), .d(n_26524), .o(x_out_63_8) );
ms00f80 x_out_63_reg_9_ ( .ck(ispd_clk), .d(n_27551), .o(x_out_63_9) );
ms00f80 x_out_6_reg_0_ ( .ck(ispd_clk), .d(n_14436), .o(x_out_6_0) );
ms00f80 x_out_6_reg_10_ ( .ck(ispd_clk), .d(n_26453), .o(x_out_6_10) );
ms00f80 x_out_6_reg_11_ ( .ck(ispd_clk), .d(n_27265), .o(x_out_6_11) );
ms00f80 x_out_6_reg_12_ ( .ck(ispd_clk), .d(n_28013), .o(x_out_6_12) );
ms00f80 x_out_6_reg_13_ ( .ck(ispd_clk), .d(n_28427), .o(x_out_6_13) );
ms00f80 x_out_6_reg_14_ ( .ck(ispd_clk), .d(n_28870), .o(x_out_6_14) );
ms00f80 x_out_6_reg_15_ ( .ck(ispd_clk), .d(n_29210), .o(x_out_6_15) );
ms00f80 x_out_6_reg_18_ ( .ck(ispd_clk), .d(n_17225), .o(x_out_6_18) );
ms00f80 x_out_6_reg_19_ ( .ck(ispd_clk), .d(n_17622), .o(x_out_6_19) );
ms00f80 x_out_6_reg_1_ ( .ck(ispd_clk), .d(n_15939), .o(x_out_6_1) );
ms00f80 x_out_6_reg_20_ ( .ck(ispd_clk), .d(n_18850), .o(x_out_6_20) );
ms00f80 x_out_6_reg_21_ ( .ck(ispd_clk), .d(n_19559), .o(x_out_6_21) );
ms00f80 x_out_6_reg_22_ ( .ck(ispd_clk), .d(n_21008), .o(x_out_6_22) );
ms00f80 x_out_6_reg_23_ ( .ck(ispd_clk), .d(n_21453), .o(x_out_6_23) );
ms00f80 x_out_6_reg_24_ ( .ck(ispd_clk), .d(n_22754), .o(x_out_6_24) );
ms00f80 x_out_6_reg_25_ ( .ck(ispd_clk), .d(n_23455), .o(x_out_6_25) );
ms00f80 x_out_6_reg_26_ ( .ck(ispd_clk), .d(n_24714), .o(x_out_6_26) );
ms00f80 x_out_6_reg_27_ ( .ck(ispd_clk), .d(n_25135), .o(x_out_6_27) );
ms00f80 x_out_6_reg_28_ ( .ck(ispd_clk), .d(n_26327), .o(x_out_6_28) );
ms00f80 x_out_6_reg_29_ ( .ck(ispd_clk), .d(n_26816), .o(x_out_6_29) );
ms00f80 x_out_6_reg_2_ ( .ck(ispd_clk), .d(n_17079), .o(x_out_6_2) );
ms00f80 x_out_6_reg_30_ ( .ck(ispd_clk), .d(n_27776), .o(x_out_6_30) );
ms00f80 x_out_6_reg_31_ ( .ck(ispd_clk), .d(n_28144), .o(x_out_6_31) );
ms00f80 x_out_6_reg_32_ ( .ck(ispd_clk), .d(n_28494), .o(x_out_6_32) );
ms00f80 x_out_6_reg_33_ ( .ck(ispd_clk), .d(n_28763), .o(x_out_6_33) );
ms00f80 x_out_6_reg_3_ ( .ck(ispd_clk), .d(n_18411), .o(x_out_6_3) );
ms00f80 x_out_6_reg_4_ ( .ck(ispd_clk), .d(n_18848), .o(x_out_6_4) );
ms00f80 x_out_6_reg_5_ ( .ck(ispd_clk), .d(n_20225), .o(x_out_6_5) );
ms00f80 x_out_6_reg_6_ ( .ck(ispd_clk), .d(n_21644), .o(x_out_6_6) );
ms00f80 x_out_6_reg_7_ ( .ck(ispd_clk), .d(n_22644), .o(x_out_6_7) );
ms00f80 x_out_6_reg_8_ ( .ck(ispd_clk), .d(n_23939), .o(x_out_6_8) );
ms00f80 x_out_6_reg_9_ ( .ck(ispd_clk), .d(n_25284), .o(x_out_6_9) );
ms00f80 x_out_7_reg_0_ ( .ck(ispd_clk), .d(n_13984), .o(x_out_7_0) );
ms00f80 x_out_7_reg_10_ ( .ck(ispd_clk), .d(n_26800), .o(x_out_7_10) );
ms00f80 x_out_7_reg_11_ ( .ck(ispd_clk), .d(n_27700), .o(x_out_7_11) );
ms00f80 x_out_7_reg_12_ ( .ck(ispd_clk), .d(n_28310), .o(x_out_7_12) );
ms00f80 x_out_7_reg_13_ ( .ck(ispd_clk), .d(n_28606), .o(x_out_7_13) );
ms00f80 x_out_7_reg_14_ ( .ck(ispd_clk), .d(n_28830), .o(x_out_7_14) );
ms00f80 x_out_7_reg_15_ ( .ck(ispd_clk), .d(n_29176), .o(x_out_7_15) );
ms00f80 x_out_7_reg_18_ ( .ck(ispd_clk), .d(n_14633), .o(x_out_7_18) );
ms00f80 x_out_7_reg_19_ ( .ck(ispd_clk), .d(n_16078), .o(x_out_7_19) );
ms00f80 x_out_7_reg_1_ ( .ck(ispd_clk), .d(n_16556), .o(x_out_7_1) );
ms00f80 x_out_7_reg_20_ ( .ck(ispd_clk), .d(n_15936), .o(x_out_7_20) );
ms00f80 x_out_7_reg_21_ ( .ck(ispd_clk), .d(n_16846), .o(x_out_7_21) );
ms00f80 x_out_7_reg_22_ ( .ck(ispd_clk), .d(n_18017), .o(x_out_7_22) );
ms00f80 x_out_7_reg_23_ ( .ck(ispd_clk), .d(n_18646), .o(x_out_7_23) );
ms00f80 x_out_7_reg_24_ ( .ck(ispd_clk), .d(n_19996), .o(x_out_7_24) );
ms00f80 x_out_7_reg_25_ ( .ck(ispd_clk), .d(n_20442), .o(x_out_7_25) );
ms00f80 x_out_7_reg_26_ ( .ck(ispd_clk), .d(n_21906), .o(x_out_7_26) );
ms00f80 x_out_7_reg_27_ ( .ck(ispd_clk), .d(n_22554), .o(x_out_7_27) );
ms00f80 x_out_7_reg_28_ ( .ck(ispd_clk), .d(n_23814), .o(x_out_7_28) );
ms00f80 x_out_7_reg_29_ ( .ck(ispd_clk), .d(n_24180), .o(x_out_7_29) );
ms00f80 x_out_7_reg_2_ ( .ck(ispd_clk), .d(n_18149), .o(x_out_7_2) );
ms00f80 x_out_7_reg_30_ ( .ck(ispd_clk), .d(n_25524), .o(x_out_7_30) );
ms00f80 x_out_7_reg_31_ ( .ck(ispd_clk), .d(n_26178), .o(x_out_7_31) );
ms00f80 x_out_7_reg_32_ ( .ck(ispd_clk), .d(n_27370), .o(x_out_7_32) );
ms00f80 x_out_7_reg_33_ ( .ck(ispd_clk), .d(n_27609), .o(x_out_7_33) );
ms00f80 x_out_7_reg_3_ ( .ck(ispd_clk), .d(n_18526), .o(x_out_7_3) );
ms00f80 x_out_7_reg_4_ ( .ck(ispd_clk), .d(n_19838), .o(x_out_7_4) );
ms00f80 x_out_7_reg_5_ ( .ck(ispd_clk), .d(n_20969), .o(x_out_7_5) );
ms00f80 x_out_7_reg_6_ ( .ck(ispd_clk), .d(n_22064), .o(x_out_7_6) );
ms00f80 x_out_7_reg_7_ ( .ck(ispd_clk), .d(n_23309), .o(x_out_7_7) );
ms00f80 x_out_7_reg_8_ ( .ck(ispd_clk), .d(n_24611), .o(x_out_7_8) );
ms00f80 x_out_7_reg_9_ ( .ck(ispd_clk), .d(n_25893), .o(x_out_7_9) );
ms00f80 x_out_8_reg_0_ ( .ck(ispd_clk), .d(n_7413), .o(x_out_8_0) );
ms00f80 x_out_8_reg_10_ ( .ck(ispd_clk), .d(n_22108), .o(x_out_8_10) );
ms00f80 x_out_8_reg_11_ ( .ck(ispd_clk), .d(n_23371), .o(x_out_8_11) );
ms00f80 x_out_8_reg_12_ ( .ck(ispd_clk), .d(n_24667), .o(x_out_8_12) );
ms00f80 x_out_8_reg_13_ ( .ck(ispd_clk), .d(n_25705), .o(x_out_8_13) );
ms00f80 x_out_8_reg_14_ ( .ck(ispd_clk), .d(n_26185), .o(x_out_8_14) );
ms00f80 x_out_8_reg_15_ ( .ck(ispd_clk), .d(n_26850), .o(x_out_8_15) );
ms00f80 x_out_8_reg_18_ ( .ck(ispd_clk), .d(n_14629), .o(x_out_8_18) );
ms00f80 x_out_8_reg_19_ ( .ck(ispd_clk), .d(n_15215), .o(x_out_8_19) );
ms00f80 x_out_8_reg_1_ ( .ck(ispd_clk), .d(n_8000), .o(x_out_8_1) );
ms00f80 x_out_8_reg_20_ ( .ck(ispd_clk), .d(n_15938), .o(x_out_8_20) );
ms00f80 x_out_8_reg_21_ ( .ck(ispd_clk), .d(n_16610), .o(x_out_8_21) );
ms00f80 x_out_8_reg_22_ ( .ck(ispd_clk), .d(n_17778), .o(x_out_8_22) );
ms00f80 x_out_8_reg_23_ ( .ck(ispd_clk), .d(n_18369), .o(x_out_8_23) );
ms00f80 x_out_8_reg_24_ ( .ck(ispd_clk), .d(n_19655), .o(x_out_8_24) );
ms00f80 x_out_8_reg_25_ ( .ck(ispd_clk), .d(n_20084), .o(x_out_8_25) );
ms00f80 x_out_8_reg_26_ ( .ck(ispd_clk), .d(n_21542), .o(x_out_8_26) );
ms00f80 x_out_8_reg_27_ ( .ck(ispd_clk), .d(n_22249), .o(x_out_8_27) );
ms00f80 x_out_8_reg_28_ ( .ck(ispd_clk), .d(n_23549), .o(x_out_8_28) );
ms00f80 x_out_8_reg_29_ ( .ck(ispd_clk), .d(n_23885), .o(x_out_8_29) );
ms00f80 x_out_8_reg_2_ ( .ck(ispd_clk), .d(n_10125), .o(x_out_8_2) );
ms00f80 x_out_8_reg_30_ ( .ck(ispd_clk), .d(n_25254), .o(x_out_8_30) );
ms00f80 x_out_8_reg_31_ ( .ck(ispd_clk), .d(n_25931), .o(x_out_8_31) );
ms00f80 x_out_8_reg_32_ ( .ck(ispd_clk), .d(n_27165), .o(x_out_8_32) );
ms00f80 x_out_8_reg_33_ ( .ck(ispd_clk), .d(n_27503), .o(x_out_8_33) );
ms00f80 x_out_8_reg_3_ ( .ck(ispd_clk), .d(n_12241), .o(x_out_8_3) );
ms00f80 x_out_8_reg_4_ ( .ck(ispd_clk), .d(n_14577), .o(x_out_8_4) );
ms00f80 x_out_8_reg_5_ ( .ck(ispd_clk), .d(n_15979), .o(x_out_8_5) );
ms00f80 x_out_8_reg_6_ ( .ck(ispd_clk), .d(n_17115), .o(x_out_8_6) );
ms00f80 x_out_8_reg_7_ ( .ck(ispd_clk), .d(n_18323), .o(x_out_8_7) );
ms00f80 x_out_8_reg_8_ ( .ck(ispd_clk), .d(n_19558), .o(x_out_8_8) );
ms00f80 x_out_8_reg_9_ ( .ck(ispd_clk), .d(n_21006), .o(x_out_8_9) );
ms00f80 x_out_9_reg_0_ ( .ck(ispd_clk), .d(n_16987), .o(x_out_9_0) );
ms00f80 x_out_9_reg_10_ ( .ck(ispd_clk), .d(n_28210), .o(x_out_9_10) );
ms00f80 x_out_9_reg_11_ ( .ck(ispd_clk), .d(n_28604), .o(x_out_9_11) );
ms00f80 x_out_9_reg_12_ ( .ck(ispd_clk), .d(n_28914), .o(x_out_9_12) );
ms00f80 x_out_9_reg_13_ ( .ck(ispd_clk), .d(n_29305), .o(x_out_9_13) );
ms00f80 x_out_9_reg_14_ ( .ck(ispd_clk), .d(n_29368), .o(x_out_9_14) );
ms00f80 x_out_9_reg_15_ ( .ck(ispd_clk), .d(n_29631), .o(x_out_9_15) );
ms00f80 x_out_9_reg_18_ ( .ck(ispd_clk), .d(n_14631), .o(x_out_9_18) );
ms00f80 x_out_9_reg_19_ ( .ck(ispd_clk), .d(n_15203), .o(x_out_9_19) );
ms00f80 x_out_9_reg_1_ ( .ck(ispd_clk), .d(n_19749), .o(x_out_9_1) );
ms00f80 x_out_9_reg_20_ ( .ck(ispd_clk), .d(n_15934), .o(x_out_9_20) );
ms00f80 x_out_9_reg_21_ ( .ck(ispd_clk), .d(n_17081), .o(x_out_9_21) );
ms00f80 x_out_9_reg_22_ ( .ck(ispd_clk), .d(n_17776), .o(x_out_9_22) );
ms00f80 x_out_9_reg_23_ ( .ck(ispd_clk), .d(n_18989), .o(x_out_9_23) );
ms00f80 x_out_9_reg_24_ ( .ck(ispd_clk), .d(n_19653), .o(x_out_9_24) );
ms00f80 x_out_9_reg_25_ ( .ck(ispd_clk), .d(n_20802), .o(x_out_9_25) );
ms00f80 x_out_9_reg_26_ ( .ck(ispd_clk), .d(n_21540), .o(x_out_9_26) );
ms00f80 x_out_9_reg_27_ ( .ck(ispd_clk), .d(n_22851), .o(x_out_9_27) );
ms00f80 x_out_9_reg_28_ ( .ck(ispd_clk), .d(n_23547), .o(x_out_9_28) );
ms00f80 x_out_9_reg_29_ ( .ck(ispd_clk), .d(n_24494), .o(x_out_9_29) );
ms00f80 x_out_9_reg_2_ ( .ck(ispd_clk), .d(n_20494), .o(x_out_9_2) );
ms00f80 x_out_9_reg_30_ ( .ck(ispd_clk), .d(n_25249), .o(x_out_9_30) );
ms00f80 x_out_9_reg_31_ ( .ck(ispd_clk), .d(n_26444), .o(x_out_9_31) );
ms00f80 x_out_9_reg_32_ ( .ck(ispd_clk), .d(n_27368), .o(x_out_9_32) );
ms00f80 x_out_9_reg_33_ ( .ck(ispd_clk), .d(n_27208), .o(x_out_9_33) );
ms00f80 x_out_9_reg_3_ ( .ck(ispd_clk), .d(n_21989), .o(x_out_9_3) );
ms00f80 x_out_9_reg_4_ ( .ck(ispd_clk), .d(n_22612), .o(x_out_9_4) );
ms00f80 x_out_9_reg_5_ ( .ck(ispd_clk), .d(n_23612), .o(x_out_9_5) );
ms00f80 x_out_9_reg_6_ ( .ck(ispd_clk), .d(n_24921), .o(x_out_9_6) );
ms00f80 x_out_9_reg_7_ ( .ck(ispd_clk), .d(n_26134), .o(x_out_9_7) );
ms00f80 x_out_9_reg_8_ ( .ck(ispd_clk), .d(n_26794), .o(x_out_9_8) );
ms00f80 x_out_9_reg_9_ ( .ck(ispd_clk), .d(n_27550), .o(x_out_9_9) );

endmodule
